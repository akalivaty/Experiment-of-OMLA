//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(KEYINPUT64), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n206), .B1(new_n207), .B2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n209), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT65), .Z(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI22_X1  g0022(.A1(new_n220), .A2(new_n221), .B1(new_n203), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n219), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G87), .ZN(new_n227));
  INV_X1    g0027(.A(G250), .ZN(new_n228));
  INV_X1    g0028(.A(G116), .ZN(new_n229));
  INV_X1    g0029(.A(G270), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(G257), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n202), .A2(new_n232), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n207), .B1(KEYINPUT67), .B2(new_n215), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n215), .A2(KEYINPUT67), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(G1), .A2(G13), .ZN(new_n237));
  INV_X1    g0037(.A(G20), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g0039(.A1(G58), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  AOI211_X1 g0043(.A(new_n214), .B(new_n236), .C1(new_n239), .C2(new_n243), .ZN(G361));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G238), .B(G244), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT68), .B(G250), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G257), .ZN(new_n250));
  XOR2_X1   g0050(.A(G264), .B(G270), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G358));
  XOR2_X1   g0053(.A(G68), .B(G77), .Z(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G58), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(G107), .B(G116), .ZN(new_n257));
  XNOR2_X1  g0057(.A(G87), .B(G97), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XOR2_X1   g0059(.A(new_n256), .B(new_n259), .Z(G351));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n238), .A2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G13), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n237), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(KEYINPUT70), .ZN(new_n269));
  AND3_X1   g0069(.A1(new_n266), .A2(KEYINPUT70), .A3(new_n237), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n269), .A2(new_n263), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n265), .B1(new_n271), .B2(new_n262), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n238), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT7), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n238), .A4(new_n277), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(KEYINPUT75), .A3(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n281), .A2(KEYINPUT75), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G68), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT76), .ZN(new_n285));
  XNOR2_X1  g0085(.A(G58), .B(G68), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n286), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT76), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n282), .A2(new_n283), .A3(new_n289), .A4(G68), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n285), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT16), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G68), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n280), .B2(new_n281), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(KEYINPUT16), .A3(new_n288), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n267), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n273), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G41), .ZN(new_n301));
  OAI211_X1 g0101(.A(G1), .B(G13), .C1(new_n275), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n276), .A2(new_n277), .ZN(new_n303));
  INV_X1    g0103(.A(G223), .ZN(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n303), .B(new_n306), .C1(G226), .C2(new_n305), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G87), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G1), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G41), .B2(G45), .ZN(new_n311));
  INV_X1    g0111(.A(G274), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n302), .A2(new_n311), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(new_n221), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n309), .A2(G190), .A3(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n309), .A2(new_n315), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G200), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT17), .B1(new_n300), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n298), .B1(new_n291), .B2(new_n292), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT17), .ZN(new_n324));
  NOR4_X1   g0124(.A1(new_n323), .A2(new_n324), .A3(new_n320), .A4(new_n273), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT18), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n317), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(G179), .B2(new_n317), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n327), .B1(new_n300), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n317), .A2(G179), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n328), .B2(new_n317), .ZN(new_n333));
  OAI211_X1 g0133(.A(KEYINPUT18), .B(new_n333), .C1(new_n323), .C2(new_n273), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G238), .A2(G1698), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n303), .B(new_n336), .C1(new_n221), .C2(G1698), .ZN(new_n337));
  INV_X1    g0137(.A(new_n302), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(G107), .C2(new_n303), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(new_n313), .C1(new_n218), .C2(new_n314), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n340), .A2(G179), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n262), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n238), .A2(G33), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT15), .B(G87), .Z(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n342), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n264), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n346), .A2(new_n267), .B1(new_n217), .B2(new_n347), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n267), .A2(new_n263), .A3(new_n217), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT72), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n340), .A2(new_n328), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n341), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n326), .A2(new_n335), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n305), .A2(G222), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n303), .B(new_n355), .C1(new_n304), .C2(new_n305), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(G77), .B2(new_n303), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT69), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n302), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n358), .B2(new_n357), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n302), .A2(G226), .A3(new_n311), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n313), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G190), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(G20), .B1(new_n241), .B2(G50), .ZN(new_n365));
  INV_X1    g0165(.A(G150), .ZN(new_n366));
  INV_X1    g0166(.A(new_n287), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n365), .B1(new_n366), .B2(new_n367), .C1(new_n343), .C2(new_n261), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n271), .A2(G50), .B1(new_n368), .B2(new_n267), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(G50), .B2(new_n264), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT9), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n362), .A2(G200), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n370), .A2(new_n371), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n364), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT10), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n362), .A2(G179), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n328), .B2(new_n362), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n370), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G97), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n221), .A2(G1698), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(G226), .B2(G1698), .ZN(new_n383));
  AND2_X1   g0183(.A1(KEYINPUT3), .A2(G33), .ZN(new_n384));
  NOR2_X1   g0184(.A1(KEYINPUT3), .A2(G33), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n381), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n338), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n302), .A2(G238), .A3(new_n311), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n389), .A2(KEYINPUT73), .A3(new_n313), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT73), .B1(new_n389), .B2(new_n313), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n388), .B(new_n394), .C1(new_n390), .C2(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT74), .A3(G169), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(G179), .A3(new_n395), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n396), .A2(KEYINPUT74), .A3(new_n400), .A4(G169), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G50), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n367), .A2(new_n403), .B1(new_n238), .B2(G68), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n343), .A2(new_n217), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n267), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT11), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n267), .A2(new_n263), .A3(new_n294), .ZN(new_n408));
  OR3_X1    g0208(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n402), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n411), .B(new_n407), .C1(new_n396), .C2(new_n363), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n319), .B1(new_n393), .B2(new_n395), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n340), .A2(new_n363), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT71), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n351), .B1(G200), .B2(new_n340), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NOR4_X1   g0223(.A1(new_n354), .A2(new_n380), .A3(new_n418), .A4(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G283), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n275), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n305), .B1(new_n276), .B2(new_n277), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n426), .B1(new_n427), .B2(G250), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n305), .B1(new_n384), .B2(new_n385), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT79), .ZN(new_n430));
  OAI21_X1  g0230(.A(G244), .B1(new_n430), .B2(KEYINPUT4), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT4), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n429), .A2(new_n431), .B1(KEYINPUT79), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n431), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n432), .A2(KEYINPUT79), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n434), .A2(new_n303), .A3(new_n305), .A4(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n428), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n338), .ZN(new_n438));
  INV_X1    g0238(.A(G45), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(G1), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  AND2_X1   g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n440), .B(G274), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n442), .B2(new_n441), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n302), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n445), .B2(new_n232), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n438), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT80), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n437), .B2(new_n338), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT80), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(G200), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n347), .A2(new_n202), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n310), .A2(G33), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n268), .A2(new_n264), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n454), .B1(new_n456), .B2(new_n202), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n282), .A2(G107), .A3(new_n283), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n287), .A2(G77), .ZN(new_n459));
  XOR2_X1   g0259(.A(KEYINPUT77), .B(KEYINPUT6), .Z(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT78), .B(G97), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n460), .A2(G107), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(G97), .B(G107), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n458), .B(new_n459), .C1(new_n465), .C2(new_n238), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n457), .B1(new_n466), .B2(new_n267), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n450), .A2(G190), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n453), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n218), .A2(G1698), .ZN(new_n470));
  OAI221_X1 g0270(.A(new_n470), .B1(G238), .B2(G1698), .C1(new_n384), .C2(new_n385), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G116), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n338), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n440), .A2(new_n312), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n228), .B1(new_n439), .B2(G1), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n302), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G200), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n344), .A2(new_n264), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(G20), .B1(new_n276), .B2(new_n277), .ZN(new_n482));
  NOR2_X1   g0282(.A1(G87), .A2(G107), .ZN(new_n483));
  AND2_X1   g0283(.A1(KEYINPUT78), .A2(G97), .ZN(new_n484));
  NOR2_X1   g0284(.A1(KEYINPUT78), .A2(G97), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT19), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n238), .B1(new_n381), .B2(new_n487), .ZN(new_n488));
  AOI22_X1  g0288(.A1(G68), .A2(new_n482), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n343), .A2(new_n484), .A3(new_n485), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT81), .B1(new_n490), .B2(KEYINPUT19), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT81), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(new_n487), .C1(new_n461), .C2(new_n343), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n267), .ZN(new_n495));
  INV_X1    g0295(.A(new_n456), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G87), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n474), .A2(G190), .A3(new_n477), .ZN(new_n498));
  AND4_X1   g0298(.A1(new_n481), .A2(new_n495), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G179), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n474), .A2(new_n500), .A3(new_n477), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n480), .B1(new_n494), .B2(new_n267), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT82), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n456), .B2(new_n345), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n267), .B1(new_n310), .B2(G33), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(KEYINPUT82), .A3(new_n264), .A4(new_n344), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n501), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n478), .A2(new_n328), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n479), .A2(new_n499), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n467), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n448), .A2(G169), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n450), .A2(G179), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n469), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n445), .A2(new_n230), .ZN(new_n517));
  OAI211_X1 g0317(.A(G264), .B(G1698), .C1(new_n384), .C2(new_n385), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(KEYINPUT84), .B1(new_n386), .B2(G303), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT84), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n303), .A2(new_n520), .A3(G264), .A4(G1698), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT83), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n429), .B2(new_n232), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n303), .A2(KEYINPUT83), .A3(G257), .A4(new_n305), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n519), .A2(new_n521), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n517), .B1(new_n525), .B2(new_n338), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(G190), .A3(new_n443), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n496), .A2(G116), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n347), .A2(new_n229), .ZN(new_n529));
  AOI21_X1  g0329(.A(G20), .B1(G33), .B2(G283), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n461), .B2(G33), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n266), .A2(new_n237), .B1(G20), .B2(new_n229), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n531), .A2(KEYINPUT20), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT20), .B1(new_n531), .B2(new_n532), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n528), .B(new_n529), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n443), .ZN(new_n537));
  AOI211_X1 g0337(.A(new_n537), .B(new_n517), .C1(new_n525), .C2(new_n338), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n527), .B(new_n536), .C1(new_n319), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(G179), .A3(new_n535), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n535), .A2(G169), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n538), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n526), .A2(new_n443), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n544), .A2(KEYINPUT21), .A3(G169), .A4(new_n535), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n539), .A2(new_n540), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n238), .A2(G107), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n547), .B(KEYINPUT23), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n238), .A2(G33), .A3(G116), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n482), .B2(G87), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n238), .B(G87), .C1(new_n384), .C2(new_n385), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(KEYINPUT22), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n548), .B(new_n549), .C1(new_n551), .C2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n482), .A2(new_n550), .A3(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(KEYINPUT22), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n559), .A2(KEYINPUT24), .A3(new_n548), .A4(new_n549), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n556), .A2(new_n267), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n496), .A2(G107), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OR3_X1    g0363(.A1(new_n264), .A2(KEYINPUT85), .A3(G107), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT85), .B1(new_n264), .B2(G107), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n564), .A2(KEYINPUT25), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT25), .B1(new_n564), .B2(new_n565), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n228), .A2(new_n305), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n232), .A2(G1698), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n570), .C1(new_n384), .C2(new_n385), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G294), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT86), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(KEYINPUT86), .A3(new_n572), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n302), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n443), .B1(new_n577), .B2(KEYINPUT87), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n445), .A2(new_n222), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n571), .A2(KEYINPUT86), .A3(new_n572), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT86), .B1(new_n571), .B2(new_n572), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n338), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT87), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(G169), .B1(new_n578), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n577), .A2(new_n579), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G179), .A3(new_n443), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n563), .A2(new_n568), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n561), .A2(new_n562), .A3(new_n568), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n579), .B1(new_n577), .B2(KEYINPUT87), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n537), .B1(new_n583), .B2(new_n584), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n363), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n583), .A2(new_n443), .A3(new_n580), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n319), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n590), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n546), .A2(new_n589), .A3(new_n596), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n424), .A2(new_n516), .A3(new_n597), .ZN(G372));
  NAND2_X1  g0398(.A1(new_n469), .A2(new_n515), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n328), .B1(new_n591), .B2(new_n592), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n594), .A2(new_n500), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n590), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n603), .A2(new_n540), .A3(new_n543), .A4(new_n545), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n502), .A2(new_n497), .A3(new_n498), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT88), .ZN(new_n606));
  NOR2_X1   g0406(.A1(G238), .A2(G1698), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n276), .B2(new_n277), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(new_n470), .B1(G33), .B2(G116), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n606), .B1(new_n609), .B2(new_n302), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n473), .A2(KEYINPUT88), .A3(new_n338), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n319), .B1(new_n612), .B2(new_n477), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n593), .A2(new_n595), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n561), .A2(new_n562), .A3(new_n568), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n600), .A2(new_n604), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT89), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n450), .A2(new_n328), .ZN(new_n620));
  AOI211_X1 g0420(.A(new_n500), .B(new_n446), .C1(new_n338), .C2(new_n437), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n512), .A2(KEYINPUT89), .A3(new_n513), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n467), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  INV_X1    g0425(.A(new_n614), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n510), .A2(new_n514), .A3(new_n511), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT26), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT88), .B1(new_n473), .B2(new_n338), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n606), .B(new_n302), .C1(new_n471), .C2(new_n472), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n477), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n328), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n508), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n618), .A2(new_n627), .A3(new_n629), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n424), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n413), .ZN(new_n637));
  INV_X1    g0437(.A(new_n353), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n637), .B1(new_n417), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n293), .A2(new_n299), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n272), .A3(new_n321), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n324), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n323), .A2(new_n273), .A3(new_n320), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n335), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n646), .A2(new_n376), .B1(new_n370), .B2(new_n378), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n636), .A2(new_n647), .ZN(G369));
  NOR2_X1   g0448(.A1(new_n589), .A2(new_n596), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n209), .A2(G20), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OR3_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .A3(G1), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT27), .B1(new_n651), .B2(G1), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT90), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n649), .B1(new_n616), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n603), .B2(new_n658), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n543), .A2(new_n545), .A3(new_n540), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n658), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n658), .A2(new_n536), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n661), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n546), .B2(new_n665), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G330), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n649), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n589), .A2(new_n658), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(G399));
  NAND3_X1  g0475(.A1(new_n461), .A2(new_n229), .A3(new_n483), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n676), .B(KEYINPUT91), .Z(new_n677));
  INV_X1    g0477(.A(new_n211), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n242), .B2(new_n680), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  INV_X1    g0484(.A(new_n546), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n516), .A2(new_n649), .A3(new_n685), .A4(new_n658), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT93), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n597), .A2(KEYINPUT93), .A3(new_n516), .A4(new_n658), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n632), .A2(KEYINPUT92), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT92), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n612), .A2(new_n692), .A3(new_n477), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n450), .B1(new_n526), .B2(new_n443), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n500), .A3(new_n594), .A4(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n587), .A2(new_n526), .A3(G179), .A4(new_n443), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n450), .A2(new_n474), .A3(new_n477), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n699), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n602), .A3(KEYINPUT30), .A4(new_n526), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(new_n704), .A3(new_n657), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n704), .B1(new_n703), .B2(new_n657), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n684), .B1(new_n690), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n635), .A2(new_n658), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n617), .B1(new_n589), .B2(new_n661), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n634), .B1(new_n714), .B2(new_n599), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n622), .A2(new_n623), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n511), .A3(new_n626), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT26), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n510), .A2(new_n625), .A3(new_n514), .A4(new_n511), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT29), .B(new_n658), .C1(new_n715), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n710), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n683), .B1(new_n724), .B2(G1), .ZN(G364));
  AOI21_X1  g0525(.A(new_n237), .B1(G20), .B2(new_n328), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n238), .A2(G190), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n500), .A2(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G311), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n238), .A2(new_n363), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n500), .A2(new_n319), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n303), .B(new_n731), .C1(G326), .C2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G322), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(new_n728), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n733), .A2(new_n727), .ZN(new_n739));
  XOR2_X1   g0539(.A(KEYINPUT33), .B(G317), .Z(new_n740));
  OAI221_X1 g0540(.A(new_n736), .B1(new_n737), .B2(new_n738), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n319), .A2(G179), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT96), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n732), .ZN(new_n744));
  INV_X1    g0544(.A(G303), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G179), .A2(G200), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n238), .B1(new_n747), .B2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(G294), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n727), .A2(new_n747), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G329), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n743), .A2(new_n727), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n753), .B1(new_n755), .B2(new_n425), .ZN(new_n756));
  NOR4_X1   g0556(.A1(new_n741), .A2(new_n746), .A3(new_n750), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n754), .A2(G107), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n758), .B1(new_n403), .B2(new_n734), .C1(new_n227), .C2(new_n744), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n303), .B1(new_n739), .B2(new_n294), .ZN(new_n760));
  INV_X1    g0560(.A(new_n748), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(G97), .B2(new_n761), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n762), .B1(new_n220), .B2(new_n738), .C1(new_n217), .C2(new_n729), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n752), .A2(G159), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT32), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n759), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n726), .B1(new_n757), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n310), .B1(new_n650), .B2(G45), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n679), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n211), .A2(G355), .A3(new_n303), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n256), .A2(new_n439), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n678), .A2(new_n303), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G45), .B2(new_n242), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n772), .B1(G116), .B2(new_n211), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n726), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT94), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n771), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT95), .ZN(new_n784));
  INV_X1    g0584(.A(new_n779), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n767), .B(new_n784), .C1(new_n667), .C2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT97), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n669), .A2(new_n770), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(G330), .B2(new_n667), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n789), .ZN(G396));
  NOR2_X1   g0590(.A1(new_n744), .A2(new_n403), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n755), .A2(new_n294), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n729), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G137), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n734), .A2(new_n796), .B1(new_n739), .B2(new_n366), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT98), .Z(new_n798));
  INV_X1    g0598(.A(new_n738), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n795), .B(new_n798), .C1(G143), .C2(new_n799), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n303), .B(new_n793), .C1(new_n800), .C2(KEYINPUT34), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n791), .B(new_n801), .C1(KEYINPUT34), .C2(new_n800), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n802), .B1(new_n220), .B2(new_n748), .C1(new_n803), .C2(new_n751), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n755), .A2(new_n227), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n739), .A2(new_n425), .B1(new_n748), .B2(new_n202), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n744), .A2(new_n203), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n734), .A2(new_n745), .B1(new_n738), .B2(new_n749), .ZN(new_n808));
  NOR4_X1   g0608(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n809), .A2(new_n386), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n810), .B1(new_n229), .B2(new_n729), .C1(new_n730), .C2(new_n751), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n804), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n771), .B1(new_n812), .B2(new_n726), .ZN(new_n813));
  INV_X1    g0613(.A(new_n726), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n778), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n353), .A2(new_n657), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n657), .A2(new_n351), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n422), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(new_n818), .B2(new_n353), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n813), .B1(G77), .B2(new_n815), .C1(new_n778), .C2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n819), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n711), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n635), .A2(new_n658), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n710), .B(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n820), .B1(new_n825), .B2(new_n770), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT99), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G384));
  INV_X1    g0628(.A(new_n288), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n292), .B1(new_n295), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n297), .A2(new_n267), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n272), .ZN(new_n832));
  INV_X1    g0632(.A(new_n655), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n331), .A2(new_n334), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n645), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n330), .A2(new_n655), .B1(new_n272), .B2(new_n831), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT37), .B1(new_n643), .B2(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n323), .A2(new_n273), .B1(new_n333), .B2(new_n833), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n641), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n837), .A2(KEYINPUT38), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n834), .B1(new_n326), .B2(new_n335), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n839), .A2(new_n842), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n844), .A2(new_n848), .A3(KEYINPUT39), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n300), .A2(new_n655), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n326), .B2(new_n335), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n641), .A2(new_n840), .A3(new_n841), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n841), .B1(new_n641), .B2(new_n840), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n845), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT39), .B1(new_n844), .B2(new_n856), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n849), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n413), .A2(new_n657), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT101), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n837), .B2(new_n843), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n846), .A2(new_n847), .A3(new_n845), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n657), .A2(new_n412), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n866), .B(new_n416), .C1(new_n402), .C2(new_n412), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n413), .A2(new_n658), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n816), .B(KEYINPUT100), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n823), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n844), .A2(new_n848), .A3(KEYINPUT101), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n865), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n335), .B2(new_n833), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n861), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n424), .A2(new_n713), .A3(new_n721), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n647), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n875), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n819), .B1(new_n867), .B2(new_n868), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n690), .B2(new_n708), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n865), .A2(new_n872), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n844), .B2(new_n856), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n880), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(G330), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n424), .A2(new_n709), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n881), .A2(new_n882), .B1(new_n884), .B2(new_n880), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n707), .B1(new_n688), .B2(new_n689), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n889), .A2(new_n424), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n878), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n310), .B2(new_n650), .ZN(new_n895));
  INV_X1    g0695(.A(new_n465), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n229), .B1(new_n896), .B2(KEYINPUT35), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(new_n239), .C1(KEYINPUT35), .C2(new_n896), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT36), .ZN(new_n899));
  OAI21_X1  g0699(.A(G77), .B1(new_n220), .B2(new_n294), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n242), .A2(new_n900), .B1(G50), .B2(new_n294), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(G1), .A3(new_n209), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n895), .A2(new_n899), .A3(new_n902), .ZN(G367));
  NAND3_X1  g0703(.A1(new_n663), .A2(new_n600), .A3(new_n649), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n600), .B1(new_n467), .B2(new_n658), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n624), .A2(new_n657), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n908), .A2(new_n589), .B1(new_n514), .B2(new_n511), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n905), .B1(new_n909), .B2(new_n657), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n910), .A2(KEYINPUT102), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(KEYINPUT102), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n502), .A2(new_n497), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n657), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n626), .A2(new_n916), .A3(new_n634), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n634), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT103), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n914), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n908), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n670), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n926), .A2(new_n673), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT45), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT44), .B1(new_n674), .B2(new_n908), .ZN(new_n932));
  OR3_X1    g0732(.A1(new_n674), .A2(KEYINPUT44), .A3(new_n908), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(new_n670), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n664), .A2(new_n671), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT104), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n668), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n670), .B(KEYINPUT105), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n723), .B1(new_n935), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n679), .B(KEYINPUT41), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n768), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n922), .A2(new_n927), .A3(new_n924), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n929), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n739), .ZN(new_n949));
  AOI22_X1  g0749(.A1(G294), .A2(new_n949), .B1(new_n752), .B2(G317), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT106), .B1(new_n744), .B2(new_n229), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(KEYINPUT46), .ZN(new_n952));
  INV_X1    g0752(.A(new_n729), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n303), .B1(new_n953), .B2(G283), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n735), .A2(G311), .B1(new_n761), .B2(G107), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(new_n755), .C2(new_n461), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n952), .B(new_n956), .C1(G303), .C2(new_n799), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n951), .A2(KEYINPUT46), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n744), .A2(new_n220), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n754), .A2(G77), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n761), .A2(G68), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n735), .A2(G143), .B1(new_n752), .B2(G137), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n386), .B1(new_n953), .B2(G50), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n960), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n959), .B(new_n964), .C1(G150), .C2(new_n799), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n949), .A2(G159), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n957), .A2(new_n958), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT47), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n726), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n918), .A2(new_n785), .ZN(new_n970));
  INV_X1    g0770(.A(new_n774), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n782), .B1(new_n211), .B2(new_n345), .C1(new_n252), .C2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n969), .A2(new_n970), .A3(new_n770), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n948), .A2(new_n973), .ZN(G387));
  NAND2_X1  g0774(.A1(new_n942), .A2(new_n724), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n680), .B1(new_n941), .B2(new_n723), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n774), .B1(new_n248), .B2(new_n439), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n211), .A2(new_n303), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n978), .B1(new_n677), .B2(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n677), .B(new_n439), .C1(new_n294), .C2(new_n217), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n262), .A2(new_n403), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT50), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n980), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n678), .A2(new_n203), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n781), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n739), .A2(new_n261), .B1(new_n729), .B2(new_n294), .ZN(new_n987));
  INV_X1    g0787(.A(new_n744), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n988), .A2(G77), .B1(G150), .B2(new_n752), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n989), .B(new_n303), .C1(new_n202), .C2(new_n755), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT107), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n987), .B(new_n991), .C1(G159), .C2(new_n735), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n761), .A2(new_n344), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n403), .C2(new_n738), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT108), .Z(new_n995));
  AOI21_X1  g0795(.A(new_n303), .B1(new_n752), .B2(G326), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n755), .B2(new_n229), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G311), .A2(new_n949), .B1(new_n799), .B2(G317), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n745), .B2(new_n729), .C1(new_n737), .C2(new_n734), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n425), .B2(new_n748), .C1(new_n749), .C2(new_n744), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT49), .Z(new_n1002));
  OAI21_X1  g0802(.A(new_n995), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n771), .B(new_n986), .C1(new_n1003), .C2(new_n726), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n660), .A2(new_n785), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n942), .A2(new_n769), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n977), .A2(new_n1006), .ZN(G393));
  INV_X1    g0807(.A(KEYINPUT109), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n935), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n934), .A2(KEYINPUT109), .A3(new_n669), .A4(new_n664), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1009), .A2(new_n975), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT111), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n975), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1011), .A2(new_n1012), .B1(new_n1013), .B2(new_n935), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n679), .C1(new_n1012), .C2(new_n1011), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n769), .ZN(new_n1017));
  INV_X1    g0817(.A(G317), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n734), .A2(new_n1018), .B1(new_n738), .B2(new_n730), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT52), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n1021), .A2(new_n1022), .A3(new_n303), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n758), .B1(new_n229), .B2(new_n748), .C1(new_n425), .C2(new_n744), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(G294), .C2(new_n953), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n745), .B2(new_n739), .C1(new_n737), .C2(new_n751), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n734), .A2(new_n366), .B1(new_n738), .B2(new_n794), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT51), .Z(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(new_n805), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n752), .A2(G143), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n739), .A2(new_n403), .B1(new_n729), .B2(new_n261), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT110), .Z(new_n1032));
  OAI21_X1  g0832(.A(new_n303), .B1(new_n744), .B2(new_n294), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G77), .B2(new_n761), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n814), .B1(new_n1026), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n211), .A2(new_n461), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1037), .B(new_n781), .C1(new_n259), .C2(new_n774), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1036), .A2(new_n771), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n908), .B2(new_n785), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1015), .A2(new_n1017), .A3(new_n1040), .ZN(G390));
  OAI22_X1  g0841(.A1(new_n849), .A2(new_n857), .B1(new_n871), .B2(new_n859), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n850), .B1(new_n836), .B2(new_n645), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n853), .A2(new_n854), .ZN(new_n1044));
  AOI21_X1  g0844(.A(KEYINPUT38), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n860), .B1(new_n1045), .B2(new_n864), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT112), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n818), .A2(new_n353), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n658), .B(new_n1048), .C1(new_n715), .C2(new_n720), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n816), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n869), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1046), .A2(new_n1047), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n869), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n859), .B1(new_n844), .B2(new_n856), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT112), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1042), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(KEYINPUT113), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n890), .A2(new_n684), .A3(new_n821), .A4(new_n869), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT113), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1042), .B(new_n1061), .C1(new_n1052), .C2(new_n1057), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1060), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1058), .A2(KEYINPUT113), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n823), .A2(new_n870), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1054), .B1(new_n709), .B2(new_n819), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n1060), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(KEYINPUT114), .ZN(new_n1070));
  OR3_X1    g0870(.A1(new_n1068), .A2(new_n1060), .A3(new_n1053), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT114), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1072), .B(new_n1067), .C1(new_n1068), .C2(new_n1060), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n876), .A2(new_n887), .A3(new_n647), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1066), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(new_n1065), .A3(new_n1063), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n679), .A3(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n988), .A2(G87), .B1(G283), .B2(new_n735), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G294), .A2(new_n752), .B1(new_n761), .B2(G77), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n793), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n386), .B1(new_n739), .B2(new_n203), .C1(new_n229), .C2(new_n738), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n729), .A2(new_n461), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT115), .Z(new_n1088));
  XOR2_X1   g0888(.A(KEYINPUT54), .B(G143), .Z(new_n1089));
  AOI22_X1  g0889(.A1(G128), .A2(new_n735), .B1(new_n953), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n794), .B2(new_n748), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n386), .B(new_n1091), .C1(G50), .C2(new_n754), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n949), .A2(G137), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n752), .A2(G125), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n744), .A2(new_n366), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT53), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G132), .B2(new_n799), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n726), .B1(new_n1088), .B2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1099), .B(new_n770), .C1(new_n262), .C2(new_n815), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n858), .B2(new_n777), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1066), .B2(new_n769), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1081), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT116), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1081), .A2(new_n1105), .A3(new_n1102), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(G378));
  INV_X1    g0907(.A(KEYINPUT57), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n886), .A2(KEYINPUT118), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT118), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n883), .A2(new_n1110), .A3(G330), .A4(new_n885), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1112));
  XOR2_X1   g0912(.A(new_n380), .B(new_n1112), .Z(new_n1113));
  NAND2_X1  g0913(.A1(new_n833), .A2(new_n370), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1113), .B(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1109), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n875), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1113), .B(new_n1114), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n886), .A2(new_n1119), .A3(KEYINPUT118), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1118), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1075), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1108), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1108), .B1(new_n1078), .B2(new_n1076), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT119), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1110), .B1(new_n889), .B2(G330), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1120), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n875), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(KEYINPUT119), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1126), .A2(new_n1128), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1125), .A2(new_n1136), .A3(new_n679), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n769), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n754), .A2(G58), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1140), .B(new_n961), .C1(new_n217), .C2(new_n744), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n734), .A2(new_n229), .B1(new_n751), .B2(new_n425), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n301), .B(new_n386), .C1(new_n739), .C2(new_n202), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n203), .B2(new_n738), .C1(new_n345), .C2(new_n729), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT117), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT58), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n403), .B1(new_n384), .B2(G41), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n988), .A2(new_n1089), .B1(G137), .B2(new_n953), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n735), .A2(G125), .B1(new_n761), .B2(G150), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(G128), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1151), .B1(new_n1152), .B2(new_n738), .C1(new_n803), .C2(new_n739), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G41), .B1(new_n1153), .B2(KEYINPUT59), .ZN(new_n1155));
  AOI21_X1  g0955(.A(G33), .B1(new_n752), .B2(G124), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n794), .C2(new_n755), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1147), .B(new_n1148), .C1(new_n1154), .C2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n771), .B1(new_n1158), .B2(new_n726), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(G50), .B2(new_n815), .C1(new_n1119), .C2(new_n778), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1139), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1137), .A2(new_n1161), .ZN(G375));
  NAND2_X1  g0962(.A1(new_n1074), .A2(new_n769), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT121), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1140), .B1(new_n403), .B2(new_n748), .C1(new_n803), .C2(new_n734), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G159), .B2(new_n988), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n386), .B1(new_n953), .B2(G150), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(new_n796), .C2(new_n738), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n949), .B2(new_n1089), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n751), .A2(new_n1152), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n949), .A2(G116), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n303), .B1(new_n953), .B2(G107), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1174), .B(new_n993), .C1(new_n749), .C2(new_n734), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n960), .B1(new_n425), .B2(new_n738), .C1(new_n745), .C2(new_n751), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(G97), .C2(new_n988), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1170), .A2(new_n1172), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n770), .B1(G68), .B2(new_n815), .C1(new_n1178), .C2(new_n814), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n869), .B2(new_n777), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1165), .A2(new_n1181), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1183), .A2(KEYINPUT120), .A3(new_n1075), .A4(new_n1071), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1070), .A2(new_n1071), .A3(new_n1075), .A4(new_n1073), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT120), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1188), .A2(new_n1077), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1182), .B1(new_n1189), .B2(new_n945), .ZN(G381));
  NOR2_X1   g0990(.A1(G375), .A2(new_n1103), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(G381), .A2(G387), .A3(G384), .ZN(new_n1192));
  INV_X1    g0992(.A(G390), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(G393), .A2(G396), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(G407));
  NAND2_X1  g0995(.A1(new_n656), .A2(G213), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT122), .Z(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1191), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(G407), .A2(G213), .A3(new_n1199), .ZN(G409));
  INV_X1    g1000(.A(KEYINPUT125), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1196), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1184), .A2(new_n1187), .B1(KEYINPUT60), .B2(new_n1079), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1185), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT60), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1203), .A2(new_n680), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1165), .A2(new_n1181), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n827), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1079), .A2(KEYINPUT60), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n679), .B(new_n1205), .C1(new_n1188), .C2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1182), .A2(new_n1211), .A3(G384), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(G378), .A2(new_n1137), .A3(new_n1161), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1135), .A2(new_n769), .A3(new_n1128), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1124), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n944), .A3(new_n1138), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1217), .A3(new_n1160), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n1102), .A3(new_n1081), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1202), .B(new_n1213), .C1(new_n1214), .C2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1201), .B1(new_n1220), .B2(KEYINPUT62), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1214), .A2(new_n1219), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1213), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1196), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(KEYINPUT125), .A3(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1222), .A2(KEYINPUT62), .A3(new_n1197), .A4(new_n1223), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1221), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1213), .B1(G2897), .B2(new_n1202), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1198), .A2(G2897), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT123), .B1(new_n1223), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT123), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1213), .A2(new_n1232), .A3(G2897), .A4(new_n1198), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1229), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1222), .A2(new_n1197), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT61), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1228), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT124), .B1(new_n948), .B2(new_n973), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(G393), .B(G396), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1239), .B1(new_n973), .B2(new_n948), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1193), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(G387), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(G390), .C1(new_n1240), .C2(new_n1238), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1237), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT63), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1235), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT61), .B1(new_n1250), .B2(new_n1223), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1222), .A2(new_n1196), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1249), .B1(new_n1234), .B2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1251), .B(new_n1246), .C1(new_n1253), .C2(new_n1220), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1248), .A2(new_n1254), .ZN(G405));
  NOR2_X1   g1055(.A1(new_n1213), .A2(KEYINPUT127), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1246), .B(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1103), .B1(new_n1137), .B2(new_n1161), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT126), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1260), .A2(new_n1214), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1261), .A2(new_n1262), .B1(KEYINPUT127), .B2(new_n1213), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1257), .B(new_n1263), .Z(G402));
endmodule


