

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(G2105), .ZN(n528) );
  XOR2_X1 U555 ( .A(KEYINPUT1), .B(n533), .Z(n793) );
  NOR2_X2 U556 ( .A1(n677), .A2(n676), .ZN(n678) );
  OR2_X1 U557 ( .A1(n694), .A2(n693), .ZN(n695) );
  OR2_X1 U558 ( .A1(n644), .A2(n643), .ZN(n647) );
  XNOR2_X1 U559 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n616) );
  XNOR2_X1 U560 ( .A(n617), .B(n616), .ZN(n664) );
  NAND2_X1 U561 ( .A1(G8), .A2(n640), .ZN(n702) );
  AND2_X2 U562 ( .A1(n528), .A2(G2104), .ZN(n883) );
  NOR2_X1 U563 ( .A1(n577), .A2(G651), .ZN(n795) );
  NOR2_X2 U564 ( .A1(n532), .A2(n531), .ZN(G160) );
  XNOR2_X1 U565 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n524) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XNOR2_X2 U567 ( .A(n524), .B(n523), .ZN(n884) );
  NAND2_X1 U568 ( .A1(n884), .A2(G137), .ZN(n527) );
  NAND2_X1 U569 ( .A1(G101), .A2(n883), .ZN(n525) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n525), .Z(n526) );
  NAND2_X1 U571 ( .A1(n527), .A2(n526), .ZN(n532) );
  NOR2_X4 U572 ( .A1(G2104), .A2(n528), .ZN(n888) );
  NAND2_X1 U573 ( .A1(G125), .A2(n888), .ZN(n530) );
  AND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U575 ( .A1(G113), .A2(n889), .ZN(n529) );
  NAND2_X1 U576 ( .A1(n530), .A2(n529), .ZN(n531) );
  INV_X1 U577 ( .A(G651), .ZN(n539) );
  NOR2_X1 U578 ( .A1(G543), .A2(n539), .ZN(n533) );
  NAND2_X1 U579 ( .A1(G63), .A2(n793), .ZN(n535) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n577) );
  NAND2_X1 U581 ( .A1(G51), .A2(n795), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U583 ( .A(KEYINPUT6), .B(n536), .ZN(n544) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n537) );
  XNOR2_X1 U585 ( .A(n537), .B(KEYINPUT64), .ZN(n790) );
  NAND2_X1 U586 ( .A1(G89), .A2(n790), .ZN(n538) );
  XNOR2_X1 U587 ( .A(n538), .B(KEYINPUT4), .ZN(n541) );
  NOR2_X1 U588 ( .A1(n577), .A2(n539), .ZN(n789) );
  NAND2_X1 U589 ( .A1(G76), .A2(n789), .ZN(n540) );
  NAND2_X1 U590 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U591 ( .A(n542), .B(KEYINPUT5), .Z(n543) );
  NOR2_X1 U592 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U593 ( .A(KEYINPUT7), .B(n545), .Z(n546) );
  XNOR2_X1 U594 ( .A(KEYINPUT76), .B(n546), .ZN(G168) );
  XOR2_X1 U595 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U596 ( .A1(G64), .A2(n793), .ZN(n548) );
  NAND2_X1 U597 ( .A1(G52), .A2(n795), .ZN(n547) );
  NAND2_X1 U598 ( .A1(n548), .A2(n547), .ZN(n553) );
  NAND2_X1 U599 ( .A1(n789), .A2(G77), .ZN(n550) );
  NAND2_X1 U600 ( .A1(G90), .A2(n790), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U602 ( .A(KEYINPUT9), .B(n551), .Z(n552) );
  NOR2_X1 U603 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U604 ( .A(KEYINPUT67), .B(n554), .ZN(G301) );
  NAND2_X1 U605 ( .A1(n789), .A2(G78), .ZN(n556) );
  NAND2_X1 U606 ( .A1(G91), .A2(n790), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U608 ( .A(KEYINPUT68), .B(n557), .Z(n563) );
  NAND2_X1 U609 ( .A1(n795), .A2(G53), .ZN(n558) );
  XOR2_X1 U610 ( .A(KEYINPUT69), .B(n558), .Z(n560) );
  NAND2_X1 U611 ( .A1(n793), .A2(G65), .ZN(n559) );
  NAND2_X1 U612 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U613 ( .A(KEYINPUT70), .B(n561), .Z(n562) );
  NAND2_X1 U614 ( .A1(n563), .A2(n562), .ZN(G299) );
  NAND2_X1 U615 ( .A1(G62), .A2(n793), .ZN(n564) );
  XNOR2_X1 U616 ( .A(n564), .B(KEYINPUT82), .ZN(n571) );
  NAND2_X1 U617 ( .A1(G75), .A2(n789), .ZN(n566) );
  NAND2_X1 U618 ( .A1(G50), .A2(n795), .ZN(n565) );
  NAND2_X1 U619 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U620 ( .A1(G88), .A2(n790), .ZN(n567) );
  XNOR2_X1 U621 ( .A(KEYINPUT83), .B(n567), .ZN(n568) );
  NOR2_X1 U622 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U623 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U624 ( .A(KEYINPUT84), .B(n572), .Z(G166) );
  XOR2_X1 U625 ( .A(KEYINPUT92), .B(G166), .Z(G303) );
  NAND2_X1 U626 ( .A1(G49), .A2(n795), .ZN(n574) );
  NAND2_X1 U627 ( .A1(G74), .A2(G651), .ZN(n573) );
  NAND2_X1 U628 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U629 ( .A(KEYINPUT80), .B(n575), .ZN(n576) );
  NOR2_X1 U630 ( .A1(n793), .A2(n576), .ZN(n579) );
  NAND2_X1 U631 ( .A1(n577), .A2(G87), .ZN(n578) );
  NAND2_X1 U632 ( .A1(n579), .A2(n578), .ZN(G288) );
  NAND2_X1 U633 ( .A1(n793), .A2(G61), .ZN(n581) );
  NAND2_X1 U634 ( .A1(G86), .A2(n790), .ZN(n580) );
  NAND2_X1 U635 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U636 ( .A1(G73), .A2(n789), .ZN(n582) );
  XNOR2_X1 U637 ( .A(n582), .B(KEYINPUT81), .ZN(n583) );
  XNOR2_X1 U638 ( .A(n583), .B(KEYINPUT2), .ZN(n584) );
  NOR2_X1 U639 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U640 ( .A1(n795), .A2(G48), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n587), .A2(n586), .ZN(G305) );
  INV_X1 U642 ( .A(KEYINPUT89), .ZN(n589) );
  NAND2_X1 U643 ( .A1(n888), .A2(G126), .ZN(n588) );
  XNOR2_X1 U644 ( .A(n589), .B(n588), .ZN(n591) );
  NAND2_X1 U645 ( .A1(n889), .A2(G114), .ZN(n590) );
  NAND2_X1 U646 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U647 ( .A(KEYINPUT90), .B(n592), .Z(n594) );
  NAND2_X1 U648 ( .A1(n884), .A2(G138), .ZN(n593) );
  NAND2_X1 U649 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U650 ( .A1(G102), .A2(n883), .ZN(n595) );
  XNOR2_X1 U651 ( .A(KEYINPUT91), .B(n595), .ZN(n596) );
  NOR2_X1 U652 ( .A1(n597), .A2(n596), .ZN(n607) );
  BUF_X1 U653 ( .A(n607), .Z(G164) );
  NAND2_X1 U654 ( .A1(n789), .A2(G72), .ZN(n599) );
  NAND2_X1 U655 ( .A1(G85), .A2(n790), .ZN(n598) );
  NAND2_X1 U656 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U657 ( .A1(G47), .A2(n795), .ZN(n600) );
  XOR2_X1 U658 ( .A(KEYINPUT66), .B(n600), .Z(n601) );
  NOR2_X1 U659 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U660 ( .A1(n793), .A2(G60), .ZN(n603) );
  NAND2_X1 U661 ( .A1(n604), .A2(n603), .ZN(G290) );
  XOR2_X1 U662 ( .A(G2078), .B(KEYINPUT25), .Z(n948) );
  NAND2_X1 U663 ( .A1(G160), .A2(G40), .ZN(n707) );
  INV_X1 U664 ( .A(n707), .ZN(n606) );
  INV_X1 U665 ( .A(G1384), .ZN(n605) );
  NAND2_X1 U666 ( .A1(n606), .A2(n605), .ZN(n608) );
  OR2_X2 U667 ( .A1(n608), .A2(n607), .ZN(n640) );
  INV_X2 U668 ( .A(n640), .ZN(n649) );
  INV_X1 U669 ( .A(n649), .ZN(n667) );
  NOR2_X1 U670 ( .A1(n948), .A2(n667), .ZN(n610) );
  NOR2_X1 U671 ( .A1(n649), .A2(G1961), .ZN(n609) );
  NOR2_X1 U672 ( .A1(n610), .A2(n609), .ZN(n660) );
  AND2_X1 U673 ( .A1(G301), .A2(n660), .ZN(n615) );
  NOR2_X1 U674 ( .A1(G2084), .A2(n667), .ZN(n679) );
  NOR2_X1 U675 ( .A1(G1966), .A2(n702), .ZN(n677) );
  NOR2_X1 U676 ( .A1(n679), .A2(n677), .ZN(n611) );
  NAND2_X1 U677 ( .A1(G8), .A2(n611), .ZN(n612) );
  XNOR2_X1 U678 ( .A(KEYINPUT30), .B(n612), .ZN(n613) );
  NOR2_X1 U679 ( .A1(n613), .A2(G168), .ZN(n614) );
  NOR2_X1 U680 ( .A1(n615), .A2(n614), .ZN(n617) );
  XOR2_X1 U681 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n619) );
  NAND2_X1 U682 ( .A1(G56), .A2(n793), .ZN(n618) );
  XNOR2_X1 U683 ( .A(n619), .B(n618), .ZN(n625) );
  NAND2_X1 U684 ( .A1(G81), .A2(n790), .ZN(n620) );
  XNOR2_X1 U685 ( .A(n620), .B(KEYINPUT12), .ZN(n622) );
  NAND2_X1 U686 ( .A1(G68), .A2(n789), .ZN(n621) );
  NAND2_X1 U687 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U688 ( .A(KEYINPUT13), .B(n623), .Z(n624) );
  NOR2_X1 U689 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U690 ( .A1(n795), .A2(G43), .ZN(n626) );
  NAND2_X1 U691 ( .A1(n627), .A2(n626), .ZN(n992) );
  INV_X1 U692 ( .A(G1996), .ZN(n947) );
  NOR2_X1 U693 ( .A1(n640), .A2(n947), .ZN(n628) );
  XOR2_X1 U694 ( .A(n628), .B(KEYINPUT26), .Z(n630) );
  NAND2_X1 U695 ( .A1(n667), .A2(G1341), .ZN(n629) );
  NAND2_X1 U696 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U697 ( .A1(n992), .A2(n631), .ZN(n644) );
  NAND2_X1 U698 ( .A1(n793), .A2(G66), .ZN(n633) );
  NAND2_X1 U699 ( .A1(G92), .A2(n790), .ZN(n632) );
  NAND2_X1 U700 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U701 ( .A1(G79), .A2(n789), .ZN(n635) );
  NAND2_X1 U702 ( .A1(G54), .A2(n795), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U705 ( .A(KEYINPUT15), .B(n638), .Z(n639) );
  XNOR2_X2 U706 ( .A(KEYINPUT73), .B(n639), .ZN(n977) );
  NAND2_X1 U707 ( .A1(G1348), .A2(n640), .ZN(n642) );
  NAND2_X1 U708 ( .A1(n649), .A2(G2067), .ZN(n641) );
  NAND2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n645) );
  NOR2_X1 U710 ( .A1(n977), .A2(n645), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n977), .A2(n645), .ZN(n646) );
  NAND2_X1 U712 ( .A1(n647), .A2(n646), .ZN(n653) );
  INV_X1 U713 ( .A(G299), .ZN(n975) );
  NAND2_X1 U714 ( .A1(n649), .A2(G2072), .ZN(n648) );
  XNOR2_X1 U715 ( .A(n648), .B(KEYINPUT27), .ZN(n651) );
  XNOR2_X1 U716 ( .A(G1956), .B(KEYINPUT97), .ZN(n1011) );
  NOR2_X1 U717 ( .A1(n1011), .A2(n649), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n975), .A2(n654), .ZN(n652) );
  NAND2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n658) );
  NOR2_X1 U721 ( .A1(n654), .A2(n975), .ZN(n655) );
  XNOR2_X1 U722 ( .A(n655), .B(KEYINPUT28), .ZN(n656) );
  INV_X1 U723 ( .A(n656), .ZN(n657) );
  NAND2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U725 ( .A(n659), .B(KEYINPUT29), .ZN(n662) );
  NOR2_X1 U726 ( .A1(G301), .A2(n660), .ZN(n661) );
  NOR2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U728 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U729 ( .A(n665), .B(KEYINPUT99), .ZN(n675) );
  NAND2_X1 U730 ( .A1(G286), .A2(n675), .ZN(n672) );
  NOR2_X1 U731 ( .A1(G1971), .A2(n702), .ZN(n666) );
  XOR2_X1 U732 ( .A(KEYINPUT101), .B(n666), .Z(n669) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n667), .ZN(n668) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U735 ( .A1(n670), .A2(G303), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U737 ( .A1(G8), .A2(n673), .ZN(n674) );
  XNOR2_X1 U738 ( .A(n674), .B(KEYINPUT32), .ZN(n683) );
  INV_X1 U739 ( .A(n675), .ZN(n676) );
  XNOR2_X1 U740 ( .A(n678), .B(KEYINPUT100), .ZN(n681) );
  NAND2_X1 U741 ( .A1(n679), .A2(G8), .ZN(n680) );
  NAND2_X1 U742 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n696) );
  NOR2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n983) );
  NOR2_X1 U745 ( .A1(G1971), .A2(G303), .ZN(n684) );
  NOR2_X1 U746 ( .A1(n983), .A2(n684), .ZN(n685) );
  NAND2_X1 U747 ( .A1(n696), .A2(n685), .ZN(n687) );
  NAND2_X1 U748 ( .A1(G288), .A2(G1976), .ZN(n686) );
  XNOR2_X1 U749 ( .A(n686), .B(KEYINPUT102), .ZN(n981) );
  NAND2_X1 U750 ( .A1(n687), .A2(n981), .ZN(n690) );
  NAND2_X1 U751 ( .A1(n983), .A2(KEYINPUT33), .ZN(n688) );
  NOR2_X1 U752 ( .A1(n688), .A2(n702), .ZN(n691) );
  OR2_X1 U753 ( .A1(n702), .A2(n691), .ZN(n689) );
  NOR2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n694) );
  INV_X1 U755 ( .A(n691), .ZN(n692) );
  AND2_X1 U756 ( .A1(n692), .A2(KEYINPUT33), .ZN(n693) );
  XOR2_X1 U757 ( .A(G1981), .B(G305), .Z(n972) );
  NAND2_X1 U758 ( .A1(n695), .A2(n972), .ZN(n706) );
  NOR2_X1 U759 ( .A1(G2090), .A2(G303), .ZN(n697) );
  NAND2_X1 U760 ( .A1(G8), .A2(n697), .ZN(n698) );
  NAND2_X1 U761 ( .A1(n696), .A2(n698), .ZN(n699) );
  AND2_X1 U762 ( .A1(n699), .A2(n702), .ZN(n704) );
  NOR2_X1 U763 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XOR2_X1 U764 ( .A(n700), .B(KEYINPUT24), .Z(n701) );
  NOR2_X1 U765 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U766 ( .A1(n704), .A2(n703), .ZN(n705) );
  AND2_X1 U767 ( .A1(n706), .A2(n705), .ZN(n740) );
  NOR2_X1 U768 ( .A1(G164), .A2(G1384), .ZN(n708) );
  NOR2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n756) );
  NAND2_X1 U770 ( .A1(G128), .A2(n888), .ZN(n710) );
  NAND2_X1 U771 ( .A1(G116), .A2(n889), .ZN(n709) );
  NAND2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U773 ( .A(n711), .B(KEYINPUT35), .ZN(n716) );
  NAND2_X1 U774 ( .A1(G104), .A2(n883), .ZN(n713) );
  NAND2_X1 U775 ( .A1(G140), .A2(n884), .ZN(n712) );
  NAND2_X1 U776 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U777 ( .A(KEYINPUT34), .B(n714), .Z(n715) );
  NAND2_X1 U778 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U779 ( .A(n717), .B(KEYINPUT36), .ZN(n874) );
  XOR2_X1 U780 ( .A(G2067), .B(KEYINPUT37), .Z(n752) );
  NAND2_X1 U781 ( .A1(n874), .A2(n752), .ZN(n718) );
  XNOR2_X1 U782 ( .A(n718), .B(KEYINPUT93), .ZN(n938) );
  NAND2_X1 U783 ( .A1(n756), .A2(n938), .ZN(n750) );
  INV_X1 U784 ( .A(n750), .ZN(n738) );
  NAND2_X1 U785 ( .A1(G107), .A2(n889), .ZN(n719) );
  XNOR2_X1 U786 ( .A(n719), .B(KEYINPUT94), .ZN(n722) );
  NAND2_X1 U787 ( .A1(G95), .A2(n883), .ZN(n720) );
  XOR2_X1 U788 ( .A(KEYINPUT95), .B(n720), .Z(n721) );
  NAND2_X1 U789 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U790 ( .A1(G119), .A2(n888), .ZN(n724) );
  NAND2_X1 U791 ( .A1(G131), .A2(n884), .ZN(n723) );
  NAND2_X1 U792 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U793 ( .A1(n726), .A2(n725), .ZN(n873) );
  INV_X1 U794 ( .A(G1991), .ZN(n945) );
  NOR2_X1 U795 ( .A1(n873), .A2(n945), .ZN(n735) );
  NAND2_X1 U796 ( .A1(G117), .A2(n889), .ZN(n728) );
  NAND2_X1 U797 ( .A1(G141), .A2(n884), .ZN(n727) );
  NAND2_X1 U798 ( .A1(n728), .A2(n727), .ZN(n731) );
  NAND2_X1 U799 ( .A1(n883), .A2(G105), .ZN(n729) );
  XOR2_X1 U800 ( .A(KEYINPUT38), .B(n729), .Z(n730) );
  NOR2_X1 U801 ( .A1(n731), .A2(n730), .ZN(n733) );
  NAND2_X1 U802 ( .A1(n888), .A2(G129), .ZN(n732) );
  NAND2_X1 U803 ( .A1(n733), .A2(n732), .ZN(n872) );
  AND2_X1 U804 ( .A1(G1996), .A2(n872), .ZN(n734) );
  NOR2_X1 U805 ( .A1(n735), .A2(n734), .ZN(n929) );
  INV_X1 U806 ( .A(n756), .ZN(n736) );
  NOR2_X1 U807 ( .A1(n929), .A2(n736), .ZN(n746) );
  XNOR2_X1 U808 ( .A(KEYINPUT96), .B(n746), .ZN(n737) );
  OR2_X1 U809 ( .A1(n738), .A2(n737), .ZN(n739) );
  OR2_X1 U810 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U811 ( .A(n741), .B(KEYINPUT103), .ZN(n743) );
  XNOR2_X1 U812 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U813 ( .A1(n756), .A2(n979), .ZN(n742) );
  NAND2_X1 U814 ( .A1(n743), .A2(n742), .ZN(n759) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n872), .ZN(n931) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n744) );
  AND2_X1 U817 ( .A1(n945), .A2(n873), .ZN(n927) );
  NOR2_X1 U818 ( .A1(n744), .A2(n927), .ZN(n745) );
  NOR2_X1 U819 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U820 ( .A(n747), .B(KEYINPUT104), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n931), .A2(n748), .ZN(n749) );
  XNOR2_X1 U822 ( .A(n749), .B(KEYINPUT39), .ZN(n751) );
  NAND2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n754) );
  NOR2_X1 U824 ( .A1(n874), .A2(n752), .ZN(n753) );
  XNOR2_X1 U825 ( .A(n753), .B(KEYINPUT105), .ZN(n924) );
  NAND2_X1 U826 ( .A1(n754), .A2(n924), .ZN(n755) );
  NAND2_X1 U827 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U828 ( .A(n757), .B(KEYINPUT106), .ZN(n758) );
  NAND2_X1 U829 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U830 ( .A(n760), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U831 ( .A(G301), .ZN(G171) );
  AND2_X1 U832 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U833 ( .A1(G135), .A2(n884), .ZN(n767) );
  NAND2_X1 U834 ( .A1(G111), .A2(n889), .ZN(n762) );
  NAND2_X1 U835 ( .A1(G99), .A2(n883), .ZN(n761) );
  NAND2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n765) );
  NAND2_X1 U837 ( .A1(n888), .A2(G123), .ZN(n763) );
  XOR2_X1 U838 ( .A(KEYINPUT18), .B(n763), .Z(n764) );
  NOR2_X1 U839 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U840 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U841 ( .A(n768), .B(KEYINPUT78), .ZN(n928) );
  XNOR2_X1 U842 ( .A(n928), .B(G2096), .ZN(n769) );
  OR2_X1 U843 ( .A1(G2100), .A2(n769), .ZN(G156) );
  INV_X1 U844 ( .A(G132), .ZN(G219) );
  INV_X1 U845 ( .A(G82), .ZN(G220) );
  INV_X1 U846 ( .A(G57), .ZN(G237) );
  XOR2_X1 U847 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n771) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n770) );
  XNOR2_X1 U849 ( .A(n771), .B(n770), .ZN(G223) );
  INV_X1 U850 ( .A(G223), .ZN(n828) );
  NAND2_X1 U851 ( .A1(n828), .A2(G567), .ZN(n772) );
  XOR2_X1 U852 ( .A(KEYINPUT11), .B(n772), .Z(G234) );
  INV_X1 U853 ( .A(G860), .ZN(n779) );
  OR2_X1 U854 ( .A1(n992), .A2(n779), .ZN(G153) );
  INV_X1 U855 ( .A(n977), .ZN(n787) );
  NOR2_X1 U856 ( .A1(n787), .A2(G868), .ZN(n773) );
  XNOR2_X1 U857 ( .A(n773), .B(KEYINPUT74), .ZN(n775) );
  INV_X1 U858 ( .A(G868), .ZN(n782) );
  NOR2_X1 U859 ( .A1(n782), .A2(G171), .ZN(n774) );
  NOR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U861 ( .A(KEYINPUT75), .B(n776), .ZN(G284) );
  NAND2_X1 U862 ( .A1(G868), .A2(G286), .ZN(n778) );
  NAND2_X1 U863 ( .A1(G299), .A2(n782), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n778), .A2(n777), .ZN(G297) );
  NAND2_X1 U865 ( .A1(n779), .A2(G559), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n780), .A2(n787), .ZN(n781) );
  XNOR2_X1 U867 ( .A(n781), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U868 ( .A1(G559), .A2(n782), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n787), .A2(n783), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n784), .B(KEYINPUT77), .ZN(n786) );
  NOR2_X1 U871 ( .A1(n992), .A2(G868), .ZN(n785) );
  NOR2_X1 U872 ( .A1(n786), .A2(n785), .ZN(G282) );
  NAND2_X1 U873 ( .A1(n787), .A2(G559), .ZN(n810) );
  XNOR2_X1 U874 ( .A(n992), .B(n810), .ZN(n788) );
  NOR2_X1 U875 ( .A1(n788), .A2(G860), .ZN(n800) );
  NAND2_X1 U876 ( .A1(n789), .A2(G80), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G93), .A2(n790), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n799) );
  NAND2_X1 U879 ( .A1(G67), .A2(n793), .ZN(n794) );
  XOR2_X1 U880 ( .A(KEYINPUT79), .B(n794), .Z(n797) );
  NAND2_X1 U881 ( .A1(n795), .A2(G55), .ZN(n796) );
  NAND2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n804) );
  XNOR2_X1 U884 ( .A(n800), .B(n804), .ZN(G145) );
  NOR2_X1 U885 ( .A1(G868), .A2(n804), .ZN(n801) );
  XNOR2_X1 U886 ( .A(n801), .B(KEYINPUT87), .ZN(n814) );
  XOR2_X1 U887 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n802) );
  XNOR2_X1 U888 ( .A(G288), .B(n802), .ZN(n806) );
  XOR2_X1 U889 ( .A(G166), .B(G305), .Z(n803) );
  XOR2_X1 U890 ( .A(n804), .B(n803), .Z(n805) );
  XNOR2_X1 U891 ( .A(n806), .B(n805), .ZN(n808) );
  XNOR2_X1 U892 ( .A(G290), .B(n975), .ZN(n807) );
  XNOR2_X1 U893 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U894 ( .A(n809), .B(n992), .ZN(n900) );
  XNOR2_X1 U895 ( .A(n900), .B(KEYINPUT86), .ZN(n811) );
  XNOR2_X1 U896 ( .A(n811), .B(n810), .ZN(n812) );
  NAND2_X1 U897 ( .A1(G868), .A2(n812), .ZN(n813) );
  NAND2_X1 U898 ( .A1(n814), .A2(n813), .ZN(G295) );
  NAND2_X1 U899 ( .A1(G2084), .A2(G2078), .ZN(n815) );
  XOR2_X1 U900 ( .A(KEYINPUT20), .B(n815), .Z(n816) );
  NAND2_X1 U901 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XNOR2_X1 U902 ( .A(KEYINPUT21), .B(n817), .ZN(n818) );
  NAND2_X1 U903 ( .A1(n818), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U904 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U905 ( .A1(G120), .A2(G69), .ZN(n819) );
  NOR2_X1 U906 ( .A1(G237), .A2(n819), .ZN(n820) );
  XNOR2_X1 U907 ( .A(KEYINPUT88), .B(n820), .ZN(n821) );
  NAND2_X1 U908 ( .A1(n821), .A2(G108), .ZN(n832) );
  NAND2_X1 U909 ( .A1(n832), .A2(G567), .ZN(n826) );
  NOR2_X1 U910 ( .A1(G220), .A2(G219), .ZN(n822) );
  XOR2_X1 U911 ( .A(KEYINPUT22), .B(n822), .Z(n823) );
  NOR2_X1 U912 ( .A1(G218), .A2(n823), .ZN(n824) );
  NAND2_X1 U913 ( .A1(G96), .A2(n824), .ZN(n833) );
  NAND2_X1 U914 ( .A1(n833), .A2(G2106), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n826), .A2(n825), .ZN(n853) );
  NAND2_X1 U916 ( .A1(G661), .A2(G483), .ZN(n827) );
  NOR2_X1 U917 ( .A1(n853), .A2(n827), .ZN(n831) );
  NAND2_X1 U918 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U921 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G108), .ZN(G238) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  INV_X1 U928 ( .A(G69), .ZN(G235) );
  NOR2_X1 U929 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U931 ( .A(G1966), .B(KEYINPUT41), .ZN(n843) );
  XOR2_X1 U932 ( .A(G1981), .B(G1956), .Z(n835) );
  XNOR2_X1 U933 ( .A(G1986), .B(G1961), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U935 ( .A(G1991), .B(G1976), .Z(n837) );
  XNOR2_X1 U936 ( .A(G1996), .B(G1971), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U938 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U939 ( .A(KEYINPUT108), .B(G2474), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(G229) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2090), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2072), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n846), .B(G2096), .Z(n848) );
  XNOR2_X1 U946 ( .A(G2084), .B(G2067), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U948 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n850) );
  XNOR2_X1 U949 ( .A(G2678), .B(G2100), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U951 ( .A(n852), .B(n851), .Z(G227) );
  INV_X1 U952 ( .A(n853), .ZN(G319) );
  NAND2_X1 U953 ( .A1(G136), .A2(n884), .ZN(n860) );
  NAND2_X1 U954 ( .A1(G112), .A2(n889), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G100), .A2(n883), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n858) );
  NAND2_X1 U957 ( .A1(n888), .A2(G124), .ZN(n856) );
  XOR2_X1 U958 ( .A(KEYINPUT44), .B(n856), .Z(n857) );
  NOR2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n861), .B(KEYINPUT109), .ZN(G162) );
  NAND2_X1 U962 ( .A1(n883), .A2(G103), .ZN(n862) );
  XOR2_X1 U963 ( .A(KEYINPUT111), .B(n862), .Z(n864) );
  NAND2_X1 U964 ( .A1(n884), .A2(G139), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U966 ( .A(KEYINPUT112), .B(n865), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G127), .A2(n888), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G115), .A2(n889), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(KEYINPUT113), .B(n868), .ZN(n869) );
  XNOR2_X1 U971 ( .A(KEYINPUT47), .B(n869), .ZN(n870) );
  NOR2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n920) );
  XNOR2_X1 U973 ( .A(n920), .B(n872), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(n880) );
  XOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n878) );
  XNOR2_X1 U977 ( .A(KEYINPUT115), .B(KEYINPUT114), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U979 ( .A(n880), .B(n879), .Z(n882) );
  XNOR2_X1 U980 ( .A(G164), .B(G160), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n898) );
  NAND2_X1 U982 ( .A1(G106), .A2(n883), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G142), .A2(n884), .ZN(n885) );
  NAND2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(KEYINPUT45), .ZN(n894) );
  NAND2_X1 U986 ( .A1(G130), .A2(n888), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G118), .A2(n889), .ZN(n890) );
  NAND2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT110), .B(n892), .Z(n893) );
  NAND2_X1 U990 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U991 ( .A(n895), .B(n928), .ZN(n896) );
  XOR2_X1 U992 ( .A(G162), .B(n896), .Z(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U994 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U995 ( .A(n900), .B(n977), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n901), .B(G286), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n902), .B(G171), .ZN(n903) );
  NOR2_X1 U998 ( .A1(G37), .A2(n903), .ZN(G397) );
  XNOR2_X1 U999 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(G229), .A2(G227), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n916) );
  XOR2_X1 U1002 ( .A(G2451), .B(G2430), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G2438), .B(G2443), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n913) );
  XOR2_X1 U1005 ( .A(G2435), .B(G2454), .Z(n909) );
  XNOR2_X1 U1006 ( .A(G1341), .B(G1348), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1008 ( .A(G2446), .B(G2427), .Z(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1010 ( .A(n913), .B(n912), .Z(n914) );
  NAND2_X1 U1011 ( .A1(G14), .A2(n914), .ZN(n919) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n919), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n919), .ZN(G401) );
  XOR2_X1 U1018 ( .A(G2072), .B(n920), .Z(n922) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n923), .B(KEYINPUT50), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n941) );
  XOR2_X1 U1023 ( .A(G2084), .B(G160), .Z(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n936) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n934) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(n932), .B(KEYINPUT51), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(n939), .B(KEYINPUT117), .ZN(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(n942), .ZN(n943) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n968) );
  NAND2_X1 U1036 ( .A1(n943), .A2(n968), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n944), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1038 ( .A(G25), .B(n945), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n946), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1040 ( .A(G32), .B(n947), .ZN(n956) );
  XNOR2_X1 U1041 ( .A(n948), .B(G27), .ZN(n954) );
  XNOR2_X1 U1042 ( .A(G2072), .B(KEYINPUT118), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(n949), .B(G33), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G26), .B(G2067), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(KEYINPUT119), .B(n952), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1050 ( .A(KEYINPUT120), .B(n959), .Z(n960) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n960), .ZN(n966) );
  XOR2_X1 U1052 ( .A(G34), .B(KEYINPUT121), .Z(n962) );
  XNOR2_X1 U1053 ( .A(G2084), .B(KEYINPUT54), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n962), .B(n961), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(n968), .B(n967), .ZN(n970) );
  INV_X1 U1059 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n971), .ZN(n1028) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT56), .ZN(n999) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G168), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(KEYINPUT57), .B(n974), .ZN(n997) );
  XNOR2_X1 U1066 ( .A(n975), .B(G1956), .ZN(n990) );
  XNOR2_X1 U1067 ( .A(G1961), .B(G171), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT122), .ZN(n985) );
  XNOR2_X1 U1069 ( .A(G1348), .B(n977), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1074 ( .A(G1971), .B(G303), .Z(n986) );
  XNOR2_X1 U1075 ( .A(KEYINPUT123), .B(n986), .ZN(n987) );
  NOR2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(KEYINPUT124), .B(n991), .ZN(n995) );
  XOR2_X1 U1079 ( .A(G1341), .B(n992), .Z(n993) );
  XNOR2_X1 U1080 ( .A(KEYINPUT125), .B(n993), .ZN(n994) );
  NOR2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1082 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1083 ( .A1(n999), .A2(n998), .ZN(n1026) );
  INV_X1 U1084 ( .A(G16), .ZN(n1024) );
  XOR2_X1 U1085 ( .A(G1976), .B(G23), .Z(n1003) );
  XNOR2_X1 U1086 ( .A(G1986), .B(G24), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(n1005), .B(n1004), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G1961), .B(G5), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1021) );
  XOR2_X1 U1096 ( .A(G1348), .B(KEYINPUT59), .Z(n1010) );
  XNOR2_X1 U1097 ( .A(G4), .B(n1010), .ZN(n1018) );
  XOR2_X1 U1098 ( .A(G1341), .B(G19), .Z(n1013) );
  XNOR2_X1 U1099 ( .A(n1011), .B(G20), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(G6), .B(G1981), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT126), .B(n1016), .Z(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(KEYINPUT60), .B(n1019), .Z(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1110 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1111 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

