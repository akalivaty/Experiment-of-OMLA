

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XNOR2_X1 U324 ( .A(n481), .B(n480), .ZN(n534) );
  XNOR2_X1 U325 ( .A(n418), .B(G92GAT), .ZN(n419) );
  NOR2_X1 U326 ( .A1(n522), .A2(n521), .ZN(n530) );
  XOR2_X1 U327 ( .A(n366), .B(n365), .Z(n525) );
  XOR2_X1 U328 ( .A(KEYINPUT102), .B(n370), .Z(n292) );
  XNOR2_X1 U329 ( .A(KEYINPUT101), .B(n367), .ZN(n293) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n356) );
  INV_X1 U331 ( .A(KEYINPUT64), .ZN(n479) );
  XNOR2_X1 U332 ( .A(n356), .B(G36GAT), .ZN(n399) );
  INV_X1 U333 ( .A(G71GAT), .ZN(n343) );
  XNOR2_X1 U334 ( .A(n479), .B(KEYINPUT48), .ZN(n480) );
  XNOR2_X1 U335 ( .A(n445), .B(KEYINPUT20), .ZN(n346) );
  XNOR2_X1 U336 ( .A(n344), .B(n343), .ZN(n445) );
  XNOR2_X1 U337 ( .A(n350), .B(n349), .ZN(n351) );
  NOR2_X1 U338 ( .A1(n523), .A2(n484), .ZN(n575) );
  OR2_X1 U339 ( .A1(n485), .A2(n527), .ZN(n355) );
  XNOR2_X1 U340 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U341 ( .A(n420), .B(n419), .ZN(n473) );
  NOR2_X1 U342 ( .A1(n538), .A2(n487), .ZN(n571) );
  XNOR2_X1 U343 ( .A(n461), .B(n460), .ZN(n507) );
  XNOR2_X1 U344 ( .A(n488), .B(G176GAT), .ZN(n489) );
  XNOR2_X1 U345 ( .A(n464), .B(KEYINPUT108), .ZN(n465) );
  XNOR2_X1 U346 ( .A(n490), .B(n489), .ZN(G1349GAT) );
  XNOR2_X1 U347 ( .A(n466), .B(n465), .ZN(G1330GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT5), .B(G57GAT), .Z(n295) );
  XNOR2_X1 U349 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n294) );
  XNOR2_X1 U350 ( .A(n295), .B(n294), .ZN(n313) );
  XOR2_X1 U351 ( .A(G148GAT), .B(G162GAT), .Z(n297) );
  XNOR2_X1 U352 ( .A(G29GAT), .B(G134GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U354 ( .A(KEYINPUT97), .B(G120GAT), .Z(n299) );
  XNOR2_X1 U355 ( .A(G155GAT), .B(G127GAT), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U357 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U358 ( .A(KEYINPUT4), .B(G1GAT), .Z(n303) );
  NAND2_X1 U359 ( .A1(G225GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U361 ( .A(KEYINPUT98), .B(n304), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT0), .B(G113GAT), .ZN(n349) );
  XNOR2_X1 U364 ( .A(n307), .B(n349), .ZN(n311) );
  XOR2_X1 U365 ( .A(KEYINPUT78), .B(G85GAT), .Z(n413) );
  XOR2_X1 U366 ( .A(G141GAT), .B(KEYINPUT2), .Z(n309) );
  XNOR2_X1 U367 ( .A(KEYINPUT3), .B(KEYINPUT95), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n413), .B(n314), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U371 ( .A(n313), .B(n312), .Z(n523) );
  XOR2_X1 U372 ( .A(G162GAT), .B(G50GAT), .Z(n410) );
  XOR2_X1 U373 ( .A(n410), .B(n314), .Z(n316) );
  NAND2_X1 U374 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n329) );
  XOR2_X1 U376 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n318) );
  XNOR2_X1 U377 ( .A(KEYINPUT90), .B(KEYINPUT23), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n320) );
  INV_X1 U379 ( .A(KEYINPUT96), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n322) );
  XOR2_X1 U381 ( .A(G155GAT), .B(G22GAT), .Z(n387) );
  XNOR2_X1 U382 ( .A(n387), .B(KEYINPUT91), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U384 ( .A(n323), .B(G204GAT), .Z(n327) );
  XOR2_X1 U385 ( .A(KEYINPUT75), .B(G78GAT), .Z(n325) );
  XNOR2_X1 U386 ( .A(G148GAT), .B(G106GAT), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n446) );
  XNOR2_X1 U388 ( .A(G211GAT), .B(n446), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n334) );
  XOR2_X1 U391 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n331) );
  XNOR2_X1 U392 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n333) );
  XOR2_X1 U394 ( .A(G218GAT), .B(KEYINPUT92), .Z(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n365) );
  XOR2_X1 U396 ( .A(n334), .B(n365), .Z(n485) );
  XOR2_X1 U397 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n336) );
  XNOR2_X1 U398 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U400 ( .A(n337), .B(G169GAT), .Z(n339) );
  XNOR2_X1 U401 ( .A(G183GAT), .B(G176GAT), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n362) );
  XOR2_X1 U403 ( .A(KEYINPUT83), .B(KEYINPUT85), .Z(n341) );
  XNOR2_X1 U404 ( .A(KEYINPUT86), .B(KEYINPUT88), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n362), .B(n342), .ZN(n354) );
  XOR2_X1 U407 ( .A(G120GAT), .B(G99GAT), .Z(n344) );
  AND2_X1 U408 ( .A1(G227GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n352) );
  XOR2_X1 U410 ( .A(G127GAT), .B(G15GAT), .Z(n386) );
  XOR2_X1 U411 ( .A(KEYINPUT84), .B(n386), .Z(n348) );
  XNOR2_X1 U412 ( .A(G134GAT), .B(G43GAT), .ZN(n398) );
  INV_X1 U413 ( .A(n398), .ZN(n400) );
  XNOR2_X1 U414 ( .A(G190GAT), .B(n400), .ZN(n347) );
  XNOR2_X1 U415 ( .A(n348), .B(n347), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n538) );
  INV_X1 U417 ( .A(n538), .ZN(n527) );
  XOR2_X1 U418 ( .A(KEYINPUT26), .B(n355), .Z(n574) );
  XOR2_X1 U419 ( .A(n399), .B(KEYINPUT99), .Z(n358) );
  NAND2_X1 U420 ( .A1(G226GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n360) );
  XNOR2_X1 U422 ( .A(G92GAT), .B(G64GAT), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n359), .B(G204GAT), .ZN(n453) );
  XOR2_X1 U424 ( .A(n360), .B(n453), .Z(n364) );
  XNOR2_X1 U425 ( .A(G211GAT), .B(G8GAT), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n361), .B(KEYINPUT79), .ZN(n383) );
  XNOR2_X1 U427 ( .A(n383), .B(n362), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n364), .B(n363), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n525), .B(KEYINPUT27), .ZN(n374) );
  AND2_X1 U430 ( .A1(n574), .A2(n374), .ZN(n367) );
  NAND2_X1 U431 ( .A1(n525), .A2(n527), .ZN(n368) );
  NAND2_X1 U432 ( .A1(n368), .A2(n485), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n369), .B(KEYINPUT25), .ZN(n370) );
  NAND2_X1 U434 ( .A1(n293), .A2(n292), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n371), .B(KEYINPUT103), .ZN(n372) );
  NOR2_X1 U436 ( .A1(n523), .A2(n372), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n373), .B(KEYINPUT104), .ZN(n379) );
  NAND2_X1 U438 ( .A1(n523), .A2(n374), .ZN(n533) );
  XNOR2_X1 U439 ( .A(KEYINPUT89), .B(n527), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n485), .B(KEYINPUT28), .ZN(n536) );
  NAND2_X1 U441 ( .A1(n375), .A2(n536), .ZN(n376) );
  NOR2_X1 U442 ( .A1(n533), .A2(n376), .ZN(n377) );
  XNOR2_X1 U443 ( .A(KEYINPUT100), .B(n377), .ZN(n378) );
  NOR2_X1 U444 ( .A1(n379), .A2(n378), .ZN(n494) );
  XOR2_X1 U445 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n381) );
  XNOR2_X1 U446 ( .A(G1GAT), .B(G71GAT), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n381), .B(n380), .ZN(n397) );
  XNOR2_X1 U448 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n382), .B(KEYINPUT73), .ZN(n454) );
  XNOR2_X1 U450 ( .A(n383), .B(n454), .ZN(n395) );
  XOR2_X1 U451 ( .A(G64GAT), .B(KEYINPUT81), .Z(n385) );
  XNOR2_X1 U452 ( .A(KEYINPUT14), .B(KEYINPUT80), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n391) );
  XOR2_X1 U454 ( .A(G183GAT), .B(G78GAT), .Z(n389) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U457 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U458 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n561) );
  NOR2_X1 U462 ( .A1(n494), .A2(n561), .ZN(n422) );
  NAND2_X1 U463 ( .A1(n399), .A2(n398), .ZN(n403) );
  INV_X1 U464 ( .A(n399), .ZN(n401) );
  NAND2_X1 U465 ( .A1(n401), .A2(n400), .ZN(n402) );
  NAND2_X1 U466 ( .A1(n403), .A2(n402), .ZN(n405) );
  NAND2_X1 U467 ( .A1(G232GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U469 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n407) );
  XNOR2_X1 U470 ( .A(KEYINPUT77), .B(G99GAT), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n415) );
  XNOR2_X1 U473 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U475 ( .A(n413), .B(n412), .Z(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n420) );
  XOR2_X1 U477 ( .A(KEYINPUT7), .B(KEYINPUT71), .Z(n417) );
  XNOR2_X1 U478 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n435) );
  XOR2_X1 U480 ( .A(n435), .B(G106GAT), .Z(n418) );
  XNOR2_X1 U481 ( .A(n473), .B(KEYINPUT105), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n421), .B(KEYINPUT36), .ZN(n588) );
  NAND2_X1 U483 ( .A1(n422), .A2(n588), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n423), .B(KEYINPUT37), .ZN(n520) );
  XOR2_X1 U485 ( .A(G197GAT), .B(G15GAT), .Z(n425) );
  XNOR2_X1 U486 ( .A(G113GAT), .B(G22GAT), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U488 ( .A(KEYINPUT70), .B(G169GAT), .Z(n427) );
  XNOR2_X1 U489 ( .A(G1GAT), .B(G8GAT), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U491 ( .A(n429), .B(n428), .Z(n434) );
  XOR2_X1 U492 ( .A(KEYINPUT68), .B(KEYINPUT72), .Z(n431) );
  NAND2_X1 U493 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U495 ( .A(KEYINPUT30), .B(n432), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n439) );
  XOR2_X1 U497 ( .A(G43GAT), .B(G36GAT), .Z(n437) );
  XNOR2_X1 U498 ( .A(G50GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U500 ( .A(n439), .B(n438), .Z(n444) );
  XOR2_X1 U501 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n441) );
  XNOR2_X1 U502 ( .A(KEYINPUT69), .B(KEYINPUT66), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U504 ( .A(G141GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U505 ( .A(n444), .B(n443), .ZN(n566) );
  XOR2_X1 U506 ( .A(n446), .B(n445), .Z(n458) );
  XOR2_X1 U507 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n448) );
  XNOR2_X1 U508 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U510 ( .A(G176GAT), .B(G85GAT), .Z(n450) );
  NAND2_X1 U511 ( .A1(G230GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U513 ( .A(n452), .B(n451), .Z(n456) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(n580) );
  NAND2_X1 U517 ( .A1(n566), .A2(n580), .ZN(n459) );
  XOR2_X1 U518 ( .A(KEYINPUT76), .B(n459), .Z(n495) );
  NAND2_X1 U519 ( .A1(n520), .A2(n495), .ZN(n461) );
  XOR2_X1 U520 ( .A(KEYINPUT38), .B(KEYINPUT106), .Z(n460) );
  NAND2_X1 U521 ( .A1(n507), .A2(n527), .ZN(n466) );
  XOR2_X1 U522 ( .A(KEYINPUT40), .B(KEYINPUT110), .Z(n463) );
  XNOR2_X1 U523 ( .A(G43GAT), .B(KEYINPUT109), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U525 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n468) );
  NAND2_X1 U526 ( .A1(n588), .A2(n561), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n468), .B(n467), .ZN(n469) );
  NOR2_X1 U528 ( .A1(n566), .A2(n469), .ZN(n470) );
  NAND2_X1 U529 ( .A1(n580), .A2(n470), .ZN(n478) );
  XOR2_X1 U530 ( .A(KEYINPUT47), .B(KEYINPUT114), .Z(n476) );
  XOR2_X1 U531 ( .A(KEYINPUT113), .B(n561), .Z(n568) );
  XNOR2_X1 U532 ( .A(KEYINPUT41), .B(n580), .ZN(n557) );
  NAND2_X1 U533 ( .A1(n566), .A2(n557), .ZN(n471) );
  XOR2_X1 U534 ( .A(KEYINPUT46), .B(n471), .Z(n472) );
  NOR2_X1 U535 ( .A1(n568), .A2(n472), .ZN(n474) );
  INV_X1 U536 ( .A(n473), .ZN(n570) );
  NAND2_X1 U537 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U538 ( .A(n476), .B(n475), .ZN(n477) );
  NAND2_X1 U539 ( .A1(n478), .A2(n477), .ZN(n481) );
  XOR2_X1 U540 ( .A(KEYINPUT124), .B(n525), .Z(n482) );
  NOR2_X1 U541 ( .A1(n534), .A2(n482), .ZN(n483) );
  XOR2_X1 U542 ( .A(KEYINPUT54), .B(n483), .Z(n484) );
  NAND2_X1 U543 ( .A1(n485), .A2(n575), .ZN(n486) );
  XOR2_X1 U544 ( .A(KEYINPUT55), .B(n486), .Z(n487) );
  NAND2_X1 U545 ( .A1(n571), .A2(n557), .ZN(n490) );
  XOR2_X1 U546 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n488) );
  NAND2_X1 U547 ( .A1(n561), .A2(n473), .ZN(n491) );
  XNOR2_X1 U548 ( .A(n491), .B(KEYINPUT82), .ZN(n492) );
  XNOR2_X1 U549 ( .A(n492), .B(KEYINPUT16), .ZN(n493) );
  NOR2_X1 U550 ( .A1(n494), .A2(n493), .ZN(n509) );
  AND2_X1 U551 ( .A1(n509), .A2(n495), .ZN(n501) );
  NAND2_X1 U552 ( .A1(n501), .A2(n523), .ZN(n496) );
  XNOR2_X1 U553 ( .A(n496), .B(KEYINPUT34), .ZN(n497) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(n497), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n525), .A2(n501), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n498), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(G15GAT), .B(KEYINPUT35), .Z(n500) );
  NAND2_X1 U558 ( .A1(n501), .A2(n527), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  INV_X1 U560 ( .A(n536), .ZN(n529) );
  NAND2_X1 U561 ( .A1(n501), .A2(n529), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U563 ( .A1(n507), .A2(n523), .ZN(n505) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(KEYINPUT39), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n525), .A2(n507), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U569 ( .A1(n529), .A2(n507), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G50GAT), .B(n508), .ZN(G1331GAT) );
  INV_X1 U571 ( .A(n566), .ZN(n576) );
  NAND2_X1 U572 ( .A1(n557), .A2(n576), .ZN(n521) );
  INV_X1 U573 ( .A(n509), .ZN(n510) );
  NOR2_X1 U574 ( .A1(n521), .A2(n510), .ZN(n516) );
  NAND2_X1 U575 ( .A1(n523), .A2(n516), .ZN(n511) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(n511), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  XOR2_X1 U578 ( .A(G64GAT), .B(KEYINPUT111), .Z(n514) );
  NAND2_X1 U579 ( .A1(n516), .A2(n525), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n527), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U584 ( .A1(n516), .A2(n529), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n519), .ZN(G1335GAT) );
  INV_X1 U587 ( .A(n520), .ZN(n522) );
  NAND2_X1 U588 ( .A1(n530), .A2(n523), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n525), .A2(n530), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n540) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U599 ( .A(KEYINPUT115), .B(n535), .Z(n551) );
  NAND2_X1 U600 ( .A1(n551), .A2(n536), .ZN(n537) );
  NOR2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n566), .A2(n547), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n542) );
  NAND2_X1 U605 ( .A1(n547), .A2(n557), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U607 ( .A(G120GAT), .B(n543), .Z(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n545) );
  NAND2_X1 U609 ( .A1(n547), .A2(n568), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n549) );
  NAND2_X1 U613 ( .A1(n547), .A2(n570), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U615 ( .A(G134GAT), .B(n550), .Z(G1343GAT) );
  NAND2_X1 U616 ( .A1(n551), .A2(n574), .ZN(n564) );
  NOR2_X1 U617 ( .A1(n576), .A2(n564), .ZN(n553) );
  XNOR2_X1 U618 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT122), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n560) );
  INV_X1 U624 ( .A(n557), .ZN(n558) );
  NOR2_X1 U625 ( .A1(n558), .A2(n564), .ZN(n559) );
  XOR2_X1 U626 ( .A(n560), .B(n559), .Z(G1345GAT) );
  INV_X1 U627 ( .A(n561), .ZN(n584) );
  NOR2_X1 U628 ( .A1(n584), .A2(n564), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G155GAT), .B(KEYINPUT123), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1346GAT) );
  NOR2_X1 U631 ( .A1(n473), .A2(n564), .ZN(n565) );
  XOR2_X1 U632 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NAND2_X1 U633 ( .A1(n571), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n568), .A2(n571), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1351GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n587) );
  NOR2_X1 U641 ( .A1(n576), .A2(n587), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n587), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n587), .ZN(n585) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n585), .Z(n586) );
  XNOR2_X1 U651 ( .A(KEYINPUT126), .B(n586), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n591) );
  INV_X1 U653 ( .A(n587), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

