

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U556 ( .A(G2104), .ZN(n526) );
  INV_X1 U557 ( .A(n664), .ZN(n618) );
  NOR2_X2 U558 ( .A1(G2105), .A2(n526), .ZN(n888) );
  AND2_X1 U559 ( .A1(n533), .A2(n532), .ZN(G160) );
  NOR2_X1 U560 ( .A1(G651), .A2(G543), .ZN(n788) );
  INV_X1 U561 ( .A(KEYINPUT28), .ZN(n608) );
  NOR2_X1 U562 ( .A1(G651), .A2(n573), .ZN(n792) );
  XNOR2_X1 U563 ( .A(n761), .B(KEYINPUT99), .ZN(n762) );
  XNOR2_X1 U564 ( .A(n763), .B(n762), .ZN(G329) );
  INV_X1 U565 ( .A(KEYINPUT67), .ZN(n523) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X2 U567 ( .A(KEYINPUT17), .B(n521), .Z(n886) );
  NAND2_X1 U568 ( .A1(n886), .A2(G137), .ZN(n522) );
  XNOR2_X1 U569 ( .A(n523), .B(n522), .ZN(n533) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(KEYINPUT66), .Z(n525) );
  NAND2_X1 U571 ( .A1(G101), .A2(n888), .ZN(n524) );
  XOR2_X1 U572 ( .A(n525), .B(n524), .Z(n531) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U574 ( .A1(G113), .A2(n882), .ZN(n529) );
  NAND2_X1 U575 ( .A1(n526), .A2(G2105), .ZN(n527) );
  XNOR2_X1 U576 ( .A(n527), .B(KEYINPUT65), .ZN(n883) );
  NAND2_X1 U577 ( .A1(G125), .A2(n883), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U580 ( .A1(G91), .A2(n788), .ZN(n535) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n573) );
  INV_X1 U582 ( .A(G651), .ZN(n537) );
  NOR2_X1 U583 ( .A1(n573), .A2(n537), .ZN(n789) );
  NAND2_X1 U584 ( .A1(G78), .A2(n789), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U586 ( .A(KEYINPUT72), .B(n536), .Z(n542) );
  NOR2_X1 U587 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n538), .Z(n794) );
  NAND2_X1 U589 ( .A1(G65), .A2(n794), .ZN(n540) );
  NAND2_X1 U590 ( .A1(G53), .A2(n792), .ZN(n539) );
  AND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(G299) );
  XNOR2_X1 U593 ( .A(KEYINPUT71), .B(KEYINPUT9), .ZN(n546) );
  NAND2_X1 U594 ( .A1(G90), .A2(n788), .ZN(n544) );
  NAND2_X1 U595 ( .A1(G77), .A2(n789), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U597 ( .A(n546), .B(n545), .ZN(n550) );
  NAND2_X1 U598 ( .A1(G64), .A2(n794), .ZN(n548) );
  NAND2_X1 U599 ( .A1(G52), .A2(n792), .ZN(n547) );
  NAND2_X1 U600 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U601 ( .A1(n550), .A2(n549), .ZN(G171) );
  NAND2_X1 U602 ( .A1(G63), .A2(n794), .ZN(n552) );
  NAND2_X1 U603 ( .A1(G51), .A2(n792), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U605 ( .A(KEYINPUT6), .B(n553), .ZN(n561) );
  NAND2_X1 U606 ( .A1(G89), .A2(n788), .ZN(n554) );
  XNOR2_X1 U607 ( .A(n554), .B(KEYINPUT74), .ZN(n555) );
  XNOR2_X1 U608 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U609 ( .A1(G76), .A2(n789), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U611 ( .A(KEYINPUT75), .B(n558), .ZN(n559) );
  XNOR2_X1 U612 ( .A(KEYINPUT5), .B(n559), .ZN(n560) );
  NOR2_X1 U613 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U614 ( .A(KEYINPUT7), .B(n562), .Z(G168) );
  NAND2_X1 U615 ( .A1(G88), .A2(n788), .ZN(n564) );
  NAND2_X1 U616 ( .A1(G75), .A2(n789), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U618 ( .A1(G62), .A2(n794), .ZN(n566) );
  NAND2_X1 U619 ( .A1(G50), .A2(n792), .ZN(n565) );
  NAND2_X1 U620 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U621 ( .A1(n568), .A2(n567), .ZN(G166) );
  XNOR2_X1 U622 ( .A(KEYINPUT83), .B(G166), .ZN(G303) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U624 ( .A1(G49), .A2(n792), .ZN(n570) );
  NAND2_X1 U625 ( .A1(G74), .A2(G651), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U627 ( .A(KEYINPUT77), .B(n571), .Z(n572) );
  NOR2_X1 U628 ( .A1(n794), .A2(n572), .ZN(n575) );
  NAND2_X1 U629 ( .A1(n573), .A2(G87), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n575), .A2(n574), .ZN(G288) );
  XOR2_X1 U631 ( .A(KEYINPUT79), .B(KEYINPUT2), .Z(n577) );
  NAND2_X1 U632 ( .A1(G73), .A2(n789), .ZN(n576) );
  XNOR2_X1 U633 ( .A(n577), .B(n576), .ZN(n584) );
  NAND2_X1 U634 ( .A1(G48), .A2(n792), .ZN(n579) );
  NAND2_X1 U635 ( .A1(G86), .A2(n788), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U637 ( .A1(n794), .A2(G61), .ZN(n580) );
  XOR2_X1 U638 ( .A(KEYINPUT78), .B(n580), .Z(n581) );
  NOR2_X1 U639 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U640 ( .A1(n584), .A2(n583), .ZN(G305) );
  NAND2_X1 U641 ( .A1(G85), .A2(n788), .ZN(n585) );
  XNOR2_X1 U642 ( .A(n585), .B(KEYINPUT68), .ZN(n593) );
  NAND2_X1 U643 ( .A1(G60), .A2(n794), .ZN(n587) );
  NAND2_X1 U644 ( .A1(G47), .A2(n792), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U646 ( .A(KEYINPUT70), .B(n588), .ZN(n591) );
  NAND2_X1 U647 ( .A1(G72), .A2(n789), .ZN(n589) );
  XNOR2_X1 U648 ( .A(KEYINPUT69), .B(n589), .ZN(n590) );
  NOR2_X1 U649 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U650 ( .A1(n593), .A2(n592), .ZN(G290) );
  NAND2_X1 U651 ( .A1(G102), .A2(n888), .ZN(n595) );
  NAND2_X1 U652 ( .A1(G138), .A2(n886), .ZN(n594) );
  NAND2_X1 U653 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U654 ( .A1(G114), .A2(n882), .ZN(n597) );
  NAND2_X1 U655 ( .A1(G126), .A2(n883), .ZN(n596) );
  NAND2_X1 U656 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U657 ( .A1(n599), .A2(n598), .ZN(G164) );
  NOR2_X1 U658 ( .A1(G164), .A2(G1384), .ZN(n697) );
  AND2_X1 U659 ( .A1(n697), .A2(G40), .ZN(n600) );
  AND2_X1 U660 ( .A1(n600), .A2(G160), .ZN(n602) );
  INV_X1 U661 ( .A(KEYINPUT64), .ZN(n601) );
  XNOR2_X2 U662 ( .A(n602), .B(n601), .ZN(n664) );
  NAND2_X1 U663 ( .A1(n664), .A2(G1956), .ZN(n603) );
  XNOR2_X1 U664 ( .A(n603), .B(KEYINPUT88), .ZN(n606) );
  NAND2_X1 U665 ( .A1(G2072), .A2(n618), .ZN(n604) );
  XOR2_X1 U666 ( .A(KEYINPUT27), .B(n604), .Z(n605) );
  NAND2_X1 U667 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U668 ( .A(n607), .B(KEYINPUT89), .ZN(n610) );
  INV_X1 U669 ( .A(G299), .ZN(n803) );
  NOR2_X1 U670 ( .A1(n610), .A2(n803), .ZN(n609) );
  XNOR2_X1 U671 ( .A(n609), .B(n608), .ZN(n646) );
  NAND2_X1 U672 ( .A1(n610), .A2(n803), .ZN(n644) );
  NAND2_X1 U673 ( .A1(G54), .A2(n792), .ZN(n612) );
  NAND2_X1 U674 ( .A1(G79), .A2(n789), .ZN(n611) );
  NAND2_X1 U675 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U676 ( .A1(G66), .A2(n794), .ZN(n614) );
  NAND2_X1 U677 ( .A1(G92), .A2(n788), .ZN(n613) );
  NAND2_X1 U678 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U679 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U680 ( .A(n617), .B(KEYINPUT15), .ZN(n994) );
  NAND2_X1 U681 ( .A1(G2067), .A2(n618), .ZN(n620) );
  NAND2_X1 U682 ( .A1(n664), .A2(G1348), .ZN(n619) );
  NAND2_X1 U683 ( .A1(n620), .A2(n619), .ZN(n636) );
  NOR2_X1 U684 ( .A1(n994), .A2(n636), .ZN(n642) );
  INV_X1 U685 ( .A(G1341), .ZN(n1004) );
  XNOR2_X1 U686 ( .A(KEYINPUT26), .B(KEYINPUT90), .ZN(n625) );
  NAND2_X1 U687 ( .A1(n1004), .A2(n625), .ZN(n621) );
  NAND2_X1 U688 ( .A1(n621), .A2(n664), .ZN(n624) );
  AND2_X1 U689 ( .A1(n618), .A2(G1996), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n622), .A2(n625), .ZN(n623) );
  NAND2_X1 U691 ( .A1(n624), .A2(n623), .ZN(n640) );
  NOR2_X1 U692 ( .A1(G1996), .A2(n625), .ZN(n635) );
  NAND2_X1 U693 ( .A1(G56), .A2(n794), .ZN(n626) );
  XOR2_X1 U694 ( .A(KEYINPUT14), .B(n626), .Z(n632) );
  NAND2_X1 U695 ( .A1(n788), .A2(G81), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n627), .B(KEYINPUT12), .ZN(n629) );
  NAND2_X1 U697 ( .A1(G68), .A2(n789), .ZN(n628) );
  NAND2_X1 U698 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U699 ( .A(KEYINPUT13), .B(n630), .Z(n631) );
  NOR2_X1 U700 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U701 ( .A1(n792), .A2(G43), .ZN(n633) );
  NAND2_X1 U702 ( .A1(n634), .A2(n633), .ZN(n978) );
  NOR2_X1 U703 ( .A1(n635), .A2(n978), .ZN(n638) );
  NAND2_X1 U704 ( .A1(n994), .A2(n636), .ZN(n637) );
  NAND2_X1 U705 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U706 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U707 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U708 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U709 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U710 ( .A(KEYINPUT29), .B(n647), .Z(n651) );
  XNOR2_X1 U711 ( .A(G2078), .B(KEYINPUT25), .ZN(n958) );
  NAND2_X1 U712 ( .A1(n618), .A2(n958), .ZN(n649) );
  INV_X1 U713 ( .A(G1961), .ZN(n1013) );
  NAND2_X1 U714 ( .A1(n664), .A2(n1013), .ZN(n648) );
  NAND2_X1 U715 ( .A1(n649), .A2(n648), .ZN(n655) );
  NAND2_X1 U716 ( .A1(G171), .A2(n655), .ZN(n650) );
  NAND2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n672) );
  NAND2_X1 U718 ( .A1(n664), .A2(G8), .ZN(n737) );
  NOR2_X1 U719 ( .A1(G1966), .A2(n737), .ZN(n660) );
  NOR2_X1 U720 ( .A1(n664), .A2(G2084), .ZN(n659) );
  NOR2_X1 U721 ( .A1(n660), .A2(n659), .ZN(n652) );
  NAND2_X1 U722 ( .A1(G8), .A2(n652), .ZN(n653) );
  XNOR2_X1 U723 ( .A(KEYINPUT30), .B(n653), .ZN(n654) );
  NOR2_X1 U724 ( .A1(G168), .A2(n654), .ZN(n657) );
  NOR2_X1 U725 ( .A1(G171), .A2(n655), .ZN(n656) );
  NOR2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U727 ( .A(KEYINPUT31), .B(n658), .Z(n670) );
  AND2_X1 U728 ( .A1(n672), .A2(n670), .ZN(n663) );
  AND2_X1 U729 ( .A1(G8), .A2(n659), .ZN(n661) );
  OR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  OR2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n680) );
  NOR2_X1 U732 ( .A1(n664), .A2(G2090), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(KEYINPUT91), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n666), .A2(G303), .ZN(n668) );
  NOR2_X1 U735 ( .A1(G1971), .A2(n737), .ZN(n667) );
  NOR2_X1 U736 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U737 ( .A(KEYINPUT92), .B(n669), .Z(n673) );
  AND2_X1 U738 ( .A1(n670), .A2(n673), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n672), .A2(n671), .ZN(n677) );
  INV_X1 U740 ( .A(n673), .ZN(n674) );
  OR2_X1 U741 ( .A1(n674), .A2(G286), .ZN(n675) );
  AND2_X1 U742 ( .A1(n675), .A2(G8), .ZN(n676) );
  NAND2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U744 ( .A(n678), .B(KEYINPUT32), .ZN(n679) );
  NAND2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n732) );
  NOR2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n690) );
  NOR2_X1 U747 ( .A1(G1971), .A2(G303), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n690), .A2(n681), .ZN(n988) );
  XOR2_X1 U749 ( .A(n988), .B(KEYINPUT93), .Z(n682) );
  NAND2_X1 U750 ( .A1(n732), .A2(n682), .ZN(n683) );
  NAND2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n984) );
  NAND2_X1 U752 ( .A1(n683), .A2(n984), .ZN(n684) );
  XNOR2_X1 U753 ( .A(KEYINPUT94), .B(n684), .ZN(n686) );
  OR2_X1 U754 ( .A1(n737), .A2(KEYINPUT95), .ZN(n685) );
  NOR2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U756 ( .A1(n687), .A2(KEYINPUT33), .ZN(n695) );
  INV_X1 U757 ( .A(KEYINPUT95), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n690), .A2(KEYINPUT33), .ZN(n688) );
  NAND2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n690), .A2(KEYINPUT95), .ZN(n691) );
  NAND2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U762 ( .A1(n737), .A2(n693), .ZN(n694) );
  NOR2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n729) );
  XOR2_X1 U764 ( .A(G1981), .B(G305), .Z(n979) );
  XNOR2_X1 U765 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n696) );
  NOR2_X1 U767 ( .A1(n697), .A2(n696), .ZN(n755) );
  NAND2_X1 U768 ( .A1(n990), .A2(n755), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n698), .B(KEYINPUT84), .ZN(n716) );
  NAND2_X1 U770 ( .A1(G131), .A2(n886), .ZN(n700) );
  NAND2_X1 U771 ( .A1(G119), .A2(n883), .ZN(n699) );
  NAND2_X1 U772 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U773 ( .A1(G95), .A2(n888), .ZN(n702) );
  NAND2_X1 U774 ( .A1(G107), .A2(n882), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U777 ( .A(n705), .B(KEYINPUT85), .ZN(n879) );
  XNOR2_X1 U778 ( .A(KEYINPUT86), .B(G1991), .ZN(n964) );
  NAND2_X1 U779 ( .A1(n879), .A2(n964), .ZN(n715) );
  NAND2_X1 U780 ( .A1(G117), .A2(n882), .ZN(n707) );
  NAND2_X1 U781 ( .A1(G129), .A2(n883), .ZN(n706) );
  NAND2_X1 U782 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U783 ( .A1(n888), .A2(G105), .ZN(n708) );
  XOR2_X1 U784 ( .A(KEYINPUT38), .B(n708), .Z(n709) );
  NOR2_X1 U785 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U786 ( .A(KEYINPUT87), .B(n711), .Z(n713) );
  NAND2_X1 U787 ( .A1(n886), .A2(G141), .ZN(n712) );
  NAND2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n866) );
  NAND2_X1 U789 ( .A1(G1996), .A2(n866), .ZN(n714) );
  NAND2_X1 U790 ( .A1(n715), .A2(n714), .ZN(n922) );
  NAND2_X1 U791 ( .A1(n755), .A2(n922), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n716), .A2(n744), .ZN(n741) );
  INV_X1 U793 ( .A(n741), .ZN(n717) );
  AND2_X1 U794 ( .A1(n979), .A2(n717), .ZN(n727) );
  NAND2_X1 U795 ( .A1(G104), .A2(n888), .ZN(n719) );
  NAND2_X1 U796 ( .A1(G140), .A2(n886), .ZN(n718) );
  NAND2_X1 U797 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U798 ( .A(KEYINPUT34), .B(n720), .ZN(n725) );
  NAND2_X1 U799 ( .A1(G116), .A2(n882), .ZN(n722) );
  NAND2_X1 U800 ( .A1(G128), .A2(n883), .ZN(n721) );
  NAND2_X1 U801 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U802 ( .A(KEYINPUT35), .B(n723), .Z(n724) );
  NOR2_X1 U803 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U804 ( .A(KEYINPUT36), .B(n726), .ZN(n896) );
  XNOR2_X1 U805 ( .A(G2067), .B(KEYINPUT37), .ZN(n753) );
  NOR2_X1 U806 ( .A1(n896), .A2(n753), .ZN(n923) );
  NAND2_X1 U807 ( .A1(n923), .A2(n755), .ZN(n752) );
  AND2_X1 U808 ( .A1(n727), .A2(n752), .ZN(n728) );
  NAND2_X1 U809 ( .A1(n729), .A2(n728), .ZN(n760) );
  INV_X1 U810 ( .A(n752), .ZN(n743) );
  NOR2_X1 U811 ( .A1(G2090), .A2(G303), .ZN(n730) );
  XNOR2_X1 U812 ( .A(n730), .B(KEYINPUT96), .ZN(n731) );
  NAND2_X1 U813 ( .A1(n731), .A2(G8), .ZN(n733) );
  NAND2_X1 U814 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U815 ( .A1(n734), .A2(n737), .ZN(n739) );
  NOR2_X1 U816 ( .A1(G1981), .A2(G305), .ZN(n735) );
  XOR2_X1 U817 ( .A(n735), .B(KEYINPUT24), .Z(n736) );
  NOR2_X1 U818 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U819 ( .A1(n739), .A2(n738), .ZN(n740) );
  OR2_X1 U820 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U821 ( .A1(n743), .A2(n742), .ZN(n758) );
  NOR2_X1 U822 ( .A1(G1996), .A2(n866), .ZN(n932) );
  INV_X1 U823 ( .A(n744), .ZN(n747) );
  NOR2_X1 U824 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U825 ( .A1(n964), .A2(n879), .ZN(n940) );
  NOR2_X1 U826 ( .A1(n745), .A2(n940), .ZN(n746) );
  NOR2_X1 U827 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U828 ( .A1(n932), .A2(n748), .ZN(n749) );
  XOR2_X1 U829 ( .A(n749), .B(KEYINPUT97), .Z(n750) );
  XNOR2_X1 U830 ( .A(KEYINPUT39), .B(n750), .ZN(n751) );
  NAND2_X1 U831 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U832 ( .A1(n896), .A2(n753), .ZN(n924) );
  NAND2_X1 U833 ( .A1(n754), .A2(n924), .ZN(n756) );
  AND2_X1 U834 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U835 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U836 ( .A1(n760), .A2(n759), .ZN(n763) );
  XOR2_X1 U837 ( .A(KEYINPUT40), .B(KEYINPUT98), .Z(n761) );
  AND2_X1 U838 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U839 ( .A(G57), .ZN(G237) );
  INV_X1 U840 ( .A(G132), .ZN(G219) );
  INV_X1 U841 ( .A(G82), .ZN(G220) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U843 ( .A(n765), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U844 ( .A(G223), .ZN(n828) );
  NAND2_X1 U845 ( .A1(n828), .A2(G567), .ZN(n766) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  XNOR2_X1 U847 ( .A(G860), .B(KEYINPUT73), .ZN(n771) );
  OR2_X1 U848 ( .A1(n978), .A2(n771), .ZN(G153) );
  INV_X1 U849 ( .A(G171), .ZN(G301) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n768) );
  INV_X1 U851 ( .A(G868), .ZN(n811) );
  NAND2_X1 U852 ( .A1(n994), .A2(n811), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(G284) );
  NOR2_X1 U854 ( .A1(G286), .A2(n811), .ZN(n770) );
  NOR2_X1 U855 ( .A1(G868), .A2(G299), .ZN(n769) );
  NOR2_X1 U856 ( .A1(n770), .A2(n769), .ZN(G297) );
  NAND2_X1 U857 ( .A1(n771), .A2(G559), .ZN(n772) );
  INV_X1 U858 ( .A(n994), .ZN(n786) );
  NAND2_X1 U859 ( .A1(n772), .A2(n786), .ZN(n773) );
  XNOR2_X1 U860 ( .A(n773), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U861 ( .A1(G868), .A2(n978), .ZN(n776) );
  NAND2_X1 U862 ( .A1(G868), .A2(n786), .ZN(n774) );
  NOR2_X1 U863 ( .A1(G559), .A2(n774), .ZN(n775) );
  NOR2_X1 U864 ( .A1(n776), .A2(n775), .ZN(G282) );
  NAND2_X1 U865 ( .A1(G99), .A2(n888), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G111), .A2(n882), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n783) );
  NAND2_X1 U868 ( .A1(G123), .A2(n883), .ZN(n779) );
  XNOR2_X1 U869 ( .A(n779), .B(KEYINPUT18), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n886), .A2(G135), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n939) );
  XNOR2_X1 U873 ( .A(G2096), .B(n939), .ZN(n785) );
  INV_X1 U874 ( .A(G2100), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(G156) );
  NAND2_X1 U876 ( .A1(n786), .A2(G559), .ZN(n809) );
  XNOR2_X1 U877 ( .A(n978), .B(n809), .ZN(n787) );
  NOR2_X1 U878 ( .A1(n787), .A2(G860), .ZN(n799) );
  NAND2_X1 U879 ( .A1(G93), .A2(n788), .ZN(n791) );
  NAND2_X1 U880 ( .A1(G80), .A2(n789), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G55), .A2(n792), .ZN(n793) );
  XNOR2_X1 U883 ( .A(n793), .B(KEYINPUT76), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n794), .A2(G67), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n797) );
  OR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n812) );
  XOR2_X1 U887 ( .A(n799), .B(n812), .Z(G145) );
  XNOR2_X1 U888 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n801) );
  XNOR2_X1 U889 ( .A(G288), .B(KEYINPUT19), .ZN(n800) );
  XNOR2_X1 U890 ( .A(n801), .B(n800), .ZN(n802) );
  XNOR2_X1 U891 ( .A(G290), .B(n802), .ZN(n805) );
  XNOR2_X1 U892 ( .A(n803), .B(G166), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n805), .B(n804), .ZN(n806) );
  XOR2_X1 U894 ( .A(n812), .B(n806), .Z(n807) );
  XNOR2_X1 U895 ( .A(n807), .B(G305), .ZN(n808) );
  XNOR2_X1 U896 ( .A(n978), .B(n808), .ZN(n900) );
  XOR2_X1 U897 ( .A(n900), .B(n809), .Z(n810) );
  NOR2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n814) );
  NOR2_X1 U899 ( .A1(G868), .A2(n812), .ZN(n813) );
  NOR2_X1 U900 ( .A1(n814), .A2(n813), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n815) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n815), .Z(n816) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n817), .ZN(n818) );
  NAND2_X1 U905 ( .A1(n818), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(KEYINPUT82), .B(G44), .ZN(n819) );
  XNOR2_X1 U907 ( .A(n819), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U910 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U911 ( .A1(G96), .A2(n822), .ZN(n919) );
  NAND2_X1 U912 ( .A1(n919), .A2(G2106), .ZN(n826) );
  NAND2_X1 U913 ( .A1(G69), .A2(G120), .ZN(n823) );
  NOR2_X1 U914 ( .A1(G237), .A2(n823), .ZN(n824) );
  NAND2_X1 U915 ( .A1(G108), .A2(n824), .ZN(n920) );
  NAND2_X1 U916 ( .A1(n920), .A2(G567), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n834) );
  NAND2_X1 U918 ( .A1(G661), .A2(G483), .ZN(n827) );
  NOR2_X1 U919 ( .A1(n834), .A2(n827), .ZN(n831) );
  NAND2_X1 U920 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n828), .ZN(G217) );
  NAND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n829) );
  XOR2_X1 U923 ( .A(KEYINPUT100), .B(n829), .Z(n830) );
  NAND2_X1 U924 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U927 ( .A(KEYINPUT101), .B(n833), .Z(G188) );
  INV_X1 U928 ( .A(n834), .ZN(G319) );
  XOR2_X1 U929 ( .A(KEYINPUT104), .B(G1981), .Z(n836) );
  XNOR2_X1 U930 ( .A(G1966), .B(G1961), .ZN(n835) );
  XNOR2_X1 U931 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U932 ( .A(n837), .B(KEYINPUT41), .Z(n839) );
  XNOR2_X1 U933 ( .A(G1996), .B(G1991), .ZN(n838) );
  XNOR2_X1 U934 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U935 ( .A(G1986), .B(G1976), .Z(n841) );
  XNOR2_X1 U936 ( .A(G1956), .B(G1971), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U938 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U939 ( .A(KEYINPUT103), .B(G2474), .ZN(n844) );
  XNOR2_X1 U940 ( .A(n845), .B(n844), .ZN(G229) );
  XOR2_X1 U941 ( .A(G2096), .B(KEYINPUT43), .Z(n847) );
  XNOR2_X1 U942 ( .A(G2072), .B(G2678), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U944 ( .A(n848), .B(KEYINPUT102), .Z(n850) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2090), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U947 ( .A(KEYINPUT42), .B(G2100), .Z(n852) );
  XNOR2_X1 U948 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(G227) );
  NAND2_X1 U951 ( .A1(n886), .A2(G136), .ZN(n855) );
  XNOR2_X1 U952 ( .A(KEYINPUT106), .B(n855), .ZN(n859) );
  XOR2_X1 U953 ( .A(KEYINPUT44), .B(KEYINPUT105), .Z(n857) );
  NAND2_X1 U954 ( .A1(G124), .A2(n883), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n858) );
  NAND2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U957 ( .A1(G100), .A2(n888), .ZN(n861) );
  NAND2_X1 U958 ( .A1(G112), .A2(n882), .ZN(n860) );
  NAND2_X1 U959 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT107), .B(n862), .Z(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(G162) );
  XOR2_X1 U962 ( .A(G160), .B(n939), .Z(n865) );
  XNOR2_X1 U963 ( .A(n866), .B(n865), .ZN(n878) );
  XOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n876) );
  NAND2_X1 U965 ( .A1(G103), .A2(n888), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G139), .A2(n886), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U968 ( .A1(G115), .A2(n882), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G127), .A2(n883), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n871), .Z(n872) );
  XNOR2_X1 U972 ( .A(KEYINPUT110), .B(n872), .ZN(n873) );
  NOR2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n927) );
  XNOR2_X1 U974 ( .A(G164), .B(n927), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n881) );
  XNOR2_X1 U977 ( .A(n879), .B(G162), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n881), .B(n880), .ZN(n898) );
  NAND2_X1 U979 ( .A1(G118), .A2(n882), .ZN(n885) );
  NAND2_X1 U980 ( .A1(G130), .A2(n883), .ZN(n884) );
  NAND2_X1 U981 ( .A1(n885), .A2(n884), .ZN(n894) );
  NAND2_X1 U982 ( .A1(n886), .A2(G142), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n887), .B(KEYINPUT108), .ZN(n890) );
  NAND2_X1 U984 ( .A1(G106), .A2(n888), .ZN(n889) );
  NAND2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U986 ( .A(KEYINPUT45), .B(n891), .ZN(n892) );
  XNOR2_X1 U987 ( .A(KEYINPUT109), .B(n892), .ZN(n893) );
  NOR2_X1 U988 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U990 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U991 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U992 ( .A(G286), .B(n994), .ZN(n901) );
  XNOR2_X1 U993 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U994 ( .A(G171), .B(n902), .Z(n903) );
  NOR2_X1 U995 ( .A1(G37), .A2(n903), .ZN(n904) );
  XOR2_X1 U996 ( .A(KEYINPUT111), .B(n904), .Z(G397) );
  XOR2_X1 U997 ( .A(G2451), .B(G2430), .Z(n906) );
  XNOR2_X1 U998 ( .A(G2438), .B(G2443), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n906), .B(n905), .ZN(n912) );
  XOR2_X1 U1000 ( .A(G2435), .B(G2454), .Z(n908) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G1348), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1003 ( .A(G2446), .B(G2427), .Z(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1005 ( .A(n912), .B(n911), .Z(n913) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n913), .ZN(n921) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n921), .ZN(n916) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(G225) );
  XOR2_X1 U1013 ( .A(KEYINPUT112), .B(G225), .Z(G308) );
  INV_X1 U1015 ( .A(G120), .ZN(G236) );
  INV_X1 U1016 ( .A(G96), .ZN(G221) );
  INV_X1 U1017 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G325) );
  INV_X1 U1019 ( .A(G325), .ZN(G261) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  INV_X1 U1021 ( .A(n921), .ZN(G401) );
  XOR2_X1 U1022 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n949) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n938) );
  XNOR2_X1 U1025 ( .A(G164), .B(G2078), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n926), .B(KEYINPUT117), .ZN(n929) );
  XOR2_X1 U1027 ( .A(G2072), .B(n927), .Z(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(KEYINPUT50), .B(n930), .ZN(n936) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  XNOR2_X1 U1033 ( .A(KEYINPUT116), .B(n934), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n947) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(KEYINPUT114), .B(n941), .ZN(n944) );
  XOR2_X1 U1038 ( .A(G160), .B(G2084), .Z(n942) );
  XNOR2_X1 U1039 ( .A(KEYINPUT113), .B(n942), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n945), .B(KEYINPUT115), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(n949), .B(n948), .ZN(n951) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n952), .A2(G29), .ZN(n953) );
  XOR2_X1 U1047 ( .A(KEYINPUT119), .B(n953), .Z(n1034) );
  XNOR2_X1 U1048 ( .A(KEYINPUT121), .B(G2067), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(n954), .B(G26), .ZN(n963) );
  XNOR2_X1 U1050 ( .A(G2072), .B(G33), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G32), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(G28), .A2(n957), .ZN(n961) );
  XOR2_X1 U1054 ( .A(G27), .B(n958), .Z(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT122), .B(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G25), .B(n964), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1060 ( .A(KEYINPUT53), .B(n967), .Z(n970) );
  XOR2_X1 U1061 ( .A(KEYINPUT54), .B(G34), .Z(n968) );
  XNOR2_X1 U1062 ( .A(G2084), .B(n968), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(KEYINPUT120), .B(G2090), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(G35), .B(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(KEYINPUT55), .B(n974), .ZN(n976) );
  INV_X1 U1068 ( .A(G29), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n977), .A2(G11), .ZN(n1032) );
  XNOR2_X1 U1071 ( .A(G16), .B(KEYINPUT56), .ZN(n1003) );
  XNOR2_X1 U1072 ( .A(n1004), .B(n978), .ZN(n1001) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(n981), .B(KEYINPUT123), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT57), .B(n982), .ZN(n999) );
  NAND2_X1 U1077 ( .A1(G1971), .A2(G303), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G1956), .B(G299), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(KEYINPUT124), .B(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G171), .B(G1961), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G1348), .B(n994), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(KEYINPUT125), .B(n997), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1030) );
  INV_X1 U1092 ( .A(G16), .ZN(n1028) );
  XNOR2_X1 U1093 ( .A(G19), .B(n1004), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G20), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT59), .B(G1348), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(KEYINPUT60), .B(n1012), .ZN(n1024) );
  XOR2_X1 U1102 ( .A(G1966), .B(G21), .Z(n1015) );
  XNOR2_X1 U1103 ( .A(n1013), .B(G5), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(G1971), .B(G22), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(G23), .B(G1976), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XOR2_X1 U1108 ( .A(G1986), .B(G24), .Z(n1018) );
  NAND2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1110 ( .A(KEYINPUT58), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(n1025), .B(KEYINPUT126), .ZN(n1026) );
  XOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1026), .Z(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1119 ( .A(n1035), .B(KEYINPUT127), .ZN(n1036) );
  XNOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1036), .ZN(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

