//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  INV_X1    g005(.A(G131), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G137), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT65), .B1(new_n188), .B2(G137), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n190), .A3(G134), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(new_n193), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G131), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT64), .A2(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT64), .A2(G143), .ZN(new_n201));
  OAI21_X1  g015(.A(G146), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n202), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n203), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT64), .A2(G143), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n203), .A2(G146), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n213), .A2(new_n214), .B1(G128), .B2(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n194), .B(new_n199), .C1(new_n208), .C2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n189), .A2(new_n193), .A3(new_n191), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n194), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT64), .B(G143), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n204), .B1(new_n221), .B2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n213), .A2(new_n214), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n220), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G116), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT2), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G113), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(KEYINPUT66), .A3(new_n237), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n239), .ZN(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n240), .A2(new_n244), .A3(KEYINPUT67), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT67), .B1(new_n240), .B2(new_n244), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n217), .B(new_n230), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n240), .A2(new_n244), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n217), .B2(new_n230), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT28), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT28), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n217), .A2(new_n230), .A3(new_n254), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n245), .A2(new_n246), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n254), .B1(new_n217), .B2(new_n230), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(G101), .ZN(new_n261));
  INV_X1    g075(.A(G237), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n261), .B(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n252), .A2(new_n259), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n265), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n217), .A2(new_n230), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT30), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n217), .A2(new_n230), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n250), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n267), .B1(new_n272), .B2(new_n248), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n266), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT70), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n245), .A2(new_n246), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n268), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n253), .B1(new_n279), .B2(new_n247), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT71), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n267), .A2(new_n274), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n281), .B(new_n282), .C1(new_n283), .C2(new_n280), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n266), .A2(new_n273), .A3(new_n285), .A4(new_n274), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n276), .A2(new_n277), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G472), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n265), .B1(new_n252), .B2(new_n259), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n247), .A2(new_n291), .A3(new_n265), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n291), .B1(new_n247), .B2(new_n265), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n217), .A2(new_n230), .A3(new_n270), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n270), .B1(new_n217), .B2(new_n230), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n249), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT31), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n265), .B1(new_n268), .B2(new_n278), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT68), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n247), .A2(new_n291), .A3(new_n265), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n297), .A3(KEYINPUT31), .A4(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n290), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n300), .A2(new_n297), .A3(new_n301), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT31), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n289), .B1(new_n310), .B2(new_n302), .ZN(new_n311));
  INV_X1    g125(.A(new_n306), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT32), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n288), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT72), .ZN(new_n316));
  XNOR2_X1  g130(.A(G125), .B(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT16), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n318), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G146), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n318), .B(new_n211), .C1(new_n323), .C2(new_n325), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT23), .B1(new_n206), .B2(G119), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT73), .B1(new_n206), .B2(G119), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G119), .B(G128), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT24), .B(G110), .Z(new_n334));
  AOI22_X1  g148(.A1(new_n332), .A2(G110), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  OAI22_X1  g150(.A1(new_n332), .A2(G110), .B1(new_n333), .B2(new_n334), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n317), .A2(new_n211), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n327), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(G137), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n343));
  XOR2_X1   g157(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n336), .A3(new_n339), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n277), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT25), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G217), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(G234), .B2(new_n277), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT25), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n352), .A2(KEYINPUT77), .A3(new_n354), .A4(new_n355), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n354), .A2(G902), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n360), .B(KEYINPUT78), .Z(new_n361));
  NAND3_X1  g175(.A1(new_n346), .A2(new_n347), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT72), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n288), .A2(new_n314), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n316), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n329), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n200), .A2(new_n201), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n262), .A2(new_n263), .A3(G214), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n203), .A2(new_n262), .A3(new_n263), .A4(G214), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n371), .A2(KEYINPUT17), .A3(G131), .A4(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT91), .ZN(new_n374));
  INV_X1    g188(.A(G214), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n375), .A2(G237), .A3(G953), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n372), .B1(new_n221), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n192), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT17), .ZN(new_n379));
  OAI211_X1 g193(.A(G131), .B(new_n372), .C1(new_n221), .C2(new_n376), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n368), .B(new_n374), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(G113), .B(G122), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT18), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n377), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n317), .B(new_n211), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n371), .A2(KEYINPUT18), .A3(G131), .A4(new_n372), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .A4(new_n378), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n388), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n317), .B(KEYINPUT19), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n211), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n378), .A2(new_n380), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n327), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n388), .B1(new_n398), .B2(new_n393), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(KEYINPUT90), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(KEYINPUT90), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(G475), .A2(G902), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n403), .B(KEYINPUT93), .Z(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT20), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n385), .A2(new_n388), .A3(new_n393), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n388), .B1(new_n385), .B2(new_n393), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n277), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G475), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n402), .A2(KEYINPUT20), .A3(new_n404), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n407), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n263), .A2(G952), .ZN(new_n414));
  NAND2_X1  g228(.A1(G234), .A2(G237), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XOR2_X1   g230(.A(KEYINPUT21), .B(G898), .Z(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(G902), .A3(G953), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G478), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(KEYINPUT15), .ZN(new_n421));
  XNOR2_X1  g235(.A(G116), .B(G122), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G107), .ZN(new_n424));
  INV_X1    g238(.A(G107), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n203), .A2(G128), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(new_n221), .B2(G128), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n424), .A2(new_n426), .B1(new_n428), .B2(new_n188), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n221), .A2(G128), .ZN(new_n430));
  INV_X1    g244(.A(new_n427), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(KEYINPUT13), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT13), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n221), .A2(new_n433), .A3(G128), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(G134), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n233), .A2(KEYINPUT14), .A3(G122), .ZN(new_n437));
  OAI211_X1 g251(.A(G107), .B(new_n437), .C1(new_n423), .C2(KEYINPUT14), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n428), .A2(new_n188), .ZN(new_n439));
  AOI211_X1 g253(.A(G134), .B(new_n427), .C1(new_n221), .C2(G128), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n426), .B(new_n438), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT9), .B(G234), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT79), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n444), .A2(new_n353), .A3(G953), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n436), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n445), .B1(new_n436), .B2(new_n441), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n277), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n421), .B1(new_n448), .B2(KEYINPUT94), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(KEYINPUT94), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT94), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n451), .B(new_n277), .C1(new_n446), .C2(new_n447), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n449), .B1(new_n453), .B2(new_n421), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n413), .A2(KEYINPUT95), .A3(new_n419), .A4(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT95), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n407), .A2(new_n454), .A3(new_n411), .A4(new_n412), .ZN(new_n457));
  INV_X1    g271(.A(new_n419), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G214), .B1(G237), .B2(G902), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n463));
  INV_X1    g277(.A(new_n225), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n226), .A2(new_n228), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n463), .B(G125), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n222), .A2(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT86), .B1(new_n467), .B2(new_n321), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n208), .A2(new_n216), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n321), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT89), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n263), .A2(G224), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT7), .A4(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n466), .A2(new_n468), .A3(new_n470), .A4(new_n473), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT89), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT3), .B1(new_n387), .B2(G107), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT3), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n425), .A3(G104), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n387), .A2(G107), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G101), .ZN(new_n484));
  INV_X1    g298(.A(G101), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n479), .A2(new_n481), .A3(new_n485), .A4(new_n482), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(KEYINPUT4), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT80), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n487), .B(new_n488), .C1(KEYINPUT4), .C2(new_n484), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n484), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n486), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n250), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT84), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n425), .A2(G104), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n387), .A2(G107), .ZN(new_n495));
  OAI21_X1  g309(.A(G101), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n486), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n232), .A2(new_n234), .A3(KEYINPUT5), .ZN(new_n498));
  OR3_X1    g312(.A1(new_n233), .A2(KEYINPUT5), .A3(G119), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(G113), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT83), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n241), .A2(new_n242), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT83), .A4(G113), .ZN(new_n504));
  AND4_X1   g318(.A1(new_n497), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n491), .A2(new_n493), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n486), .A2(new_n496), .ZN(new_n507));
  AND4_X1   g321(.A1(new_n507), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n493), .A2(KEYINPUT8), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n493), .A2(KEYINPUT8), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n503), .B2(new_n500), .ZN(new_n511));
  NOR4_X1   g325(.A1(new_n508), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT88), .B(KEYINPUT7), .Z(new_n514));
  AOI22_X1  g328(.A1(new_n513), .A2(new_n470), .B1(new_n473), .B2(new_n514), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n506), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n478), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n471), .B(new_n473), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n484), .A2(KEYINPUT4), .A3(new_n486), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n488), .B1(new_n484), .B2(KEYINPUT4), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n490), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n505), .B1(new_n522), .B2(new_n249), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n493), .A2(KEYINPUT85), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n524), .ZN(new_n526));
  OAI211_X1 g340(.A(KEYINPUT6), .B(new_n526), .C1(new_n491), .C2(new_n505), .ZN(new_n527));
  INV_X1    g341(.A(new_n493), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT87), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n518), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n518), .B2(new_n530), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n517), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G210), .B1(G237), .B2(G902), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n517), .B(new_n535), .C1(new_n532), .C2(new_n533), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n462), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G469), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT81), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n497), .A2(KEYINPUT10), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n469), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT10), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n507), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n545), .B(KEYINPUT81), .C1(new_n216), .C2(new_n208), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n522), .A2(new_n467), .ZN(new_n548));
  INV_X1    g362(.A(new_n220), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n206), .B1(new_n213), .B2(KEYINPUT1), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(new_n222), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n497), .B1(new_n551), .B2(new_n208), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n544), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G140), .ZN(new_n555));
  INV_X1    g369(.A(G227), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(G953), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n555), .B(new_n557), .Z(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n469), .A2(new_n507), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT12), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n549), .B2(KEYINPUT82), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n561), .A2(new_n220), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n563), .B1(new_n561), .B2(new_n220), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n547), .A2(new_n548), .A3(new_n553), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n220), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n558), .B1(new_n569), .B2(new_n554), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n540), .B(new_n277), .C1(new_n567), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(G469), .A2(G902), .ZN(new_n572));
  INV_X1    g386(.A(new_n558), .ZN(new_n573));
  INV_X1    g387(.A(new_n554), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n573), .B1(new_n566), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n569), .A2(new_n554), .A3(new_n558), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(G469), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(G221), .B1(new_n444), .B2(G902), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n460), .A2(new_n539), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n367), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(new_n485), .ZN(G3));
  NAND2_X1  g398(.A1(new_n537), .A2(new_n538), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n407), .A2(new_n411), .A3(new_n412), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n436), .A2(new_n441), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT33), .B1(new_n587), .B2(KEYINPUT96), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n446), .A2(new_n447), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(G478), .A3(new_n277), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n448), .A2(new_n420), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n585), .A2(new_n419), .A3(new_n596), .A4(new_n461), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT98), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n539), .A2(new_n599), .A3(new_n419), .A4(new_n596), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G472), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n304), .B2(new_n277), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n304), .B2(new_n306), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n364), .A2(new_n581), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(new_n387), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n607), .B(new_n609), .ZN(G6));
  INV_X1    g424(.A(new_n454), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n611), .A2(new_n407), .A3(new_n411), .A4(new_n412), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT100), .B1(new_n612), .B2(new_n458), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n413), .A2(new_n614), .A3(new_n419), .A4(new_n611), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n539), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n539), .A2(new_n613), .A3(KEYINPUT101), .A4(new_n615), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n606), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT102), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n621), .B(new_n623), .ZN(G9));
  NAND4_X1  g438(.A1(new_n460), .A2(new_n539), .A3(new_n581), .A4(new_n605), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n345), .A2(KEYINPUT36), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n340), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n361), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n358), .A2(new_n359), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT37), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G110), .ZN(G12));
  AND3_X1   g447(.A1(new_n288), .A2(new_n314), .A3(new_n365), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n365), .B1(new_n288), .B2(new_n314), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n539), .A2(new_n581), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n418), .A2(G900), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n416), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n612), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n636), .A2(new_n637), .A3(new_n629), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G128), .ZN(G30));
  XOR2_X1   g457(.A(new_n639), .B(KEYINPUT39), .Z(new_n644));
  NOR2_X1   g458(.A1(new_n580), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n645), .A2(KEYINPUT40), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(KEYINPUT40), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n462), .B(new_n629), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n585), .B(KEYINPUT38), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n413), .A2(new_n454), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n265), .B1(new_n279), .B2(new_n247), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n297), .B2(new_n294), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n652), .B2(G902), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n314), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n648), .A2(new_n649), .A3(new_n650), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n369), .ZN(G45));
  NAND2_X1  g470(.A1(new_n596), .A2(new_n639), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n636), .A2(new_n637), .A3(new_n629), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G146), .ZN(G48));
  INV_X1    g474(.A(new_n570), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n559), .A2(new_n566), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n540), .B1(new_n663), .B2(new_n277), .ZN(new_n664));
  INV_X1    g478(.A(new_n571), .ZN(new_n665));
  INV_X1    g479(.A(new_n579), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n316), .A2(new_n364), .A3(new_n366), .A4(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n601), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT41), .B(G113), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G15));
  AOI21_X1  g485(.A(new_n668), .B1(new_n618), .B2(new_n619), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT103), .B(G116), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G18));
  AND2_X1   g488(.A1(new_n455), .A2(new_n459), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n539), .A2(new_n667), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n634), .A2(new_n635), .A3(new_n630), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n231), .ZN(G21));
  NAND2_X1  g494(.A1(new_n585), .A2(new_n461), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n664), .A2(new_n665), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n579), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n306), .B(KEYINPUT104), .Z(new_n685));
  OAI21_X1  g499(.A(new_n281), .B1(new_n283), .B2(new_n280), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n686), .A2(new_n267), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n298), .A2(new_n303), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n604), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n363), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n684), .A2(new_n419), .A3(new_n650), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G122), .ZN(G24));
  NOR2_X1   g508(.A1(new_n630), .A2(new_n640), .ZN(new_n695));
  INV_X1    g509(.A(new_n596), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n691), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n684), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n537), .A2(new_n461), .A3(new_n538), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n580), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(new_n316), .A3(new_n364), .A4(new_n366), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n700), .B1(new_n703), .B2(new_n657), .ZN(new_n704));
  AOI22_X1  g518(.A1(G472), .A2(new_n287), .B1(new_n307), .B2(new_n313), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT105), .B1(new_n705), .B2(new_n363), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n364), .A2(new_n315), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n657), .A2(new_n701), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(KEYINPUT42), .A3(new_n581), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G131), .ZN(G33));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n641), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n703), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n641), .A2(new_n714), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G134), .ZN(G36));
  AND2_X1   g533(.A1(new_n575), .A2(new_n576), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n720), .A2(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(KEYINPUT45), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(G469), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n572), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n665), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(KEYINPUT46), .A3(new_n572), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n666), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n644), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n413), .A2(new_n595), .ZN(new_n731));
  NAND2_X1  g545(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n734));
  OAI21_X1  g548(.A(new_n733), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n605), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n629), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n701), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n730), .B(new_n739), .C1(new_n738), .C2(new_n737), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G137), .ZN(G39));
  OR2_X1    g555(.A1(new_n728), .A2(KEYINPUT47), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n728), .A2(KEYINPUT47), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n636), .A2(new_n364), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n710), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G140), .ZN(G42));
  XNOR2_X1  g561(.A(new_n682), .B(KEYINPUT108), .ZN(new_n748));
  NOR2_X1   g562(.A1(KEYINPUT109), .A2(KEYINPUT49), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n363), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n649), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n750), .A2(new_n579), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n748), .A2(new_n749), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n731), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n654), .B1(KEYINPUT109), .B2(KEYINPUT49), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n461), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n416), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n735), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n735), .A2(KEYINPUT114), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n762), .A2(new_n692), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n684), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n667), .A2(KEYINPUT115), .A3(new_n462), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n667), .A2(new_n462), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n649), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n763), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT50), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n763), .A2(new_n772), .A3(new_n766), .A4(new_n769), .ZN(new_n773));
  INV_X1    g587(.A(new_n691), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n683), .A2(new_n701), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n762), .A2(new_n629), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n654), .A2(new_n416), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n364), .A3(new_n777), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n778), .A2(new_n586), .A3(new_n595), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n771), .A2(new_n773), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n748), .A2(new_n666), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n742), .A2(new_n743), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n701), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n763), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n765), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n773), .A2(new_n776), .A3(new_n779), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT51), .A3(new_n784), .A4(new_n771), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n778), .A2(new_n696), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n786), .A2(new_n788), .A3(new_n414), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n762), .A2(new_n709), .A3(new_n775), .ZN(new_n791));
  XNOR2_X1  g605(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  OAI22_X1  g608(.A1(new_n367), .A2(new_n582), .B1(new_n625), .B2(new_n630), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n681), .A2(new_n458), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n696), .A2(new_n612), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n796), .A2(new_n606), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n634), .A2(new_n635), .A3(new_n457), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n695), .B(new_n702), .C1(new_n800), .C2(new_n697), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n799), .A2(new_n712), .A3(new_n718), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n693), .B1(new_n601), .B2(new_n668), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n668), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n620), .A2(new_n805), .B1(new_n678), .B2(new_n677), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g622(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n809));
  NOR2_X1   g623(.A1(new_n629), .A2(new_n640), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n637), .A2(new_n650), .A3(new_n654), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n642), .A2(new_n659), .A3(new_n698), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT110), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n678), .B(new_n637), .C1(new_n641), .C2(new_n658), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT110), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n815), .A2(new_n816), .A3(new_n698), .A4(new_n811), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n814), .B1(new_n813), .B2(new_n817), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n808), .B(new_n809), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n812), .A2(new_n814), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT53), .B1(new_n824), .B2(new_n808), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT54), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n804), .B2(new_n806), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n802), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n803), .A2(new_n672), .A3(new_n679), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(new_n827), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n704), .A2(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n831), .A2(new_n835), .A3(new_n799), .A4(new_n801), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n813), .A2(new_n817), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n836), .B1(new_n838), .B2(new_n822), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n833), .B(new_n834), .C1(new_n839), .C2(new_n809), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n826), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT113), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n826), .A2(new_n843), .A3(new_n840), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n764), .A2(new_n794), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(G952), .A2(G953), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n756), .B1(new_n845), .B2(new_n846), .ZN(G75));
  OAI21_X1  g661(.A(new_n833), .B1(new_n839), .B2(new_n809), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n277), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(G210), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n530), .B(KEYINPUT117), .Z(new_n853));
  XNOR2_X1  g667(.A(new_n518), .B(KEYINPUT55), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n856), .B2(KEYINPUT56), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n851), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n857), .B1(new_n851), .B2(new_n852), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n263), .A2(G952), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(G51));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n572), .B(KEYINPUT57), .Z(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n865), .B2(new_n840), .ZN(new_n866));
  INV_X1    g680(.A(new_n663), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n840), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n808), .B1(new_n818), .B2(new_n819), .ZN(new_n870));
  INV_X1    g684(.A(new_n809), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n834), .B1(new_n872), .B2(new_n833), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n863), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(KEYINPUT119), .A3(new_n663), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n849), .A2(new_n277), .A3(new_n723), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n868), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n860), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(G54));
  NAND3_X1  g693(.A1(new_n850), .A2(KEYINPUT58), .A3(G475), .ZN(new_n880));
  INV_X1    g694(.A(new_n402), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(new_n860), .ZN(G60));
  XOR2_X1   g698(.A(new_n590), .B(KEYINPUT120), .Z(new_n885));
  NAND2_X1  g699(.A1(G478), .A2(G902), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT59), .Z(new_n887));
  AOI211_X1 g701(.A(new_n885), .B(new_n887), .C1(new_n865), .C2(new_n840), .ZN(new_n888));
  INV_X1    g702(.A(new_n887), .ZN(new_n889));
  INV_X1    g703(.A(new_n844), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n843), .B1(new_n826), .B2(new_n840), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n860), .B(new_n888), .C1(new_n892), .C2(new_n885), .ZN(G63));
  NAND2_X1  g707(.A1(G217), .A2(G902), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT60), .ZN(new_n895));
  INV_X1    g709(.A(new_n347), .ZN(new_n896));
  INV_X1    g710(.A(new_n346), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n849), .A2(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n895), .B1(new_n872), .B2(new_n833), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n860), .B1(new_n899), .B2(new_n627), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n900), .B2(KEYINPUT121), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n901), .B(new_n903), .ZN(G66));
  AOI21_X1  g718(.A(new_n263), .B1(new_n417), .B2(G224), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n831), .A2(new_n799), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n906), .B2(new_n263), .ZN(new_n907));
  INV_X1    g721(.A(G898), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n853), .B1(new_n908), .B2(G953), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n907), .B(new_n909), .ZN(G69));
  AOI21_X1  g724(.A(new_n263), .B1(G227), .B2(G900), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT124), .Z(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT126), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n263), .A2(G900), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n815), .A2(new_n698), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n746), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n730), .A2(new_n539), .A3(new_n650), .A4(new_n709), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n835), .B(KEYINPUT125), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n916), .A2(new_n740), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n919), .B2(new_n263), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n295), .A2(new_n296), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n395), .ZN(new_n922));
  INV_X1    g736(.A(new_n367), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n645), .A3(new_n783), .A4(new_n797), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n746), .A2(new_n740), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n655), .A2(new_n915), .A3(new_n926), .ZN(new_n927));
  OR3_X1    g741(.A1(new_n927), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n925), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n263), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n922), .B(KEYINPUT122), .ZN(new_n932));
  OAI221_X1 g746(.A(new_n913), .B1(new_n920), .B2(new_n922), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n912), .A2(KEYINPUT126), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G72));
  NAND2_X1  g749(.A1(G472), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT63), .Z(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n930), .B2(new_n906), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n938), .B(new_n265), .C1(new_n248), .C2(new_n272), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n919), .B2(new_n906), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n940), .A2(new_n247), .A3(new_n267), .A4(new_n297), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n941), .A3(new_n878), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n821), .A2(new_n825), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n308), .B2(new_n273), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n937), .B2(new_n944), .ZN(G57));
endmodule


