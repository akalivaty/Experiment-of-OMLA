

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  XNOR2_X1 U321 ( .A(n430), .B(n402), .ZN(n403) );
  XNOR2_X1 U322 ( .A(n401), .B(n400), .ZN(n402) );
  NOR2_X1 U323 ( .A1(n465), .A2(n464), .ZN(n467) );
  XNOR2_X1 U324 ( .A(n445), .B(n444), .ZN(n524) );
  XOR2_X1 U325 ( .A(n406), .B(n405), .Z(n512) );
  AND2_X1 U326 ( .A1(n524), .A2(n512), .ZN(n453) );
  XNOR2_X1 U327 ( .A(KEYINPUT25), .B(KEYINPUT102), .ZN(n455) );
  XNOR2_X1 U328 ( .A(n456), .B(n455), .ZN(n457) );
  INV_X1 U329 ( .A(G134GAT), .ZN(n294) );
  XNOR2_X1 U330 ( .A(n295), .B(n294), .ZN(n296) );
  INV_X1 U331 ( .A(KEYINPUT103), .ZN(n466) );
  XNOR2_X1 U332 ( .A(n364), .B(n296), .ZN(n297) );
  XNOR2_X1 U333 ( .A(n467), .B(n466), .ZN(n479) );
  INV_X1 U334 ( .A(G190GAT), .ZN(n447) );
  XOR2_X1 U335 ( .A(n552), .B(KEYINPUT75), .Z(n536) );
  XOR2_X1 U336 ( .A(KEYINPUT38), .B(n484), .Z(n493) );
  XNOR2_X1 U337 ( .A(n447), .B(KEYINPUT58), .ZN(n448) );
  XNOR2_X1 U338 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n291) );
  XOR2_X1 U340 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  XNOR2_X1 U341 ( .A(G36GAT), .B(G190GAT), .ZN(n289) );
  XNOR2_X1 U342 ( .A(n289), .B(G218GAT), .ZN(n401) );
  XNOR2_X1 U343 ( .A(n422), .B(n401), .ZN(n290) );
  XNOR2_X1 U344 ( .A(n291), .B(n290), .ZN(n298) );
  XOR2_X1 U345 ( .A(G29GAT), .B(G43GAT), .Z(n293) );
  XNOR2_X1 U346 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n292) );
  XNOR2_X1 U347 ( .A(n293), .B(n292), .ZN(n364) );
  NAND2_X1 U348 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U349 ( .A(n298), .B(n297), .Z(n306) );
  XOR2_X1 U350 ( .A(KEYINPUT70), .B(G92GAT), .Z(n300) );
  XNOR2_X1 U351 ( .A(G99GAT), .B(G85GAT), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U353 ( .A(G106GAT), .B(n301), .Z(n333) );
  XOR2_X1 U354 ( .A(KEYINPUT74), .B(KEYINPUT10), .Z(n303) );
  XNOR2_X1 U355 ( .A(KEYINPUT64), .B(KEYINPUT65), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n333), .B(n304), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n552) );
  XNOR2_X1 U359 ( .A(G127GAT), .B(G134GAT), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n307), .B(KEYINPUT81), .ZN(n308) );
  XOR2_X1 U361 ( .A(n308), .B(KEYINPUT0), .Z(n310) );
  XNOR2_X1 U362 ( .A(G113GAT), .B(G120GAT), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n445) );
  XOR2_X1 U364 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n312) );
  NAND2_X1 U365 ( .A1(G225GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U367 ( .A(KEYINPUT95), .B(n313), .ZN(n328) );
  XOR2_X1 U368 ( .A(KEYINPUT6), .B(G57GAT), .Z(n315) );
  XNOR2_X1 U369 ( .A(G1GAT), .B(G155GAT), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U371 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n317) );
  XNOR2_X1 U372 ( .A(KEYINPUT1), .B(KEYINPUT92), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U374 ( .A(n319), .B(n318), .Z(n326) );
  XOR2_X1 U375 ( .A(KEYINPUT88), .B(KEYINPUT3), .Z(n321) );
  XNOR2_X1 U376 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n426) );
  XOR2_X1 U378 ( .A(G85GAT), .B(G148GAT), .Z(n323) );
  XNOR2_X1 U379 ( .A(G29GAT), .B(G162GAT), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n426), .B(n324), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n445), .B(n329), .ZN(n509) );
  INV_X1 U385 ( .A(KEYINPUT54), .ZN(n409) );
  XOR2_X1 U386 ( .A(KEYINPUT69), .B(KEYINPUT33), .Z(n331) );
  XNOR2_X1 U387 ( .A(G120GAT), .B(KEYINPUT72), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n344) );
  XOR2_X1 U390 ( .A(KEYINPUT68), .B(KEYINPUT13), .Z(n335) );
  XNOR2_X1 U391 ( .A(G71GAT), .B(G57GAT), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n351) );
  XOR2_X1 U393 ( .A(G148GAT), .B(G78GAT), .Z(n418) );
  XOR2_X1 U394 ( .A(n351), .B(n418), .Z(n337) );
  NAND2_X1 U395 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U397 ( .A(n338), .B(KEYINPUT31), .Z(n342) );
  XOR2_X1 U398 ( .A(G64GAT), .B(KEYINPUT71), .Z(n340) );
  XNOR2_X1 U399 ( .A(G176GAT), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n390) );
  XNOR2_X1 U401 ( .A(n390), .B(KEYINPUT32), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n569) );
  XOR2_X1 U404 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n346) );
  XNOR2_X1 U405 ( .A(KEYINPUT78), .B(KEYINPUT12), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n361) );
  XOR2_X1 U407 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n348) );
  NAND2_X1 U408 ( .A1(G231GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U410 ( .A(n349), .B(KEYINPUT77), .Z(n353) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(G183GAT), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n350), .B(KEYINPUT76), .ZN(n389) );
  XNOR2_X1 U413 ( .A(n389), .B(n351), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U415 ( .A(G64GAT), .B(G78GAT), .Z(n355) );
  XNOR2_X1 U416 ( .A(G127GAT), .B(G211GAT), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U418 ( .A(n357), .B(n356), .Z(n359) );
  XOR2_X1 U419 ( .A(G15GAT), .B(G1GAT), .Z(n363) );
  XOR2_X1 U420 ( .A(G22GAT), .B(G155GAT), .Z(n417) );
  XNOR2_X1 U421 ( .A(n363), .B(n417), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U423 ( .A(n361), .B(n360), .Z(n468) );
  INV_X1 U424 ( .A(n468), .ZN(n573) );
  XNOR2_X1 U425 ( .A(KEYINPUT36), .B(n536), .ZN(n578) );
  NOR2_X1 U426 ( .A1(n573), .A2(n578), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n362), .B(KEYINPUT45), .ZN(n379) );
  XOR2_X1 U428 ( .A(n364), .B(n363), .Z(n366) );
  NAND2_X1 U429 ( .A1(G229GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U431 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n368) );
  XNOR2_X1 U432 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U434 ( .A(n370), .B(n369), .Z(n378) );
  XOR2_X1 U435 ( .A(G113GAT), .B(G36GAT), .Z(n372) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(G50GAT), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U438 ( .A(G8GAT), .B(G197GAT), .Z(n374) );
  XNOR2_X1 U439 ( .A(G141GAT), .B(G22GAT), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U442 ( .A(n378), .B(n377), .Z(n527) );
  INV_X1 U443 ( .A(n527), .ZN(n565) );
  NAND2_X1 U444 ( .A1(n379), .A2(n565), .ZN(n380) );
  NOR2_X1 U445 ( .A1(n569), .A2(n380), .ZN(n381) );
  XOR2_X1 U446 ( .A(KEYINPUT117), .B(n381), .Z(n387) );
  NAND2_X1 U447 ( .A1(n552), .A2(n573), .ZN(n384) );
  XNOR2_X1 U448 ( .A(KEYINPUT41), .B(n569), .ZN(n543) );
  NOR2_X1 U449 ( .A1(n565), .A2(n543), .ZN(n382) );
  XNOR2_X1 U450 ( .A(n382), .B(KEYINPUT46), .ZN(n383) );
  NOR2_X1 U451 ( .A1(n384), .A2(n383), .ZN(n385) );
  XOR2_X1 U452 ( .A(KEYINPUT47), .B(n385), .Z(n386) );
  NOR2_X1 U453 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n388), .B(KEYINPUT48), .ZN(n522) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n406) );
  XOR2_X1 U456 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n392) );
  XNOR2_X1 U457 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U459 ( .A(G169GAT), .B(n393), .ZN(n439) );
  XOR2_X1 U460 ( .A(KEYINPUT96), .B(G92GAT), .Z(n395) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U463 ( .A(n439), .B(n396), .Z(n404) );
  XOR2_X1 U464 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n398) );
  XNOR2_X1 U465 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U467 ( .A(G197GAT), .B(n399), .Z(n430) );
  XOR2_X1 U468 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n400) );
  XNOR2_X1 U469 ( .A(n404), .B(n403), .ZN(n405) );
  INV_X1 U470 ( .A(n512), .ZN(n407) );
  NOR2_X1 U471 ( .A1(n522), .A2(n407), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n410) );
  NOR2_X1 U473 ( .A1(n509), .A2(n410), .ZN(n564) );
  XOR2_X1 U474 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n412) );
  XNOR2_X1 U475 ( .A(G218GAT), .B(G106GAT), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U477 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n414) );
  XNOR2_X1 U478 ( .A(KEYINPUT91), .B(KEYINPUT24), .ZN(n413) );
  XNOR2_X1 U479 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U480 ( .A(n416), .B(n415), .Z(n424) );
  XOR2_X1 U481 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U486 ( .A(n425), .B(G204GAT), .Z(n428) );
  XNOR2_X1 U487 ( .A(n426), .B(KEYINPUT89), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n460) );
  NAND2_X1 U490 ( .A1(n564), .A2(n460), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n431), .B(KEYINPUT55), .ZN(n446) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XOR2_X1 U493 ( .A(KEYINPUT84), .B(G176GAT), .Z(n433) );
  XNOR2_X1 U494 ( .A(G190GAT), .B(G71GAT), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U496 ( .A(G43GAT), .B(G99GAT), .Z(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U500 ( .A(G183GAT), .B(KEYINPUT82), .Z(n441) );
  XNOR2_X1 U501 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n444) );
  NAND2_X1 U504 ( .A1(n446), .A2(n524), .ZN(n561) );
  NOR2_X1 U505 ( .A1(n536), .A2(n561), .ZN(n449) );
  NOR2_X1 U506 ( .A1(n565), .A2(n569), .ZN(n450) );
  XOR2_X1 U507 ( .A(KEYINPUT73), .B(n450), .Z(n483) );
  NOR2_X1 U508 ( .A1(n524), .A2(n460), .ZN(n451) );
  XOR2_X1 U509 ( .A(KEYINPUT26), .B(n451), .Z(n540) );
  INV_X1 U510 ( .A(n540), .ZN(n563) );
  XNOR2_X1 U511 ( .A(n512), .B(KEYINPUT27), .ZN(n461) );
  AND2_X1 U512 ( .A1(n563), .A2(n461), .ZN(n452) );
  XNOR2_X1 U513 ( .A(KEYINPUT100), .B(n452), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n453), .B(KEYINPUT101), .ZN(n454) );
  NAND2_X1 U515 ( .A1(n454), .A2(n460), .ZN(n456) );
  NOR2_X1 U516 ( .A1(n458), .A2(n457), .ZN(n459) );
  NOR2_X1 U517 ( .A1(n509), .A2(n459), .ZN(n465) );
  XOR2_X1 U518 ( .A(KEYINPUT28), .B(n460), .Z(n516) );
  INV_X1 U519 ( .A(n516), .ZN(n525) );
  NAND2_X1 U520 ( .A1(n461), .A2(n509), .ZN(n521) );
  NOR2_X1 U521 ( .A1(n524), .A2(n521), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n525), .A2(n462), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n463), .B(KEYINPUT99), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n468), .A2(n536), .ZN(n469) );
  XNOR2_X1 U525 ( .A(KEYINPUT16), .B(n469), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n479), .A2(n470), .ZN(n497) );
  AND2_X1 U527 ( .A1(n483), .A2(n497), .ZN(n476) );
  NAND2_X1 U528 ( .A1(n509), .A2(n476), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT34), .ZN(n472) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n472), .ZN(G1324GAT) );
  NAND2_X1 U531 ( .A1(n512), .A2(n476), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U534 ( .A1(n476), .A2(n524), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  NAND2_X1 U536 ( .A1(n516), .A2(n476), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(KEYINPUT104), .ZN(n478) );
  XNOR2_X1 U538 ( .A(G22GAT), .B(n478), .ZN(G1327GAT) );
  XOR2_X1 U539 ( .A(G29GAT), .B(KEYINPUT39), .Z(n486) );
  NOR2_X1 U540 ( .A1(n479), .A2(n578), .ZN(n480) );
  NAND2_X1 U541 ( .A1(n480), .A2(n573), .ZN(n482) );
  XOR2_X1 U542 ( .A(KEYINPUT105), .B(KEYINPUT37), .Z(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(n508) );
  NAND2_X1 U544 ( .A1(n508), .A2(n483), .ZN(n484) );
  NAND2_X1 U545 ( .A1(n493), .A2(n509), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n488) );
  NAND2_X1 U548 ( .A1(n493), .A2(n512), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U550 ( .A(G36GAT), .B(n489), .ZN(G1329GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n491) );
  NAND2_X1 U552 ( .A1(n493), .A2(n524), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U554 ( .A(n492), .B(G43GAT), .Z(G1330GAT) );
  XOR2_X1 U555 ( .A(G50GAT), .B(KEYINPUT109), .Z(n495) );
  NAND2_X1 U556 ( .A1(n493), .A2(n516), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1331GAT) );
  XNOR2_X1 U558 ( .A(KEYINPUT110), .B(n543), .ZN(n557) );
  NOR2_X1 U559 ( .A1(n557), .A2(n527), .ZN(n496) );
  XOR2_X1 U560 ( .A(KEYINPUT111), .B(n496), .Z(n507) );
  AND2_X1 U561 ( .A1(n507), .A2(n497), .ZN(n502) );
  NAND2_X1 U562 ( .A1(n502), .A2(n509), .ZN(n498) );
  XNOR2_X1 U563 ( .A(KEYINPUT42), .B(n498), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NAND2_X1 U565 ( .A1(n512), .A2(n502), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n500), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U567 ( .A1(n524), .A2(n502), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n501), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n504) );
  NAND2_X1 U570 ( .A1(n502), .A2(n516), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(n506) );
  XOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT112), .Z(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(G1335GAT) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(KEYINPUT114), .ZN(n511) );
  AND2_X1 U575 ( .A1(n508), .A2(n507), .ZN(n517) );
  NAND2_X1 U576 ( .A1(n517), .A2(n509), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n517), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U580 ( .A(G99GAT), .B(KEYINPUT115), .Z(n515) );
  NAND2_X1 U581 ( .A1(n517), .A2(n524), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT116), .B(KEYINPUT44), .Z(n519) );
  NAND2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U586 ( .A(G106GAT), .B(n520), .Z(G1339GAT) );
  XOR2_X1 U587 ( .A(G113GAT), .B(KEYINPUT119), .Z(n529) );
  NOR2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U589 ( .A(KEYINPUT118), .B(n523), .Z(n539) );
  NAND2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U591 ( .A1(n539), .A2(n526), .ZN(n530) );
  NAND2_X1 U592 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  INV_X1 U594 ( .A(n530), .ZN(n535) );
  NOR2_X1 U595 ( .A1(n557), .A2(n535), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U598 ( .A1(n573), .A2(n535), .ZN(n533) );
  XOR2_X1 U599 ( .A(KEYINPUT50), .B(n533), .Z(n534) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  NOR2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n538) );
  XNOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U605 ( .A(KEYINPUT120), .B(n541), .Z(n551) );
  NOR2_X1 U606 ( .A1(n565), .A2(n551), .ZN(n542) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n542), .Z(G1344GAT) );
  NOR2_X1 U608 ( .A1(n551), .A2(n543), .ZN(n548) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(KEYINPUT121), .B(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n551), .A2(n573), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(KEYINPUT123), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n553), .Z(G1347GAT) );
  NOR2_X1 U619 ( .A1(n565), .A2(n561), .ZN(n556) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT125), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1348GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n561), .ZN(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(n560), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n573), .A2(n561), .ZN(n562) );
  XOR2_X1 U628 ( .A(G183GAT), .B(n562), .Z(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n577) );
  NOR2_X1 U630 ( .A1(n565), .A2(n577), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  INV_X1 U635 ( .A(n577), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n577), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

