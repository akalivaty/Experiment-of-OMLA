//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  INV_X1    g005(.A(G131), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G137), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n188), .A2(G137), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n190), .A2(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(G131), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT69), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n197), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n205), .B2(G146), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT65), .B1(new_n211), .B2(G143), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n205), .A3(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(KEYINPUT64), .A3(G143), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n210), .A2(new_n212), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n208), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n194), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n203), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n216), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(new_n224), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n202), .A2(new_n219), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT66), .A2(G116), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT66), .A2(G116), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(G119), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G119), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G113), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT2), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT2), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G113), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT66), .A2(G116), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT66), .A2(G116), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n234), .B1(new_n244), .B2(G119), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n240), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT67), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AND4_X1   g061(.A1(KEYINPUT67), .A2(new_n232), .A3(new_n235), .A4(new_n246), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n241), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n232), .A2(new_n235), .A3(new_n246), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT68), .A3(new_n241), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n229), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT73), .ZN(new_n260));
  OR2_X1    g074(.A1(KEYINPUT71), .A2(G237), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT71), .A2(G237), .ZN(new_n262));
  AOI21_X1  g076(.A(G953), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n260), .B(new_n264), .ZN(new_n265));
  XOR2_X1   g079(.A(KEYINPUT72), .B(KEYINPUT27), .Z(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n229), .A2(new_n251), .A3(new_n255), .A4(KEYINPUT70), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n258), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n269), .A2(KEYINPUT74), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n249), .A2(new_n250), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT68), .B1(new_n254), .B2(new_n241), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n229), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(KEYINPUT30), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n228), .A2(new_n222), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n219), .A2(new_n194), .A3(new_n197), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(KEYINPUT30), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n274), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n258), .A2(new_n267), .A3(new_n282), .A4(new_n268), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT31), .B1(new_n270), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n279), .B1(new_n271), .B2(new_n272), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n258), .A2(new_n268), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT28), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n256), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n267), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n269), .A2(KEYINPUT74), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT31), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n283), .A4(new_n281), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n285), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT75), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n297), .A2(new_n302), .A3(new_n298), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n299), .A2(new_n301), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n281), .A2(new_n258), .A3(new_n268), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n292), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n288), .A2(new_n267), .A3(new_n290), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT76), .B(G902), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n275), .B1(new_n271), .B2(new_n272), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n258), .A2(new_n313), .A3(new_n268), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT28), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n290), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n267), .A2(KEYINPUT29), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G472), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n304), .A2(new_n306), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n321));
  OAI22_X1  g135(.A1(new_n217), .A2(G119), .B1(KEYINPUT78), .B2(KEYINPUT23), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT79), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n326));
  INV_X1    g140(.A(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G128), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n326), .A2(new_n328), .A3(new_n329), .A4(new_n323), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n217), .A2(G119), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G110), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n328), .A2(new_n331), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT24), .B(G110), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n336), .B1(new_n335), .B2(new_n339), .ZN(new_n342));
  XNOR2_X1  g156(.A(G125), .B(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT16), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT16), .ZN(new_n345));
  INV_X1    g159(.A(G140), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(G125), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(G146), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n211), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n341), .A2(new_n342), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n332), .A2(new_n334), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G110), .ZN(new_n353));
  AOI21_X1  g167(.A(G146), .B1(new_n344), .B2(new_n347), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n348), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n337), .A2(new_n338), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT80), .A4(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n346), .A2(G125), .ZN(new_n360));
  INV_X1    g174(.A(G125), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G140), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n347), .B1(new_n363), .B2(new_n345), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(new_n211), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n357), .B1(new_n365), .B2(new_n354), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n333), .B1(new_n332), .B2(new_n334), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n359), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n358), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n321), .B1(new_n351), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n335), .A2(new_n339), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT81), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n372), .A2(new_n340), .A3(new_n349), .A4(new_n348), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(KEYINPUT82), .A3(new_n368), .A4(new_n358), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT22), .B(G137), .ZN(new_n375));
  INV_X1    g189(.A(G953), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n376), .A2(G221), .A3(G234), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n375), .B(new_n377), .Z(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n370), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n321), .B(new_n378), .C1(new_n351), .C2(new_n369), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G217), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n312), .B2(G234), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G902), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT25), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(new_n387), .A3(new_n312), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n384), .B(KEYINPUT77), .Z(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n312), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n380), .B2(new_n381), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(new_n387), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n386), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n263), .A2(G143), .A3(G214), .ZN(new_n399));
  AND2_X1   g213(.A1(KEYINPUT71), .A2(G237), .ZN(new_n400));
  NOR2_X1   g214(.A1(KEYINPUT71), .A2(G237), .ZN(new_n401));
  OAI211_X1 g215(.A(G214), .B(new_n376), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n205), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT18), .A2(G131), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT88), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT88), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n399), .A2(new_n403), .A3(new_n408), .A4(new_n405), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n399), .A2(new_n403), .A3(KEYINPUT87), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n406), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n363), .A2(G146), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n349), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n404), .A2(G131), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT17), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n399), .A2(new_n403), .A3(new_n192), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n356), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n404), .A2(KEYINPUT17), .A3(G131), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n398), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n417), .A2(new_n398), .A3(new_n424), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT89), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT89), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n417), .A2(new_n424), .A3(new_n428), .A4(new_n398), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n425), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G475), .B1(new_n430), .B2(G902), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n427), .A2(new_n429), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n418), .A2(new_n420), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n343), .B(KEYINPUT19), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n434), .B(new_n348), .C1(G146), .C2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n398), .B1(new_n417), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n432), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n438), .B1(new_n427), .B2(new_n429), .ZN(new_n443));
  INV_X1    g257(.A(new_n441), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n443), .A2(KEYINPUT20), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n431), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT90), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT91), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n233), .B2(G122), .ZN(new_n450));
  INV_X1    g264(.A(G122), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT91), .A3(G116), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n230), .A2(G122), .A3(new_n231), .ZN(new_n454));
  INV_X1    g268(.A(G107), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n205), .A2(G128), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n217), .A2(G143), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT93), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT93), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n188), .ZN(new_n464));
  OR3_X1    g278(.A1(new_n454), .A2(KEYINPUT95), .A3(KEYINPUT14), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT95), .B1(new_n454), .B2(KEYINPUT14), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n454), .A2(KEYINPUT14), .ZN(new_n467));
  AND4_X1   g281(.A1(new_n453), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n456), .B(new_n464), .C1(new_n468), .C2(new_n455), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT9), .B(G234), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n470), .A2(new_n383), .A3(G953), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n453), .A2(new_n454), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G107), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n473), .A2(new_n456), .B1(new_n463), .B2(new_n188), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n458), .A2(KEYINPUT13), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT92), .A3(new_n457), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT13), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n457), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT92), .B1(new_n475), .B2(new_n457), .ZN(new_n479));
  OAI21_X1  g293(.A(G134), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT94), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n474), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n474), .B2(new_n480), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n469), .B(new_n471), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT96), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n484), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n482), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n489), .A2(KEYINPUT96), .A3(new_n469), .A4(new_n471), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n469), .B1(new_n483), .B2(new_n484), .ZN(new_n491));
  INV_X1    g305(.A(new_n471), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n487), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n312), .ZN(new_n495));
  INV_X1    g309(.A(G478), .ZN(new_n496));
  NOR2_X1   g310(.A1(KEYINPUT97), .A2(KEYINPUT15), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(KEYINPUT97), .A2(KEYINPUT15), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n500), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n494), .A2(new_n312), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(G234), .A2(G237), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n505), .A2(G952), .A3(new_n376), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n391), .A2(G953), .A3(new_n505), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT21), .B(G898), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(KEYINPUT90), .B(new_n431), .C1(new_n442), .C2(new_n445), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n448), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G214), .B1(G237), .B2(G902), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n514), .B(G113), .C1(KEYINPUT5), .C2(new_n235), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n254), .ZN(new_n516));
  INV_X1    g330(.A(G101), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n397), .A2(G107), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n455), .A2(KEYINPUT3), .A3(G104), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT3), .B1(new_n455), .B2(G104), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n517), .B(new_n518), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n397), .A2(G107), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT83), .B1(new_n455), .B2(G104), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT83), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n397), .A3(G107), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n522), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n521), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n516), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G110), .B(G122), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G101), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT4), .A3(new_n521), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT4), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n533), .A3(G101), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n528), .B(new_n529), .C1(new_n273), .C2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n529), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n535), .B1(new_n251), .B2(new_n255), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n516), .A2(new_n527), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n536), .A2(KEYINPUT6), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT6), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n542), .B(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n216), .A2(new_n218), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n361), .A3(new_n208), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n361), .B2(new_n228), .ZN(new_n546));
  INV_X1    g360(.A(G224), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(G953), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n546), .B(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n541), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT7), .B1(new_n547), .B2(G953), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n546), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n516), .B(new_n527), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n529), .B(KEYINPUT8), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(G902), .B1(new_n555), .B2(new_n536), .ZN(new_n556));
  OAI21_X1  g370(.A(G210), .B1(G237), .B2(G902), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n550), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n557), .B1(new_n550), .B2(new_n556), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n513), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G221), .B1(new_n470), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G110), .B(G140), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n376), .A2(G227), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n526), .A2(new_n517), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n216), .A2(new_n207), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n216), .A2(new_n218), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n521), .B(new_n568), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n544), .A2(new_n527), .A3(new_n208), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n222), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT84), .B(new_n567), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT84), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n574), .B1(new_n571), .B2(new_n572), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(KEYINPUT12), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(KEYINPUT12), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n571), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n532), .A2(new_n228), .A3(new_n534), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n219), .A2(new_n568), .A3(KEYINPUT10), .A4(new_n521), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n582), .A2(new_n574), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n566), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n566), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n222), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT85), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(KEYINPUT85), .A3(new_n222), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G469), .B1(new_n594), .B2(G902), .ZN(new_n595));
  INV_X1    g409(.A(G469), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n592), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n566), .B1(new_n597), .B2(new_n585), .ZN(new_n598));
  INV_X1    g412(.A(new_n587), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n580), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n596), .B(new_n312), .C1(new_n598), .C2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n563), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n512), .A2(new_n561), .A3(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n320), .A2(new_n395), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(new_n517), .ZN(G3));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n485), .A2(KEYINPUT33), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n494), .A2(new_n607), .B1(new_n493), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(G478), .A3(new_n312), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n495), .A2(new_n496), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n511), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT20), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n440), .A2(new_n614), .A3(new_n441), .ZN(new_n615));
  INV_X1    g429(.A(new_n432), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n443), .B2(new_n444), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT90), .B1(new_n618), .B2(new_n431), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n612), .B1(new_n613), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n509), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n558), .B1(new_n560), .B2(new_n622), .ZN(new_n623));
  AOI211_X1 g437(.A(KEYINPUT98), .B(new_n557), .C1(new_n550), .C2(new_n556), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n621), .B(new_n513), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n297), .A2(new_n302), .A3(new_n298), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n302), .B1(new_n297), .B2(new_n298), .ZN(new_n628));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n297), .B2(new_n312), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n603), .A2(new_n394), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n626), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  NAND3_X1  g449(.A1(new_n440), .A2(new_n441), .A3(new_n432), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n617), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n504), .A2(new_n431), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n625), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n631), .A3(new_n632), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n351), .A2(new_n369), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n379), .A2(KEYINPUT36), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT99), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n646), .A2(new_n385), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n390), .B2(new_n393), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT100), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n652), .B(new_n649), .C1(new_n390), .C2(new_n393), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n604), .A2(new_n631), .A3(new_n651), .A4(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n506), .B1(new_n507), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n431), .A2(new_n504), .A3(new_n637), .A4(new_n659), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n602), .A2(new_n651), .A3(new_n660), .A4(new_n653), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n513), .B1(new_n623), .B2(new_n624), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n320), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  NOR2_X1   g479(.A1(new_n559), .A2(new_n560), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT38), .ZN(new_n667));
  INV_X1    g481(.A(new_n513), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n667), .A2(new_n668), .A3(new_n650), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n658), .B(KEYINPUT39), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n602), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT40), .Z(new_n672));
  INV_X1    g486(.A(new_n284), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n673), .A2(new_n294), .B1(new_n292), .B2(new_n314), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n674), .B2(G902), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n304), .A2(new_n306), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n504), .B1(new_n613), .B2(new_n619), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n669), .A2(new_n672), .A3(new_n676), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  NAND2_X1  g494(.A1(new_n651), .A2(new_n653), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n603), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n612), .B(new_n659), .C1(new_n613), .C2(new_n619), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n320), .A2(new_n682), .A3(new_n663), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  NOR2_X1   g500(.A1(new_n596), .A2(KEYINPUT101), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n588), .A2(KEYINPUT85), .A3(new_n222), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT85), .B1(new_n588), .B2(new_n222), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n585), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n566), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n690), .A2(new_n691), .B1(new_n599), .B2(new_n580), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n687), .B1(new_n692), .B2(new_n391), .ZN(new_n693));
  INV_X1    g507(.A(new_n687), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n312), .B(new_n694), .C1(new_n598), .C2(new_n600), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n693), .A2(new_n562), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n320), .A2(new_n395), .A3(new_n626), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NOR2_X1   g513(.A1(new_n627), .A2(new_n628), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n305), .B1(new_n700), .B2(new_n301), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n394), .B1(new_n701), .B2(new_n319), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n702), .A2(new_n703), .A3(new_n639), .A4(new_n696), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n320), .A2(new_n395), .A3(new_n639), .A4(new_n696), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT102), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NAND4_X1  g522(.A1(new_n696), .A2(new_n448), .A3(new_n511), .A4(new_n510), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n681), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n320), .A2(new_n710), .A3(new_n663), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NAND2_X1  g526(.A1(new_n696), .A2(new_n621), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n677), .A2(new_n713), .A3(new_n662), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n298), .B(KEYINPUT103), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n294), .A2(new_n283), .A3(new_n281), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n716), .A2(KEYINPUT31), .B1(new_n316), .B2(new_n292), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n715), .B1(new_n717), .B2(new_n296), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n630), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT104), .B1(new_n719), .B2(new_n395), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n630), .A2(new_n394), .A3(new_n718), .A4(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n714), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  NAND2_X1  g538(.A1(new_n717), .A2(new_n296), .ZN(new_n725));
  INV_X1    g539(.A(new_n715), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n297), .A2(new_n312), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n650), .B(new_n727), .C1(new_n728), .C2(new_n629), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n683), .ZN(new_n730));
  INV_X1    g544(.A(new_n696), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n662), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  NAND2_X1  g548(.A1(new_n299), .A2(new_n301), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n306), .A2(new_n319), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n736), .A2(new_n395), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n602), .A2(new_n666), .A3(new_n513), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(KEYINPUT42), .A3(new_n684), .A4(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n320), .A2(new_n395), .A3(new_n684), .A4(new_n739), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(KEYINPUT105), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n741), .B2(KEYINPUT105), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n740), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  NAND4_X1  g560(.A1(new_n320), .A2(new_n395), .A3(new_n660), .A4(new_n739), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT106), .B(G134), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G36));
  XOR2_X1   g563(.A(new_n594), .B(KEYINPUT45), .Z(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(G469), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(G469), .A2(G902), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n601), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT46), .B1(new_n753), .B2(new_n754), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n562), .B(new_n670), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n666), .A2(new_n513), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n448), .A2(new_n511), .A3(new_n612), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(KEYINPUT43), .Z(new_n762));
  INV_X1    g576(.A(new_n631), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n650), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n759), .B(new_n766), .C1(new_n765), .C2(new_n764), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  OAI21_X1  g582(.A(new_n562), .B1(new_n756), .B2(new_n757), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n320), .A2(new_n395), .A3(new_n683), .A4(new_n760), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT108), .B(G140), .Z(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G42));
  AND2_X1   g591(.A1(new_n762), .A2(new_n506), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n731), .A2(new_n760), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n729), .ZN(new_n781));
  INV_X1    g595(.A(new_n676), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n395), .A3(new_n506), .A4(new_n779), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n448), .A2(new_n511), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n783), .A2(new_n784), .A3(new_n612), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT51), .B1(new_n787), .B2(KEYINPUT114), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n788), .B1(KEYINPUT114), .B2(new_n787), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n720), .A2(new_n722), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n778), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n668), .A3(new_n667), .A4(new_n696), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT50), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n693), .A2(new_n695), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n563), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n771), .A2(new_n772), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n760), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n791), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n798), .B2(new_n799), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n789), .B(new_n795), .C1(new_n800), .C2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT48), .ZN(new_n805));
  INV_X1    g619(.A(new_n737), .ZN(new_n806));
  OAI211_X1 g620(.A(KEYINPUT117), .B(new_n805), .C1(new_n780), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n791), .A2(new_n732), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT116), .Z(new_n809));
  NOR2_X1   g623(.A1(new_n780), .A2(new_n806), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n805), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n376), .A2(G952), .ZN(new_n814));
  INV_X1    g628(.A(new_n783), .ZN(new_n815));
  INV_X1    g629(.A(new_n620), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n807), .A2(new_n809), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n786), .B1(new_n798), .B2(new_n802), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n795), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n804), .B(new_n818), .C1(new_n820), .C2(KEYINPUT51), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n697), .A2(new_n723), .A3(new_n711), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n704), .B2(new_n706), .ZN(new_n824));
  INV_X1    g638(.A(new_n561), .ZN(new_n825));
  INV_X1    g639(.A(new_n504), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n784), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n621), .B(new_n825), .C1(new_n816), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n631), .A2(new_n632), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n654), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n605), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n431), .A2(new_n826), .A3(new_n637), .A4(new_n659), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n320), .A2(new_n682), .A3(new_n801), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT110), .B1(new_n730), .B2(new_n739), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n729), .A2(new_n683), .A3(new_n738), .A4(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n747), .B(new_n833), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n745), .A2(new_n824), .A3(new_n831), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n677), .A2(new_n662), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n603), .A2(new_n650), .A3(new_n658), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n676), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n685), .A2(new_n664), .A3(new_n842), .A4(new_n733), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n822), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n664), .A2(new_n733), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(KEYINPUT52), .A3(new_n685), .A4(new_n842), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n843), .A2(new_n844), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(KEYINPUT111), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT111), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT105), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n702), .A2(new_n857), .A3(new_n684), .A4(new_n739), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n741), .A2(KEYINPUT105), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n743), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n837), .B1(new_n860), .B2(new_n740), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n705), .B(new_n703), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT112), .B1(new_n862), .B2(new_n823), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n824), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n831), .A2(KEYINPUT53), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n861), .A2(new_n863), .A3(new_n865), .A4(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n848), .B(new_n849), .C1(new_n856), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n823), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n707), .A2(new_n831), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n851), .A2(new_n852), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n861), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT53), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n861), .A3(new_n822), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n874), .B1(new_n875), .B2(new_n856), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n869), .B1(new_n876), .B2(new_n849), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n821), .A2(new_n877), .B1(G952), .B2(G953), .ZN(new_n878));
  INV_X1    g692(.A(new_n667), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n796), .B(KEYINPUT49), .Z(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n880), .A3(new_n761), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n395), .A2(new_n513), .A3(new_n562), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT109), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n782), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n376), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n861), .A2(new_n863), .A3(new_n865), .A4(new_n867), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT111), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n845), .B2(new_n846), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n853), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n888), .A2(new_n891), .B1(new_n822), .B2(new_n873), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n312), .ZN(new_n893));
  INV_X1    g707(.A(new_n557), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT56), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n541), .A2(new_n543), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n549), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT55), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n887), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n895), .B2(new_n898), .ZN(G51));
  OAI21_X1  g714(.A(KEYINPUT119), .B1(new_n892), .B2(new_n849), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n848), .B1(new_n856), .B2(new_n868), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT54), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n869), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n824), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n866), .B1(new_n907), .B2(KEYINPUT112), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n891), .A2(new_n861), .A3(new_n908), .A4(new_n865), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(KEYINPUT118), .A3(new_n849), .A4(new_n848), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n901), .A2(new_n904), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n754), .B(KEYINPUT57), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT120), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n914));
  INV_X1    g728(.A(new_n912), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT54), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n903), .B1(new_n902), .B2(KEYINPUT54), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n906), .A2(new_n910), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n914), .B(new_n915), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n692), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n913), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n753), .B(KEYINPUT121), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n893), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n886), .B1(new_n922), .B2(new_n924), .ZN(G54));
  AND3_X1   g739(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n887), .B1(new_n926), .B2(new_n440), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n440), .B2(new_n926), .ZN(G60));
  XNOR2_X1  g742(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n609), .B1(new_n877), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n911), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n609), .A2(new_n931), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n886), .B(new_n932), .C1(new_n933), .C2(new_n934), .ZN(G63));
  INV_X1    g749(.A(G902), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT60), .B1(new_n383), .B2(new_n936), .ZN(new_n937));
  OR3_X1    g751(.A1(new_n383), .A2(new_n936), .A3(KEYINPUT60), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n902), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n887), .B1(new_n939), .B2(new_n382), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n646), .A2(new_n647), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n939), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT61), .ZN(G66));
  NOR3_X1   g757(.A1(new_n508), .A2(new_n547), .A3(new_n376), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n871), .B2(new_n376), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n896), .B1(G898), .B2(new_n376), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  NOR2_X1   g761(.A1(new_n276), .A2(new_n280), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n436), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(G227), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n950), .A2(new_n657), .A3(new_n376), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n850), .A2(new_n685), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n767), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n737), .A2(new_n840), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n747), .B1(new_n758), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n773), .B2(new_n774), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n745), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n949), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n961), .A2(KEYINPUT123), .ZN(new_n962));
  XNOR2_X1  g776(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n952), .A2(new_n679), .ZN(new_n964));
  MUX2_X1   g778(.A(new_n962), .B(new_n963), .S(new_n964), .Z(new_n965));
  NOR2_X1   g779(.A1(new_n816), .A2(new_n827), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n966), .A2(new_n671), .A3(new_n760), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n967), .A2(new_n702), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT124), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n965), .A2(new_n767), .A3(new_n775), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n960), .B1(new_n949), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n951), .B1(new_n971), .B2(new_n376), .ZN(G72));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT63), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT126), .ZN(new_n975));
  INV_X1    g789(.A(new_n871), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n970), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n267), .A3(new_n307), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n308), .A2(new_n716), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n979), .A2(new_n974), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n876), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n955), .A2(new_n745), .A3(new_n871), .A4(new_n958), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n983), .A2(new_n975), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n307), .A2(new_n267), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n982), .B(new_n887), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n983), .B2(new_n975), .ZN(new_n988));
  OAI21_X1  g802(.A(KEYINPUT127), .B1(new_n988), .B2(new_n886), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n981), .B1(new_n987), .B2(new_n989), .ZN(G57));
endmodule


