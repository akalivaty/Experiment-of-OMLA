//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n637,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1219, new_n1220, new_n1221;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G137), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n466), .B(new_n470), .C1(new_n472), .C2(new_n467), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n465), .A2(new_n475), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n483), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n467), .B1(new_n462), .B2(new_n464), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n484), .A2(new_n485), .B1(G124), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n479), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT72), .Z(G162));
  NAND2_X1  g064(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n460), .A2(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(new_n467), .A3(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT76), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n493), .A2(new_n467), .A3(G138), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n471), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n462), .A2(new_n464), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n467), .A2(G138), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n495), .A2(new_n498), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n486), .A2(G126), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n467), .B1(KEYINPUT73), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G114), .ZN(new_n509));
  AOI211_X1 g084(.A(KEYINPUT74), .B(new_n505), .C1(new_n507), .C2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(KEYINPUT73), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n509), .A2(new_n512), .A3(G2105), .ZN(new_n513));
  INV_X1    g088(.A(new_n505), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n504), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT75), .ZN(new_n517));
  OAI21_X1  g092(.A(G2105), .B1(new_n508), .B2(G114), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n506), .A2(KEYINPUT73), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n513), .A2(new_n511), .A3(new_n514), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(new_n504), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n503), .B1(new_n517), .B2(new_n525), .ZN(G164));
  AND2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G50), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n537), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G651), .ZN(new_n539));
  INV_X1    g114(.A(G88), .ZN(new_n540));
  AND2_X1   g115(.A1(KEYINPUT5), .A2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(KEYINPUT5), .A2(G543), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n528), .A2(new_n527), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n534), .A2(new_n544), .ZN(G166));
  NOR2_X1   g120(.A1(new_n541), .A2(new_n542), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n539), .ZN(new_n547));
  AOI22_X1  g122(.A1(G51), .A2(new_n531), .B1(new_n547), .B2(G63), .ZN(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT7), .ZN(new_n550));
  INV_X1    g125(.A(G89), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n551), .B2(new_n543), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n548), .B1(KEYINPUT78), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n552), .A2(KEYINPUT78), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(G168));
  OR2_X1    g130(.A1(new_n527), .A2(new_n528), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G52), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT79), .B(G90), .Z(new_n559));
  OAI22_X1  g134(.A1(new_n557), .A2(new_n558), .B1(new_n543), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n537), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(new_n539), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n560), .A2(new_n562), .ZN(G171));
  AOI22_X1  g138(.A1(new_n537), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n539), .ZN(new_n565));
  INV_X1    g140(.A(G43), .ZN(new_n566));
  INV_X1    g141(.A(G81), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n557), .A2(new_n566), .B1(new_n567), .B2(new_n543), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT80), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n565), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  NAND4_X1  g149(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND4_X1  g152(.A1(G319), .A2(G483), .A3(G661), .A4(new_n577), .ZN(G188));
  NAND2_X1  g153(.A1(new_n531), .A2(G53), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g155(.A1(G78), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G65), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n546), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n543), .ZN(new_n584));
  AOI22_X1  g159(.A1(G651), .A2(new_n583), .B1(new_n584), .B2(G91), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n580), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  INV_X1    g162(.A(G168), .ZN(G286));
  OR2_X1    g163(.A1(new_n534), .A2(new_n544), .ZN(G303));
  AOI22_X1  g164(.A1(G87), .A2(new_n584), .B1(new_n531), .B2(G49), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n591));
  NAND2_X1  g166(.A1(G74), .A2(G651), .ZN(new_n592));
  OAI211_X1 g167(.A(KEYINPUT81), .B(new_n592), .C1(new_n546), .C2(new_n539), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n594), .B(G651), .C1(new_n537), .C2(G74), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n590), .A2(new_n591), .A3(new_n593), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n531), .A2(G49), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n556), .A2(G87), .A3(new_n537), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n597), .A2(new_n593), .A3(new_n595), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT82), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G288));
  OAI21_X1  g177(.A(G61), .B1(new_n541), .B2(new_n542), .ZN(new_n603));
  NAND2_X1  g178(.A1(G73), .A2(G543), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n539), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n605), .A2(new_n606), .B1(new_n531), .B2(G48), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n608));
  INV_X1    g183(.A(G86), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n543), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n556), .A2(KEYINPUT84), .A3(G86), .A4(new_n537), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G61), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n535), .B2(new_n536), .ZN(new_n614));
  INV_X1    g189(.A(new_n604), .ZN(new_n615));
  OAI21_X1  g190(.A(G651), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT83), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n607), .A2(new_n612), .A3(new_n617), .ZN(G305));
  AOI22_X1  g193(.A1(G85), .A2(new_n584), .B1(new_n531), .B2(G47), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n537), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n539), .B2(new_n620), .ZN(G290));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NOR2_X1   g197(.A1(G301), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n584), .A2(G92), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(G79), .A2(G543), .ZN(new_n627));
  INV_X1    g202(.A(G66), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n546), .B2(new_n628), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n629), .A2(G651), .B1(new_n531), .B2(G54), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT85), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n623), .B1(new_n632), .B2(new_n622), .ZN(G284));
  AOI21_X1  g208(.A(new_n623), .B1(new_n632), .B2(new_n622), .ZN(G321));
  AND2_X1   g209(.A1(new_n580), .A2(new_n585), .ZN(new_n635));
  OAI21_X1  g210(.A(KEYINPUT86), .B1(new_n635), .B2(G868), .ZN(new_n636));
  NOR2_X1   g211(.A1(G168), .A2(new_n622), .ZN(new_n637));
  MUX2_X1   g212(.A(new_n636), .B(KEYINPUT86), .S(new_n637), .Z(G297));
  MUX2_X1   g213(.A(new_n636), .B(KEYINPUT86), .S(new_n637), .Z(G280));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n632), .B1(new_n640), .B2(G860), .ZN(G148));
  NAND2_X1  g216(.A1(new_n572), .A2(new_n622), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT85), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n631), .B(new_n643), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n644), .A2(G559), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n642), .B1(new_n645), .B2(new_n622), .ZN(G323));
  XNOR2_X1  g221(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g222(.A1(new_n486), .A2(G123), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n467), .A2(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n478), .B2(G135), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT87), .B(G2096), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT12), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT13), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n658), .ZN(G156));
  XOR2_X1   g234(.A(KEYINPUT15), .B(G2435), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2438), .ZN(new_n661));
  XOR2_X1   g236(.A(G2427), .B(G2430), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT88), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(KEYINPUT14), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2451), .B(G2454), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n666), .B(new_n670), .Z(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(new_n674), .A3(G14), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G401));
  XNOR2_X1  g251(.A(G2084), .B(G2090), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT89), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2072), .B(G2078), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT18), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT90), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n680), .B1(new_n683), .B2(new_n679), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n683), .B2(new_n679), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n685), .A2(new_n678), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n679), .B(KEYINPUT17), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n678), .B2(new_n680), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n678), .A2(new_n680), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n682), .B1(new_n686), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2096), .B(G2100), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(G227));
  XNOR2_X1  g270(.A(G1956), .B(G2474), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT91), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1961), .B(G1966), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1971), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT19), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT20), .Z(new_n704));
  OR2_X1    g279(.A1(new_n697), .A2(new_n699), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(new_n702), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n702), .A3(new_n700), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n714), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(G229));
  NAND2_X1  g292(.A1(new_n478), .A2(G131), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  INV_X1    g294(.A(G107), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G2105), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n486), .B2(G119), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G29), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G25), .B2(G29), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G24), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT92), .Z(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G290), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1986), .ZN(new_n733));
  AOI21_X1  g308(.A(KEYINPUT93), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n728), .B(new_n734), .C1(new_n733), .C2(new_n732), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n729), .A2(G22), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G166), .B2(new_n729), .ZN(new_n737));
  INV_X1    g312(.A(G1971), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(G6), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G305), .B2(new_n729), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT32), .B(G1981), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  MUX2_X1   g319(.A(G23), .B(new_n599), .S(G16), .Z(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT33), .B(G1976), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n739), .A2(new_n743), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n727), .B(new_n735), .C1(new_n748), .C2(KEYINPUT34), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(KEYINPUT34), .B2(new_n748), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT36), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G35), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G162), .B2(new_n752), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT29), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G2090), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT102), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n752), .A2(G27), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G164), .B2(new_n752), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT101), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n478), .A2(G139), .ZN(new_n763));
  NAND2_X1  g338(.A1(G115), .A2(G2104), .ZN(new_n764));
  INV_X1    g339(.A(G127), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n492), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n766), .A2(KEYINPUT96), .A3(G2105), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT25), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT96), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n763), .A2(new_n767), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  MUX2_X1   g348(.A(G33), .B(new_n773), .S(G29), .Z(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G2072), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n478), .A2(G141), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT26), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT98), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n778), .B(new_n780), .C1(G129), .C2(new_n486), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(new_n752), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n752), .B2(G32), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G2084), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT24), .B(G34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(new_n752), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT97), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n473), .B2(new_n752), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n775), .B(new_n787), .C1(new_n788), .C2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n761), .A2(KEYINPUT101), .ZN(new_n797));
  AND4_X1   g372(.A1(new_n762), .A2(new_n795), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT100), .B1(G16), .B2(G21), .ZN(new_n799));
  NAND2_X1  g374(.A1(G168), .A2(G16), .ZN(new_n800));
  MUX2_X1   g375(.A(KEYINPUT100), .B(new_n799), .S(new_n800), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1966), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n785), .A2(new_n786), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n729), .A2(G20), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT23), .Z(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G299), .B2(G16), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G1956), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n729), .A2(G5), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G171), .B2(new_n729), .ZN(new_n809));
  INV_X1    g384(.A(G1961), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n792), .A2(new_n788), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT31), .B(G11), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT30), .B(G28), .Z(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G29), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n652), .B2(G29), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n811), .A2(new_n812), .A3(new_n816), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n803), .A2(new_n807), .A3(new_n817), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n802), .B(new_n818), .C1(new_n755), .C2(G2090), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n752), .A2(G26), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT28), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n478), .A2(G140), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n823));
  INV_X1    g398(.A(G116), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(G2105), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n486), .B2(G128), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n821), .B1(new_n827), .B2(G29), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G2067), .ZN(new_n829));
  NOR2_X1   g404(.A1(G16), .A2(G19), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n573), .B2(G16), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT94), .B(G1341), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n632), .A2(G16), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G4), .B2(G16), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(G1348), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(G1348), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n829), .B(new_n833), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT95), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(KEYINPUT95), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n819), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND4_X1   g416(.A1(new_n751), .A2(new_n757), .A3(new_n798), .A4(new_n841), .ZN(G311));
  NAND4_X1  g417(.A1(new_n751), .A2(new_n757), .A3(new_n798), .A4(new_n841), .ZN(G150));
  INV_X1    g418(.A(G55), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n557), .A2(new_n844), .B1(new_n845), .B2(new_n543), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n537), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n539), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  OAI21_X1  g427(.A(KEYINPUT103), .B1(new_n644), .B2(new_n640), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n632), .A2(new_n854), .A3(G559), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT38), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n572), .A2(new_n850), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n565), .B(new_n849), .C1(new_n570), .C2(new_n571), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n863), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n857), .A2(new_n859), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(KEYINPUT39), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT104), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT39), .B1(new_n864), .B2(new_n866), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n852), .B1(new_n868), .B2(new_n870), .ZN(G145));
  NAND2_X1  g446(.A1(new_n773), .A2(KEYINPUT105), .ZN(new_n872));
  INV_X1    g447(.A(G126), .ZN(new_n873));
  AOI211_X1 g448(.A(new_n873), .B(new_n467), .C1(new_n462), .C2(new_n464), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n521), .B2(new_n522), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n492), .A2(KEYINPUT76), .A3(new_n494), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n497), .B1(new_n471), .B2(new_n496), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n500), .B1(new_n462), .B2(new_n464), .ZN(new_n878));
  OAI22_X1  g453(.A1(new_n876), .A2(new_n877), .B1(new_n493), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n872), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n486), .A2(G130), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n467), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n478), .B2(G142), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n656), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n881), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n782), .B(new_n827), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n723), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n890), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G162), .B(new_n652), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n473), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n891), .A2(new_n895), .A3(new_n892), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g476(.A(G303), .B(G305), .ZN(new_n902));
  XNOR2_X1  g477(.A(G290), .B(new_n599), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n903), .A2(new_n904), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n907), .A3(new_n905), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT42), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT109), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n645), .A2(new_n863), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n635), .A2(new_n626), .A3(new_n630), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n631), .A2(G299), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n865), .B1(new_n644), .B2(G559), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n912), .A2(new_n917), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n913), .A2(KEYINPUT41), .A3(new_n914), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT107), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n922), .A2(new_n930), .A3(new_n927), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n920), .A2(new_n921), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n910), .A2(KEYINPUT109), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n911), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n935));
  INV_X1    g510(.A(new_n910), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n921), .A2(new_n920), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n929), .A2(new_n931), .ZN(new_n938));
  AND4_X1   g513(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n850), .A2(new_n622), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(G295));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n941), .ZN(G331));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n906), .A2(new_n908), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n946));
  NAND2_X1  g521(.A1(G301), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n861), .B2(new_n862), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(G286), .B1(KEYINPUT110), .B2(G171), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n861), .A2(new_n862), .A3(new_n947), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n950), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n861), .A2(new_n862), .A3(new_n947), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(new_n948), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n927), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(new_n955), .A3(new_n916), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n945), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT111), .B1(new_n959), .B2(G37), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(new_n945), .A3(new_n958), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n958), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n926), .B1(new_n952), .B2(new_n955), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n909), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n967), .A3(new_n898), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n960), .A2(new_n963), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n961), .A3(new_n898), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n944), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n960), .A2(new_n968), .A3(new_n961), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n959), .A2(G37), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n973), .A2(KEYINPUT43), .B1(new_n974), .B2(new_n963), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n972), .B1(new_n975), .B2(new_n944), .ZN(G397));
  AOI21_X1  g551(.A(G1384), .B1(new_n875), .B2(new_n879), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n472), .A2(new_n467), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n978), .A2(G40), .A3(new_n466), .A4(new_n470), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n977), .A2(new_n979), .A3(KEYINPUT45), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n723), .A2(new_n726), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n723), .A2(new_n726), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G2067), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n827), .B(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n980), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n987), .B(KEYINPUT113), .Z(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n986), .A2(new_n989), .A3(new_n783), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n980), .A2(new_n989), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(new_n782), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT112), .ZN(new_n994));
  NOR2_X1   g569(.A1(G290), .A2(G1986), .ZN(new_n995));
  AND2_X1   g570(.A1(G290), .A2(G1986), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n980), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND4_X1   g572(.A1(new_n983), .A2(new_n991), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1000), .B(new_n1001), .C1(new_n516), .C2(new_n503), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n977), .A2(KEYINPUT114), .A3(new_n1000), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G40), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n473), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n999), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n810), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(G164), .B2(G1384), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n979), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n760), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1008), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G164), .A2(G1384), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1018), .B2(KEYINPUT45), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1015), .A2(G2078), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1010), .A2(new_n1016), .A3(new_n1021), .A4(G301), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1022), .A2(KEYINPUT54), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1001), .B1(new_n516), .B2(new_n503), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n979), .B1(new_n1024), .B2(new_n1011), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1020), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1025), .A2(new_n1027), .A3(KEYINPUT124), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT124), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1010), .A2(new_n1016), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT125), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1031), .A2(new_n1032), .A3(G171), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1031), .B2(G171), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1023), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI211_X1 g610(.A(KEYINPUT75), .B(new_n874), .C1(new_n521), .C2(new_n522), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n524), .B1(new_n523), .B2(new_n504), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n879), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT45), .B1(new_n1038), .B2(new_n1001), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1008), .B1(new_n1024), .B2(new_n1011), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n738), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G2090), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n999), .A2(new_n1006), .A3(new_n1042), .A4(new_n1008), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G8), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G166), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(G8), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n977), .A2(new_n1008), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n599), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(G8), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT52), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1045), .B1(new_n977), .B2(new_n1008), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n596), .A2(new_n600), .A3(new_n1051), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1052), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n584), .A2(G86), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n606), .B(G651), .C1(new_n614), .C2(new_n615), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n531), .A2(G48), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n617), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G1981), .ZN(new_n1064));
  INV_X1    g639(.A(G1981), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n607), .A2(new_n612), .A3(new_n1065), .A4(new_n617), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(KEYINPUT49), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT116), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1064), .A2(new_n1069), .A3(KEYINPUT49), .A4(new_n1066), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT49), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1068), .A2(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1059), .B1(new_n1073), .B2(new_n1055), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1049), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1048), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1038), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n979), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1077), .A2(new_n1042), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1971), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT119), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1077), .A2(new_n1042), .A3(new_n1078), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1041), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(G8), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1075), .B1(new_n1076), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n979), .A2(G2084), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n999), .A2(new_n1006), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1038), .A2(KEYINPUT45), .A3(new_n1001), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1966), .B1(new_n1089), .B2(new_n1025), .ZN(new_n1090));
  OAI211_X1 g665(.A(G8), .B(G168), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1966), .ZN(new_n1092));
  NOR3_X1   g667(.A1(G164), .A2(new_n1011), .A3(G1384), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1092), .B1(new_n1093), .B2(new_n1017), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n999), .A2(new_n1006), .A3(new_n1087), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1045), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G168), .A2(new_n1045), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1091), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(KEYINPUT51), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1031), .A2(G171), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1014), .A2(new_n1015), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1106));
  AOI21_X1  g681(.A(G301), .B1(new_n1106), .B2(new_n1010), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1104), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1035), .A2(new_n1086), .A3(new_n1103), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1038), .A2(new_n1001), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1040), .B1(new_n1110), .B2(new_n1011), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(G1956), .ZN(new_n1115));
  NAND2_X1  g690(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n635), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(G299), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1115), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1122), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1113), .B(new_n1124), .C1(G1956), .C2(new_n1114), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT61), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT58), .B(G1341), .Z(new_n1127));
  AOI22_X1  g702(.A1(new_n1111), .A2(new_n989), .B1(new_n1050), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(KEYINPUT59), .A3(new_n573), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1128), .B2(new_n572), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1126), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1050), .A2(G2067), .ZN(new_n1135));
  INV_X1    g710(.A(G1348), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n1009), .B2(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1137), .A2(new_n644), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n644), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1138), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1123), .A2(KEYINPUT61), .A3(new_n1125), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1134), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1138), .A2(new_n1123), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1125), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1109), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1085), .A2(new_n1076), .ZN(new_n1151));
  AOI211_X1 g726(.A(new_n1045), .B(G286), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(new_n1055), .A3(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1045), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1048), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1151), .A2(new_n1152), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1157), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1155), .A2(KEYINPUT117), .A3(new_n1156), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1158), .A2(new_n1048), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1091), .A2(new_n1161), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1166), .A2(new_n1049), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1100), .B1(new_n1171), .B2(G8), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(new_n1152), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1098), .B(G8), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1097), .ZN(new_n1175));
  AOI21_X1  g750(.A(KEYINPUT51), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT62), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1101), .B(new_n1178), .C1(new_n1102), .C2(KEYINPUT51), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1177), .A2(new_n1086), .A3(new_n1107), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT118), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1049), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1055), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1184), .A2(new_n1051), .A3(new_n601), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1183), .B1(new_n1185), .B2(new_n1066), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1181), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1066), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1055), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1155), .A2(new_n1156), .A3(KEYINPUT117), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT117), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g767(.A(KEYINPUT118), .B(new_n1189), .C1(new_n1192), .C2(new_n1049), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1187), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1170), .A2(new_n1180), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n998), .B1(new_n1150), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n991), .A2(new_n981), .A3(new_n994), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n822), .A2(new_n984), .A3(new_n826), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n986), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT46), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n992), .A2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT126), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n985), .B(new_n783), .C1(new_n1200), .C2(G1996), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n980), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  XOR2_X1   g780(.A(new_n1205), .B(KEYINPUT47), .Z(new_n1206));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n995), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT48), .ZN(new_n1208));
  AND4_X1   g783(.A1(new_n983), .A2(new_n991), .A3(new_n994), .A4(new_n1208), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1199), .A2(new_n1206), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1196), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g786(.A1(new_n693), .A2(G319), .A3(new_n694), .ZN(new_n1213));
  XOR2_X1   g787(.A(new_n1213), .B(KEYINPUT127), .Z(new_n1214));
  NAND2_X1  g788(.A1(new_n1214), .A2(new_n675), .ZN(new_n1215));
  AOI21_X1  g789(.A(new_n1215), .B1(new_n715), .B2(new_n716), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1216), .A2(new_n900), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n975), .A2(new_n1217), .ZN(G308));
  NAND2_X1  g792(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n963), .A2(new_n974), .ZN(new_n1220));
  NAND2_X1  g794(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g795(.A1(new_n1221), .A2(new_n900), .A3(new_n1216), .ZN(G225));
endmodule


