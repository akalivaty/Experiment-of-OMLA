//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(G234), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT25), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT73), .A2(G125), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(KEYINPUT73), .A2(G125), .A3(G140), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(KEYINPUT16), .A3(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT16), .B1(new_n195), .B2(G125), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n193), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n193), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n204), .A2(G128), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n205), .B(new_n207), .C1(new_n208), .C2(KEYINPUT23), .ZN(new_n209));
  OR2_X1    g023(.A1(new_n209), .A2(G110), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT71), .B1(new_n204), .B2(G128), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT71), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n206), .A3(G119), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n213), .A3(new_n205), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT74), .ZN(new_n215));
  INV_X1    g029(.A(G110), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT24), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G110), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT72), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n217), .B2(new_n219), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n214), .B(new_n215), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n210), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n217), .A2(new_n219), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT72), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n215), .B1(new_n228), .B2(new_n214), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n203), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n209), .A2(G110), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n198), .A2(new_n193), .A3(new_n200), .ZN(new_n232));
  OAI221_X1 g046(.A(new_n231), .B1(new_n228), .B2(new_n214), .C1(new_n232), .C2(new_n201), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT22), .B(G137), .ZN(new_n235));
  INV_X1    g049(.A(G953), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(G221), .A3(G234), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n235), .B(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n230), .A2(new_n233), .A3(new_n238), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n192), .B1(new_n242), .B2(G902), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n230), .A2(new_n233), .A3(new_n238), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n238), .B1(new_n230), .B2(new_n233), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT25), .A3(new_n189), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n191), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n190), .A2(G902), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n187), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT25), .B1(new_n246), .B2(new_n189), .ZN(new_n253));
  NOR4_X1   g067(.A1(new_n244), .A2(new_n245), .A3(new_n192), .A4(G902), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n190), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n250), .A3(KEYINPUT75), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G116), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(G119), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(KEYINPUT67), .A3(G119), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT67), .B1(new_n258), .B2(G119), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT2), .B(G113), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n266), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n204), .B2(G116), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n259), .B1(new_n270), .B2(new_n261), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n268), .B1(new_n271), .B2(KEYINPUT66), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  OR2_X1    g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  INV_X1    g089(.A(G143), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G146), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n193), .A2(G143), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n274), .B(new_n275), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n193), .A2(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(G146), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT0), .A4(G128), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G137), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT65), .B1(new_n284), .B2(G134), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n286));
  INV_X1    g100(.A(G134), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(G137), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT64), .B1(new_n287), .B2(G137), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT11), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT11), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT64), .B(new_n292), .C1(new_n287), .C2(G137), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G131), .ZN(new_n295));
  INV_X1    g109(.A(G131), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n289), .A2(new_n291), .A3(new_n296), .A4(new_n293), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n283), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n297), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT1), .B1(new_n276), .B2(G146), .ZN(new_n300));
  OAI211_X1 g114(.A(G128), .B(new_n300), .C1(new_n277), .C2(new_n278), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n280), .B(new_n281), .C1(KEYINPUT1), .C2(new_n206), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n284), .A2(G134), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n287), .A2(G137), .ZN(new_n304));
  OAI21_X1  g118(.A(G131), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n273), .B1(new_n298), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n295), .A2(new_n297), .ZN(new_n309));
  INV_X1    g123(.A(new_n283), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n301), .A2(new_n302), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n297), .A3(new_n305), .ZN(new_n314));
  INV_X1    g128(.A(new_n273), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n308), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n298), .A2(new_n307), .A3(new_n273), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT28), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(G237), .A2(G953), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G210), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT27), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G101), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT30), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n311), .A2(new_n329), .A3(new_n314), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT30), .B1(new_n298), .B2(new_n307), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n319), .B1(new_n332), .B2(new_n273), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n328), .B1(new_n333), .B2(new_n326), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n315), .B1(new_n330), .B2(new_n331), .ZN(new_n335));
  INV_X1    g149(.A(new_n326), .ZN(new_n336));
  NOR4_X1   g150(.A1(new_n335), .A2(KEYINPUT68), .A3(new_n336), .A4(new_n319), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT31), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n329), .B1(new_n311), .B2(new_n314), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n298), .A2(new_n307), .A3(KEYINPUT30), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n273), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n326), .A3(new_n316), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT31), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n327), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(G472), .A2(G902), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT32), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n327), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n342), .A2(KEYINPUT68), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n333), .A2(new_n328), .A3(new_n326), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n343), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n344), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n349), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT32), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(new_n346), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n348), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n321), .A2(new_n326), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n333), .A2(new_n326), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n189), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT69), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n298), .A2(new_n307), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(new_n315), .ZN(new_n365));
  NOR4_X1   g179(.A1(new_n298), .A2(new_n307), .A3(new_n273), .A4(KEYINPUT69), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT70), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n308), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(KEYINPUT70), .B(new_n273), .C1(new_n298), .C2(new_n307), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n317), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NOR4_X1   g186(.A1(new_n372), .A2(new_n359), .A3(new_n336), .A4(new_n320), .ZN(new_n373));
  OAI21_X1  g187(.A(G472), .B1(new_n362), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n257), .B1(new_n357), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n236), .A2(G227), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT76), .ZN(new_n377));
  XOR2_X1   g191(.A(G110), .B(G140), .Z(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G107), .ZN(new_n383));
  OR2_X1    g197(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n383), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n382), .A2(G107), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n384), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G101), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(new_n388), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n383), .A4(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n392), .A2(KEYINPUT4), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n399), .B(G101), .C1(new_n387), .C2(new_n391), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n310), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n381), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n385), .A2(G104), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n388), .B2(new_n389), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n395), .B1(new_n404), .B2(new_n394), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n283), .B1(new_n405), .B2(new_n399), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n392), .A2(KEYINPUT4), .A3(new_n397), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(KEYINPUT79), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G101), .B1(new_n389), .B2(new_n403), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n397), .A2(new_n302), .A3(new_n301), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT10), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT10), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n313), .A2(new_n412), .A3(new_n397), .A4(new_n409), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n402), .A2(new_n408), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n309), .A2(KEYINPUT80), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n295), .A2(new_n416), .A3(new_n297), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n380), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT81), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n309), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n411), .A2(new_n413), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n406), .A2(KEYINPUT79), .A3(new_n407), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT79), .B1(new_n406), .B2(new_n407), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n420), .B(new_n422), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n419), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n397), .A2(new_n409), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n312), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n410), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n309), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT12), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(KEYINPUT12), .A3(new_n309), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n418), .B(new_n422), .C1(new_n423), .C2(new_n424), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n379), .B(KEYINPUT77), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(G902), .B1(new_n427), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G469), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT82), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT81), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n309), .A3(new_n425), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n379), .B1(new_n445), .B2(new_n436), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n435), .A2(new_n379), .A3(new_n436), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n441), .B(new_n189), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n445), .A2(new_n419), .B1(new_n437), .B2(new_n438), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n449), .B(G469), .C1(new_n450), .C2(G902), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n442), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G214), .B1(G237), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n236), .A2(G952), .ZN(new_n455));
  NAND2_X1  g269(.A1(G234), .A2(G237), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT92), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(G898), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(G902), .A3(G953), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G210), .B1(G237), .B2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n273), .A2(new_n407), .A3(new_n400), .ZN(new_n466));
  OAI211_X1 g280(.A(KEYINPUT5), .B(new_n260), .C1(new_n262), .C2(new_n263), .ZN(new_n467));
  INV_X1    g281(.A(G113), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT5), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n259), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n271), .A2(new_n268), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n471), .A2(new_n397), .A3(new_n409), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G122), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n466), .A2(new_n473), .A3(new_n475), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n283), .A2(G125), .ZN(new_n480));
  INV_X1    g294(.A(G125), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n312), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G224), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(G953), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n480), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n481), .B1(new_n279), .B2(new_n282), .ZN(new_n487));
  AOI21_X1  g301(.A(G125), .B1(new_n301), .B2(new_n302), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n474), .A2(new_n491), .A3(new_n476), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n479), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n189), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n485), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n475), .B(KEYINPUT8), .ZN(new_n498));
  INV_X1    g312(.A(new_n473), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n471), .A2(new_n472), .B1(new_n397), .B2(new_n409), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT83), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n496), .B1(new_n482), .B2(new_n480), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n497), .A2(new_n501), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n478), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n503), .B1(new_n490), .B2(new_n496), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n502), .B1(new_n507), .B2(new_n501), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n465), .B1(new_n494), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n501), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT83), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n478), .A3(new_n505), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n513), .A2(new_n189), .A3(new_n464), .A4(new_n493), .ZN(new_n514));
  AOI211_X1 g328(.A(new_n454), .B(new_n463), .C1(new_n510), .C2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n232), .B2(new_n201), .ZN(new_n517));
  AND3_X1   g331(.A1(KEYINPUT73), .A2(G125), .A3(G140), .ZN(new_n518));
  AOI21_X1  g332(.A(G140), .B1(KEYINPUT73), .B2(G125), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT16), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(G146), .B1(new_n521), .B2(new_n199), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n198), .A2(new_n193), .A3(new_n200), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(KEYINPUT88), .A3(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(KEYINPUT84), .A2(G143), .ZN(new_n525));
  NAND2_X1  g339(.A1(KEYINPUT84), .A2(G143), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n525), .A2(new_n526), .B1(new_n322), .B2(G214), .ZN(new_n527));
  INV_X1    g341(.A(G237), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n236), .A3(G214), .ZN(new_n529));
  NOR2_X1   g343(.A1(KEYINPUT84), .A2(G143), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(G131), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n533));
  INV_X1    g347(.A(new_n526), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n529), .B1(new_n534), .B2(new_n530), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n525), .A2(G214), .A3(new_n322), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n296), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n296), .B1(new_n535), .B2(new_n536), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT17), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n517), .A2(new_n524), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(G113), .B(G122), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n382), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT18), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT85), .ZN(new_n545));
  OAI211_X1 g359(.A(G131), .B(new_n545), .C1(new_n527), .C2(new_n531), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n535), .B(new_n536), .C1(KEYINPUT85), .C2(new_n544), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n202), .A2(new_n193), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n196), .A2(G146), .A3(new_n197), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n546), .A2(new_n547), .A3(new_n550), .A4(new_n537), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n541), .A2(new_n543), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n543), .B1(new_n541), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n189), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G475), .ZN(new_n555));
  OR2_X1    g369(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n556));
  NAND2_X1  g370(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n202), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n196), .A2(KEYINPUT19), .A3(new_n197), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n193), .A3(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n535), .A2(new_n296), .A3(new_n536), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n522), .B(new_n560), .C1(new_n561), .C2(new_n539), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n551), .ZN(new_n563));
  INV_X1    g377(.A(new_n543), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT87), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n541), .A2(new_n543), .A3(new_n551), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(KEYINPUT87), .A3(new_n564), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT20), .ZN(new_n571));
  NOR2_X1   g385(.A1(G475), .A2(G902), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n571), .B1(new_n570), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n555), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n206), .A2(G143), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n276), .A2(G128), .ZN(new_n577));
  OR3_X1    g391(.A1(new_n576), .A2(new_n577), .A3(G134), .ZN(new_n578));
  INV_X1    g392(.A(G122), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G116), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n258), .A2(G122), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n580), .A2(new_n581), .A3(new_n385), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n385), .B1(new_n580), .B2(new_n581), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n276), .A2(G128), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n577), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n576), .A2(KEYINPUT13), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n287), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT89), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n588), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G134), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT89), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n582), .A2(new_n583), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n578), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT90), .B1(new_n581), .B2(KEYINPUT14), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n581), .A2(KEYINPUT14), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n580), .A3(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n581), .A2(KEYINPUT90), .A3(KEYINPUT14), .ZN(new_n599));
  OAI21_X1  g413(.A(G107), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(G134), .B1(new_n576), .B2(new_n577), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n582), .B1(new_n578), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n590), .A2(new_n595), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT9), .B(G234), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n605), .A2(new_n188), .A3(G953), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n590), .A2(new_n595), .A3(new_n603), .A4(new_n606), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT91), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G478), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(KEYINPUT15), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n610), .B(new_n611), .C1(KEYINPUT15), .C2(new_n613), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n575), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(G221), .B1(new_n605), .B2(G902), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n452), .A2(new_n515), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n375), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  AND3_X1   g437(.A1(new_n452), .A2(new_n515), .A3(new_n619), .ZN(new_n624));
  INV_X1    g438(.A(G472), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n354), .B2(new_n189), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n338), .A2(new_n344), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n347), .B1(new_n627), .B2(new_n349), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n626), .A2(new_n628), .A3(new_n257), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n608), .A2(new_n609), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n630), .A2(KEYINPUT33), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(KEYINPUT33), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(G478), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n613), .A2(new_n189), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n610), .B2(new_n613), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n575), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n624), .A2(new_n629), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NAND3_X1  g455(.A1(new_n452), .A2(new_n515), .A3(new_n619), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n345), .B2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n354), .A2(new_n346), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n252), .A2(new_n256), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT93), .B1(new_n573), .B2(new_n574), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT87), .B1(new_n563), .B2(new_n564), .ZN(new_n648));
  AOI211_X1 g462(.A(new_n566), .B(new_n543), .C1(new_n562), .C2(new_n551), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n552), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n572), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT20), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT93), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n647), .A2(new_n655), .A3(new_n555), .A4(new_n617), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n642), .A2(new_n646), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT35), .B(G107), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NOR2_X1   g473(.A1(new_n239), .A2(KEYINPUT36), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT94), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n230), .A2(new_n662), .A3(new_n233), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n662), .B1(new_n230), .B2(new_n233), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n665), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n660), .A3(new_n663), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n249), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT95), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n669), .A2(KEYINPUT95), .A3(new_n249), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n255), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n643), .A2(new_n644), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n620), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT37), .B(G110), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT96), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n676), .B(new_n678), .ZN(G12));
  INV_X1    g493(.A(new_n674), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n357), .B2(new_n374), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n454), .B1(new_n510), .B2(new_n514), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n452), .A2(new_n619), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n647), .A2(new_n555), .A3(new_n655), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n458), .B(KEYINPUT97), .Z(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n686), .B1(new_n687), .B2(new_n462), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n684), .A2(KEYINPUT98), .A3(new_n617), .A4(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT98), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(new_n656), .B2(new_n688), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n681), .A2(new_n682), .A3(new_n683), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  NOR2_X1   g509(.A1(new_n334), .A2(new_n337), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n326), .B1(new_n367), .B2(new_n371), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT100), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n625), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n369), .A2(new_n370), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n319), .A2(new_n363), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n316), .A2(KEYINPUT69), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n336), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT100), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n696), .A2(new_n699), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(G472), .A2(G902), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT101), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT101), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n706), .A2(new_n710), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n712), .A2(new_n357), .A3(KEYINPUT102), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT102), .B1(new_n712), .B2(new_n357), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n510), .A2(new_n514), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n680), .A2(new_n575), .A3(new_n617), .A4(new_n453), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n688), .B(KEYINPUT39), .Z(new_n721));
  NAND3_X1  g535(.A1(new_n452), .A2(new_n619), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT40), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n452), .A2(new_n724), .A3(new_n619), .A4(new_n721), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n720), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n715), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n276), .ZN(G45));
  NOR2_X1   g542(.A1(new_n637), .A2(new_n688), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n681), .A2(new_n682), .A3(new_n683), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  NOR3_X1   g545(.A1(new_n345), .A2(KEYINPUT32), .A3(new_n347), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n355), .B1(new_n354), .B2(new_n346), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n374), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n448), .A2(new_n619), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n189), .B1(new_n446), .B2(new_n447), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n441), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI211_X1 g552(.A(KEYINPUT103), .B(new_n189), .C1(new_n446), .C2(new_n447), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n735), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n463), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n682), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n637), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n734), .A2(new_n645), .A3(new_n740), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NOR2_X1   g560(.A1(new_n742), .A2(new_n656), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n734), .A2(new_n645), .A3(new_n740), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT104), .B(G116), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G18));
  NAND2_X1  g564(.A1(new_n618), .A2(new_n741), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT105), .B1(new_n740), .B2(new_n682), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n436), .B1(new_n421), .B2(new_n426), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n447), .B1(new_n754), .B2(new_n380), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n737), .B1(new_n755), .B2(G902), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(G469), .A3(new_n739), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n448), .A2(new_n619), .ZN(new_n758));
  AND4_X1   g572(.A1(KEYINPUT105), .A2(new_n757), .A3(new_n682), .A4(new_n758), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n681), .B(new_n752), .C1(new_n753), .C2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G119), .ZN(G21));
  OAI21_X1  g575(.A(KEYINPUT106), .B1(new_n372), .B2(new_n320), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT28), .B1(new_n700), .B2(new_n703), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n764));
  INV_X1    g578(.A(new_n320), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n766), .A3(new_n336), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n347), .B1(new_n767), .B2(new_n627), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n248), .A2(new_n251), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n626), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n652), .A2(new_n654), .B1(G475), .B2(new_n554), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n615), .A2(new_n616), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n575), .A2(new_n617), .A3(KEYINPUT107), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(new_n515), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n771), .A2(new_n778), .A3(KEYINPUT108), .A4(new_n740), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n777), .A2(new_n757), .A3(new_n515), .A4(new_n758), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n767), .A2(new_n627), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n346), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n643), .A3(new_n769), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n780), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G122), .ZN(G24));
  AND4_X1   g601(.A1(new_n643), .A2(new_n783), .A3(new_n729), .A4(new_n674), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(new_n753), .B2(new_n759), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G125), .ZN(G27));
  NAND2_X1  g604(.A1(new_n734), .A2(new_n769), .ZN(new_n791));
  INV_X1    g605(.A(new_n619), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n454), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n510), .A2(new_n514), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n414), .A2(new_n418), .B1(new_n433), .B2(new_n434), .ZN(new_n796));
  INV_X1    g610(.A(new_n438), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT109), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT109), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n437), .A2(new_n799), .A3(new_n438), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n427), .A3(new_n800), .A4(G469), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n441), .A2(new_n189), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT110), .B1(new_n805), .B2(new_n448), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n448), .A2(KEYINPUT110), .A3(new_n803), .A4(new_n801), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n729), .B(new_n795), .C1(new_n806), .C2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT42), .B1(new_n791), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n811));
  INV_X1    g625(.A(new_n448), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(new_n812), .B2(new_n804), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n794), .B1(new_n813), .B2(new_n807), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n637), .A2(KEYINPUT42), .A3(new_n688), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n375), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g631(.A(KEYINPUT111), .B(G131), .Z(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(G33));
  NAND4_X1  g633(.A1(new_n693), .A2(new_n814), .A3(new_n734), .A4(new_n645), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G134), .ZN(G36));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n427), .A2(new_n439), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT45), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n798), .A2(new_n427), .A3(new_n800), .A4(KEYINPUT45), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n822), .A2(new_n825), .A3(G469), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n441), .B1(new_n823), .B2(new_n824), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n822), .B1(new_n828), .B2(new_n826), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n803), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT46), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n448), .ZN(new_n833));
  OAI211_X1 g647(.A(KEYINPUT46), .B(new_n803), .C1(new_n827), .C2(new_n829), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n619), .B(new_n721), .C1(new_n833), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n626), .A2(new_n628), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n633), .A2(new_n635), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n575), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT43), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT43), .B1(new_n575), .B2(new_n838), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n674), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT44), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n837), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n837), .B2(new_n843), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n716), .A2(new_n454), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n836), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n284), .ZN(G39));
  NAND3_X1  g664(.A1(new_n729), .A2(new_n257), .A3(new_n847), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n734), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(KEYINPUT47), .B(new_n619), .C1(new_n833), .C2(new_n835), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n812), .B1(new_n830), .B2(new_n831), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n792), .B1(new_n855), .B2(new_n834), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(KEYINPUT47), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n852), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(G140), .ZN(G42));
  NAND4_X1  g673(.A1(new_n718), .A2(new_n769), .A3(new_n793), .A4(new_n839), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT49), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n757), .A2(new_n448), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n860), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n864), .B(new_n715), .C1(new_n861), .C2(new_n863), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n689), .A2(new_n619), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n674), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n777), .A2(new_n868), .A3(new_n682), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n813), .B2(new_n807), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n713), .B2(new_n714), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n694), .A3(new_n730), .A4(new_n789), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT52), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n773), .A2(new_n617), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n642), .A2(new_n646), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n875), .A2(new_n876), .A3(new_n676), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n620), .A2(new_n675), .ZN(new_n878));
  INV_X1    g692(.A(new_n874), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n624), .A2(new_n629), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT113), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n786), .A2(new_n760), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n622), .A2(new_n744), .A3(new_n748), .A4(new_n639), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n617), .A2(new_n688), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n847), .A2(new_n684), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n734), .A2(new_n683), .A3(new_n887), .A4(new_n674), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n788), .A2(new_n814), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n820), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n817), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n873), .A2(new_n882), .A3(new_n885), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n872), .A2(KEYINPUT52), .ZN(new_n894));
  OR4_X1    g708(.A1(new_n866), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n814), .A2(new_n734), .A3(new_n645), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n814), .A2(new_n734), .A3(new_n769), .A4(new_n729), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n897), .A2(new_n815), .B1(new_n898), .B2(KEYINPUT42), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n820), .A2(new_n888), .A3(new_n889), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n877), .A2(new_n881), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n642), .A2(new_n646), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n638), .A2(new_n903), .B1(new_n375), .B2(new_n621), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n375), .B(new_n740), .C1(new_n743), .C2(new_n747), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n786), .A3(new_n760), .A4(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n901), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n894), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n907), .A2(KEYINPUT53), .A3(new_n908), .A4(new_n873), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n896), .A2(new_n909), .A3(new_n866), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n895), .A2(KEYINPUT54), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n896), .A2(new_n909), .A3(KEYINPUT115), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n913), .B(new_n893), .C1(new_n892), .C2(new_n894), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n911), .B1(new_n915), .B2(KEYINPUT54), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n854), .A2(new_n857), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n863), .A2(new_n792), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n919), .A2(KEYINPUT119), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n841), .A2(new_n686), .A3(new_n842), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n784), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n922), .A2(new_n847), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n919), .A2(KEYINPUT119), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n740), .A2(new_n847), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n926), .A2(new_n257), .A3(new_n458), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n715), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n928), .A2(KEYINPUT118), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(KEYINPUT118), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n773), .A3(new_n838), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n926), .A2(new_n921), .ZN(new_n933));
  NOR4_X1   g747(.A1(new_n933), .A2(new_n626), .A3(new_n680), .A4(new_n768), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT50), .ZN(new_n935));
  INV_X1    g749(.A(new_n922), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n718), .A2(new_n740), .A3(new_n454), .ZN(new_n937));
  OAI211_X1 g751(.A(KEYINPUT117), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n937), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n935), .A2(KEYINPUT117), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n922), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n934), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n925), .A2(KEYINPUT51), .A3(new_n932), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n933), .A2(new_n791), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT48), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n753), .A2(new_n759), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n455), .B1(new_n947), .B2(new_n936), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n945), .B(new_n948), .C1(new_n931), .C2(new_n638), .ZN(new_n949));
  XNOR2_X1  g763(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n932), .A2(new_n942), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n919), .A2(new_n923), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n943), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n916), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(G952), .A2(G953), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n865), .B1(new_n955), .B2(new_n956), .ZN(G75));
  NAND4_X1  g771(.A1(new_n912), .A2(G210), .A3(G902), .A4(new_n914), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n479), .A2(new_n492), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n490), .ZN(new_n960));
  XNOR2_X1  g774(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g776(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n958), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT56), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n236), .A2(G952), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(G51));
  XNOR2_X1  g782(.A(new_n802), .B(KEYINPUT57), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n912), .A2(KEYINPUT54), .A3(new_n914), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT54), .B1(new_n912), .B2(new_n914), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n755), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n912), .A2(new_n914), .ZN(new_n975));
  OR4_X1    g789(.A1(new_n189), .A2(new_n975), .A3(new_n827), .A4(new_n829), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n967), .B1(new_n974), .B2(new_n976), .ZN(G54));
  AND2_X1   g791(.A1(KEYINPUT58), .A2(G475), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n912), .A2(G902), .A3(new_n914), .A4(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(new_n650), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n650), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n980), .A2(new_n981), .A3(new_n967), .ZN(G60));
  NAND2_X1  g796(.A1(new_n631), .A2(new_n632), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n634), .B(KEYINPUT59), .Z(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n916), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n970), .B2(new_n971), .ZN(new_n987));
  INV_X1    g801(.A(new_n967), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n985), .A2(new_n989), .ZN(G63));
  XNOR2_X1  g804(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n188), .A2(new_n189), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n242), .B1(new_n975), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n912), .A2(new_n669), .A3(new_n914), .A4(new_n993), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n988), .A3(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT61), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n995), .A2(KEYINPUT61), .A3(new_n988), .A4(new_n996), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(G66));
  INV_X1    g815(.A(new_n460), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n236), .B1(new_n1002), .B2(G224), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n882), .A2(new_n885), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n236), .ZN(new_n1005));
  INV_X1    g819(.A(G898), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n959), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1005), .B(new_n1007), .ZN(G69));
  INV_X1    g822(.A(KEYINPUT124), .ZN(new_n1009));
  AOI211_X1 g823(.A(new_n454), .B(new_n716), .C1(new_n637), .C2(new_n874), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n375), .A2(new_n683), .A3(new_n721), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(new_n836), .B2(new_n848), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n856), .B(KEYINPUT47), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(new_n852), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n789), .A2(new_n694), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n720), .A2(new_n723), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1016), .B(new_n725), .C1(new_n714), .C2(new_n713), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1015), .A2(new_n1017), .A3(KEYINPUT62), .A4(new_n730), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT62), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n694), .A2(new_n789), .A3(new_n730), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1019), .B1(new_n1020), .B2(new_n727), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1014), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT123), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1014), .A2(new_n1022), .A3(KEYINPUT123), .ZN(new_n1026));
  AOI21_X1  g840(.A(G953), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n558), .A2(new_n559), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n332), .B(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1009), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1026), .ZN(new_n1031));
  AOI21_X1  g845(.A(KEYINPUT123), .B1(new_n1014), .B2(new_n1022), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n236), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1029), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1033), .A2(KEYINPUT124), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n236), .B1(G227), .B2(G900), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1034), .B1(G900), .B2(G953), .ZN(new_n1038));
  AND4_X1   g852(.A1(new_n734), .A2(new_n769), .A3(new_n682), .A4(new_n777), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n856), .A2(new_n721), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(KEYINPUT125), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT125), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n856), .A2(new_n1042), .A3(new_n721), .A4(new_n1039), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n810), .A2(new_n816), .A3(new_n820), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n849), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1020), .ZN(new_n1047));
  NAND4_X1  g861(.A1(new_n1044), .A2(new_n1046), .A3(new_n858), .A4(new_n1047), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1038), .B1(new_n1048), .B2(G953), .ZN(new_n1049));
  NAND4_X1  g863(.A1(new_n1030), .A2(new_n1035), .A3(new_n1037), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT126), .ZN(new_n1051));
  XNOR2_X1  g865(.A(new_n1049), .B(new_n1051), .ZN(new_n1052));
  AND3_X1   g866(.A1(new_n1030), .A2(new_n1052), .A3(new_n1035), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1050), .B1(new_n1053), .B2(new_n1037), .ZN(G72));
  XNOR2_X1  g868(.A(new_n707), .B(KEYINPUT63), .ZN(new_n1055));
  INV_X1    g869(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1056), .B1(new_n1048), .B2(new_n1004), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n1057), .B(KEYINPUT127), .ZN(new_n1058));
  AND3_X1   g872(.A1(new_n1058), .A2(new_n336), .A3(new_n333), .ZN(new_n1059));
  NAND4_X1  g873(.A1(new_n1025), .A2(new_n882), .A3(new_n885), .A4(new_n1026), .ZN(new_n1060));
  AOI211_X1 g874(.A(new_n336), .B(new_n333), .C1(new_n1060), .C2(new_n1056), .ZN(new_n1061));
  INV_X1    g875(.A(new_n361), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1055), .B1(new_n696), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n895), .A2(new_n910), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1064), .A2(new_n988), .ZN(new_n1065));
  NOR3_X1   g879(.A1(new_n1059), .A2(new_n1061), .A3(new_n1065), .ZN(G57));
endmodule


