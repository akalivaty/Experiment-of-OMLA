//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(G902), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G110), .B(G140), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G227), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n194), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G137), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT11), .A3(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G131), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n201), .A2(new_n203), .A3(new_n207), .A4(new_n204), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(G143), .B2(new_n210), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n211), .A2(new_n213), .A3(new_n215), .A4(G128), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT74), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT74), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G107), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G104), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G107), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n226), .A2(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n222), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n229), .A2(G107), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n227), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G101), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT10), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT10), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n220), .A2(new_n234), .A3(new_n240), .A4(new_n237), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n230), .B1(new_n222), .B2(new_n224), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n227), .A2(new_n235), .B1(new_n221), .B2(KEYINPUT3), .ZN(new_n243));
  OAI21_X1  g057(.A(G101), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n234), .A3(KEYINPUT4), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT75), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT75), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n244), .A2(new_n234), .A3(new_n247), .A4(KEYINPUT4), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n211), .A2(new_n213), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT0), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n217), .A3(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(KEYINPUT0), .B2(G128), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n255), .B2(new_n250), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n251), .B1(new_n214), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n259), .B(G101), .C1(new_n242), .C2(new_n243), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT76), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n228), .A2(new_n232), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT76), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n259), .A4(G101), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n258), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  AOI221_X4 g079(.A(new_n209), .B1(new_n239), .B2(new_n241), .C1(new_n249), .C2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n209), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n227), .A2(new_n225), .B1(new_n236), .B2(new_n222), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n259), .B1(new_n268), .B2(new_n233), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n247), .B1(new_n269), .B2(new_n244), .ZN(new_n270));
  INV_X1    g084(.A(new_n248), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n265), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n239), .A2(new_n241), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n267), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n198), .B1(new_n266), .B2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n220), .A2(new_n234), .A3(new_n237), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n220), .B1(new_n234), .B2(new_n237), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n209), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT12), .B(new_n209), .C1(new_n276), .C2(new_n277), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(KEYINPUT77), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n272), .A2(new_n267), .A3(new_n273), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT77), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n278), .A2(new_n284), .A3(new_n279), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n282), .A2(new_n283), .A3(new_n197), .A4(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(G902), .B1(new_n275), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n193), .B1(new_n287), .B2(new_n191), .ZN(new_n288));
  OR3_X1    g102(.A1(new_n266), .A2(new_n274), .A3(new_n198), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n198), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n291), .A3(G469), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n190), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n212), .A2(G128), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT84), .B1(new_n217), .B2(G143), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT84), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(new_n212), .A3(G128), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(new_n200), .ZN(new_n300));
  INV_X1    g114(.A(G116), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G122), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT14), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT14), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n301), .A3(G122), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n301), .A2(G122), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT85), .A3(G107), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n226), .A3(new_n302), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(G107), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT85), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n300), .A2(new_n308), .A3(new_n309), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n299), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n295), .A2(KEYINPUT13), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(new_n200), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n306), .A2(new_n302), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G107), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n314), .A2(new_n316), .B1(new_n318), .B2(new_n309), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n314), .B2(new_n316), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n187), .A2(G217), .A3(new_n195), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n322), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n313), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n192), .ZN(new_n327));
  INV_X1    g141(.A(G478), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT15), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n326), .B(new_n192), .C1(KEYINPUT15), .C2(new_n328), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(G475), .A2(G902), .ZN(new_n335));
  INV_X1    g149(.A(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G125), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G140), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT16), .ZN(new_n340));
  OR3_X1    g154(.A1(new_n338), .A2(KEYINPUT16), .A3(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n210), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n341), .A3(G146), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT69), .A4(G146), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G237), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n195), .A3(G214), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(new_n212), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT17), .A3(G131), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(G131), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n350), .B(G143), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n207), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT17), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n348), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G113), .B(G122), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT82), .B(G104), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT18), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n354), .B1(new_n363), .B2(new_n207), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n351), .A2(KEYINPUT18), .A3(G131), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n337), .A2(new_n339), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(new_n210), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n358), .A2(new_n362), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n366), .B(KEYINPUT19), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n210), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n353), .A2(new_n355), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n345), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n362), .B1(new_n374), .B2(new_n368), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n335), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT20), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n362), .B1(new_n358), .B2(new_n368), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n192), .B1(new_n370), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT83), .B(new_n192), .C1(new_n370), .C2(new_n378), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G475), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n334), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n195), .A2(G952), .ZN(new_n387));
  NAND2_X1  g201(.A1(G234), .A2(G237), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(KEYINPUT87), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT21), .B(G898), .Z(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n388), .A2(G902), .A3(G953), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(G214), .B1(G237), .B2(G902), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n396), .B(KEYINPUT78), .Z(new_n397));
  AND2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G210), .B1(G237), .B2(G902), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT81), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G116), .B(G119), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT2), .B(G113), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT2), .B(G113), .Z(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n402), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n261), .B2(new_n264), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n249), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n402), .A2(KEYINPUT5), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n301), .A2(KEYINPUT5), .A3(G119), .ZN(new_n413));
  INV_X1    g227(.A(G113), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n412), .A2(new_n415), .B1(new_n406), .B2(new_n402), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n234), .A3(new_n237), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G122), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT79), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(KEYINPUT6), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n417), .ZN(new_n424));
  AOI211_X1 g238(.A(new_n424), .B(new_n420), .C1(new_n249), .C2(new_n410), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n249), .B2(new_n410), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(new_n421), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G143), .B(G146), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n252), .A2(new_n217), .ZN(new_n432));
  NAND2_X1  g246(.A1(KEYINPUT0), .A2(G128), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n254), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n431), .B1(new_n434), .B2(new_n253), .ZN(new_n435));
  OAI21_X1  g249(.A(G125), .B1(new_n435), .B2(new_n251), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n218), .A2(new_n338), .A3(new_n219), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n195), .A2(G224), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n438), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n430), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(KEYINPUT7), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n256), .A2(new_n214), .ZN(new_n444));
  INV_X1    g258(.A(new_n251), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n338), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n218), .A2(new_n338), .A3(new_n219), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n436), .A2(KEYINPUT7), .A3(new_n437), .A4(new_n439), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n234), .A2(new_n237), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n412), .A2(new_n415), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n407), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT80), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n454), .A2(new_n417), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n416), .A2(new_n234), .A3(KEYINPUT80), .A4(new_n237), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n419), .B(KEYINPUT8), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n450), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n192), .B1(new_n425), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n401), .B1(new_n442), .B2(new_n461), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n400), .B(new_n460), .C1(new_n430), .C2(new_n441), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n398), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n294), .A2(new_n386), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n209), .A2(new_n257), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n200), .A2(G137), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n202), .A2(G134), .ZN(new_n468));
  OAI21_X1  g282(.A(G131), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n208), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n220), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n466), .A2(new_n471), .A3(KEYINPUT30), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n408), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n349), .A2(new_n195), .A3(G210), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(G101), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n209), .A2(new_n257), .B1(new_n470), .B2(new_n220), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n409), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n476), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n466), .A2(new_n409), .A3(new_n471), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n409), .B1(new_n466), .B2(new_n471), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT28), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT28), .B1(new_n481), .B2(new_n409), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n480), .B(KEYINPUT65), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI22_X1  g305(.A1(KEYINPUT31), .A2(new_n483), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT31), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n476), .A2(new_n493), .A3(new_n480), .A4(new_n482), .ZN(new_n494));
  AOI21_X1  g308(.A(G902), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G472), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT32), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n483), .A2(KEYINPUT31), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n489), .A2(new_n491), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n494), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n500), .A2(KEYINPUT32), .A3(new_n496), .A4(new_n192), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n480), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n466), .A2(KEYINPUT30), .A3(new_n471), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT30), .B1(new_n466), .B2(new_n471), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n504), .A2(new_n505), .A3(new_n409), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n503), .B1(new_n506), .B2(new_n484), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT66), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n472), .A2(new_n408), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n482), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n487), .B1(new_n511), .B2(KEYINPUT28), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT29), .B1(new_n512), .B2(new_n490), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n476), .A2(new_n482), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(KEYINPUT66), .A3(new_n503), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n509), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n480), .A2(KEYINPUT29), .ZN(new_n517));
  AOI21_X1  g331(.A(G902), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n496), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n497), .A2(new_n502), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G234), .ZN(new_n521));
  OAI21_X1  g335(.A(G217), .B1(new_n521), .B2(G902), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT67), .Z(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT71), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT22), .B(G137), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OR2_X1    g343(.A1(KEYINPUT24), .A2(G110), .ZN(new_n530));
  INV_X1    g344(.A(G119), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G128), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n217), .A2(G119), .ZN(new_n533));
  NAND2_X1  g347(.A1(KEYINPUT24), .A2(G110), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n530), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(KEYINPUT24), .A2(G110), .ZN(new_n538));
  NOR2_X1   g352(.A1(KEYINPUT24), .A2(G110), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n540), .A2(KEYINPUT68), .A3(new_n532), .A4(new_n533), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(G119), .B2(new_n217), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n531), .A2(KEYINPUT23), .A3(G128), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n532), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n537), .A2(new_n541), .B1(new_n545), .B2(G110), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n346), .A2(new_n546), .A3(new_n347), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n366), .A2(new_n210), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n545), .A2(G110), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n540), .B1(new_n532), .B2(new_n533), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n345), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n548), .B1(new_n547), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n529), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n547), .A2(new_n552), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(new_n529), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n192), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT25), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n555), .A2(KEYINPUT25), .A3(new_n558), .A4(new_n192), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n524), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n556), .A2(KEYINPUT70), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n557), .B1(new_n566), .B2(new_n529), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n522), .A2(new_n192), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n568), .B(KEYINPUT72), .Z(new_n569));
  AND2_X1   g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT73), .B1(new_n563), .B2(new_n570), .ZN(new_n571));
  OR3_X1    g385(.A1(new_n563), .A2(KEYINPUT73), .A3(new_n570), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n520), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n465), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT88), .B(G101), .Z(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(G3));
  INV_X1    g390(.A(new_n396), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT89), .B1(new_n462), .B2(new_n463), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n460), .B1(new_n430), .B2(new_n441), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n401), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n577), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n313), .B(new_n320), .C1(KEYINPUT91), .C2(new_n324), .ZN(new_n583));
  OAI211_X1 g397(.A(KEYINPUT33), .B(new_n583), .C1(new_n323), .C2(KEYINPUT91), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n328), .A2(G902), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT90), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n326), .B2(new_n587), .ZN(new_n588));
  AOI211_X1 g402(.A(KEYINPUT90), .B(KEYINPUT33), .C1(new_n323), .C2(new_n325), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n584), .B(new_n585), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n327), .A2(new_n328), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n377), .A2(new_n383), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n582), .A2(new_n395), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n496), .B1(new_n500), .B2(new_n192), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n500), .A2(new_n496), .A3(new_n192), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n572), .B2(new_n571), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n293), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT34), .B(G104), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  NOR2_X1   g416(.A1(new_n334), .A2(new_n384), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n582), .A2(new_n395), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n599), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT35), .B(G107), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G9));
  AOI21_X1  g421(.A(KEYINPUT25), .B1(new_n567), .B2(new_n192), .ZN(new_n608));
  INV_X1    g422(.A(new_n562), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n523), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT93), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n528), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT92), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n566), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n613), .A2(KEYINPUT92), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(KEYINPUT92), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(new_n564), .A3(new_n565), .A4(new_n617), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n615), .A2(new_n569), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n610), .A2(new_n611), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT93), .B1(new_n563), .B2(new_n619), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n597), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n465), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  NOR2_X1   g441(.A1(new_n520), .A2(new_n623), .ZN(new_n628));
  INV_X1    g442(.A(G900), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT94), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n629), .A2(KEYINPUT94), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n393), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n390), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT95), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n334), .A2(new_n384), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n628), .A2(new_n582), .A3(new_n293), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  XNOR2_X1  g451(.A(new_n580), .B(new_n401), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n638), .B(new_n639), .Z(new_n640));
  NOR3_X1   g454(.A1(new_n334), .A2(new_n385), .A3(new_n577), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT32), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n596), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n491), .A2(new_n511), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n644), .A2(new_n483), .ZN(new_n645));
  OAI21_X1  g459(.A(G472), .B1(new_n645), .B2(G902), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n643), .A2(new_n501), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n640), .A2(new_n623), .A3(new_n641), .A4(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT97), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n634), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n293), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT40), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(new_n212), .ZN(G45));
  INV_X1    g471(.A(new_n634), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n592), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n628), .A2(new_n582), .A3(new_n293), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  NAND2_X1  g476(.A1(new_n275), .A2(new_n286), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n192), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(G469), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n287), .B2(new_n191), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n664), .A2(new_n666), .A3(G469), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n189), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n190), .B1(new_n668), .B2(new_n669), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n593), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n676), .A2(new_n677), .A3(KEYINPUT101), .A4(new_n573), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT100), .B1(new_n670), .B2(new_n189), .ZN(new_n680));
  AOI211_X1 g494(.A(new_n672), .B(new_n190), .C1(new_n668), .C2(new_n669), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n573), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n679), .B1(new_n682), .B2(new_n593), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n687), .B1(new_n682), .B2(new_n604), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n582), .A2(new_n395), .A3(new_n603), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n676), .A2(new_n689), .A3(KEYINPUT102), .A4(new_n573), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  INV_X1    g506(.A(new_n395), .ZN(new_n693));
  NOR4_X1   g507(.A1(new_n520), .A2(new_n386), .A3(new_n623), .A4(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n582), .A2(new_n674), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n500), .A2(new_n496), .A3(new_n192), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n698), .B1(new_n699), .B2(new_n594), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n595), .A2(KEYINPUT103), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n563), .A2(new_n570), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n703), .A3(new_n395), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n578), .A2(new_n581), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n641), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n676), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT104), .B(G122), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G24));
  AND4_X1   g524(.A1(new_n622), .A2(new_n700), .A3(new_n701), .A4(new_n621), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n582), .A3(new_n660), .A4(new_n674), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT105), .B(G125), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G27));
  NAND2_X1  g528(.A1(new_n289), .A2(new_n291), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT106), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n289), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n716), .A2(G469), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n190), .B1(new_n719), .B2(new_n288), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n462), .A2(new_n463), .A3(new_n577), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n659), .A2(KEYINPUT42), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n573), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n720), .A2(new_n660), .A3(new_n721), .ZN(new_n726));
  INV_X1    g540(.A(new_n520), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n703), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT42), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n207), .ZN(G33));
  NAND3_X1  g545(.A1(new_n723), .A2(new_n573), .A3(new_n635), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  NAND2_X1  g547(.A1(new_n590), .A2(new_n591), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n384), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT43), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(KEYINPUT43), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n623), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n597), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n721), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n716), .A2(KEYINPUT45), .A3(new_n718), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n746), .A2(KEYINPUT107), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n289), .A2(new_n291), .ZN(new_n748));
  OAI21_X1  g562(.A(G469), .B1(new_n748), .B2(KEYINPUT45), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(new_n746), .B2(KEYINPUT107), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n193), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n752), .A2(KEYINPUT46), .B1(new_n191), .B2(new_n287), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n190), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n653), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT108), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n758), .A3(new_n653), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n745), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n202), .ZN(G39));
  NAND2_X1  g575(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n287), .A2(new_n191), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n189), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT47), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n755), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n572), .A2(new_n571), .ZN(new_n770));
  AND4_X1   g584(.A1(new_n520), .A2(new_n770), .A3(new_n660), .A4(new_n721), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n767), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n390), .B1(new_n737), .B2(new_n738), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n674), .A2(new_n775), .A3(new_n711), .A4(new_n721), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n640), .A2(new_n396), .A3(new_n671), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n703), .A3(new_n702), .ZN(new_n778));
  NOR2_X1   g592(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n779), .B1(new_n777), .B2(new_n778), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n674), .A2(new_n721), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n783), .A2(new_n770), .A3(new_n390), .A4(new_n647), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n385), .A3(new_n735), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT116), .Z(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT117), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n767), .A2(new_n769), .B1(new_n190), .B2(new_n670), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n778), .A2(new_n638), .A3(new_n577), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT114), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n789), .A2(KEYINPUT114), .A3(new_n791), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n774), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n782), .A2(KEYINPUT51), .A3(new_n786), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n789), .B2(new_n791), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT118), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n796), .B(new_n799), .C1(new_n789), .C2(new_n791), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n775), .A2(new_n674), .A3(new_n721), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n728), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT48), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(KEYINPUT48), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n784), .A2(new_n592), .ZN(new_n805));
  INV_X1    g619(.A(new_n695), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n805), .B(new_n387), .C1(new_n806), .C2(new_n778), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n798), .A2(new_n800), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n795), .A2(new_n809), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n707), .A2(new_n676), .B1(new_n694), .B2(new_n695), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n725), .A2(new_n732), .A3(new_n729), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n684), .A2(new_n691), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n711), .A2(new_n660), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n332), .A2(new_n634), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n293), .A2(new_n721), .A3(new_n385), .A4(new_n816), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n815), .A2(new_n723), .B1(new_n817), .B2(new_n628), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n465), .B1(new_n573), .B2(new_n624), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n385), .A2(new_n332), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n464), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n598), .A2(new_n821), .A3(new_n293), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n592), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT111), .B1(new_n824), .B2(new_n464), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n638), .A2(new_n826), .A3(new_n398), .A4(new_n592), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n825), .A2(new_n827), .A3(new_n293), .A4(new_n598), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n818), .A2(new_n819), .A3(new_n823), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n636), .A2(new_n712), .A3(new_n661), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n563), .A2(new_n619), .A3(new_n634), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n647), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n641), .A2(new_n833), .A3(new_n705), .A4(new_n720), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(KEYINPUT52), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n636), .A2(new_n712), .A3(new_n661), .A4(new_n834), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n829), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n813), .A2(new_n839), .B1(KEYINPUT112), .B2(KEYINPUT53), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(KEYINPUT112), .B2(KEYINPUT53), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n819), .A2(new_n828), .A3(new_n823), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n817), .A2(new_n628), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n814), .B2(new_n722), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n836), .A2(new_n837), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n836), .A2(new_n837), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n684), .A2(new_n691), .A3(new_n811), .A4(new_n812), .ZN(new_n849));
  OR4_X1    g663(.A1(KEYINPUT112), .A2(new_n848), .A3(new_n849), .A4(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n841), .A2(new_n850), .A3(KEYINPUT54), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n732), .A2(KEYINPUT113), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n813), .B(new_n839), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n845), .B(new_n853), .C1(new_n846), .C2(new_n847), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n855), .B(KEYINPUT53), .C1(new_n848), .C2(new_n849), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n851), .A2(new_n859), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n810), .A2(new_n860), .B1(G952), .B2(G953), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n640), .A2(new_n647), .ZN(new_n862));
  INV_X1    g676(.A(new_n670), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT49), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n736), .A2(new_n189), .A3(new_n397), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n703), .A3(new_n865), .ZN(new_n866));
  OAI221_X1 g680(.A(new_n862), .B1(KEYINPUT49), .B2(new_n863), .C1(KEYINPUT109), .C2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(KEYINPUT109), .B2(new_n866), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT110), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n861), .A2(new_n869), .ZN(G75));
  NOR2_X1   g684(.A1(new_n857), .A2(new_n192), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT56), .B1(new_n871), .B2(new_n400), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n430), .B(new_n441), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT55), .Z(new_n874));
  AND2_X1   g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n872), .A2(new_n874), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n195), .A2(G952), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G51));
  NAND2_X1  g692(.A1(new_n871), .A2(new_n751), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n663), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n193), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n854), .A2(new_n856), .A3(KEYINPUT54), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT54), .B1(new_n854), .B2(new_n856), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(KEYINPUT120), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n880), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT121), .B1(new_n890), .B2(new_n877), .ZN(new_n891));
  INV_X1    g705(.A(new_n883), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n854), .A2(new_n856), .A3(KEYINPUT54), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n859), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n663), .B1(new_n894), .B2(KEYINPUT120), .ZN(new_n895));
  INV_X1    g709(.A(new_n889), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n879), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n898));
  INV_X1    g712(.A(new_n877), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n891), .A2(new_n900), .ZN(G54));
  NAND2_X1  g715(.A1(KEYINPUT58), .A2(G475), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT122), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n871), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n370), .A2(new_n375), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n877), .ZN(G60));
  OR2_X1    g722(.A1(new_n588), .A2(new_n589), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n909), .A2(new_n584), .ZN(new_n910));
  NAND2_X1  g724(.A1(G478), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT59), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n910), .B1(new_n860), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n859), .A2(new_n893), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n910), .A2(new_n912), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n877), .B(new_n913), .C1(new_n914), .C2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT60), .Z(new_n918));
  AND3_X1   g732(.A1(new_n854), .A2(new_n856), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n618), .A3(new_n615), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n920), .B(new_n899), .C1(new_n567), .C2(new_n919), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g736(.A(new_n195), .B1(new_n391), .B2(G224), .ZN(new_n923));
  INV_X1    g737(.A(new_n842), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n684), .A2(new_n691), .A3(new_n924), .A4(new_n811), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n925), .B2(new_n195), .ZN(new_n926));
  INV_X1    g740(.A(G898), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n430), .B1(new_n927), .B2(G953), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n926), .B(new_n928), .ZN(G69));
  NAND2_X1  g743(.A1(new_n474), .A2(new_n475), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(new_n371), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n772), .A2(new_n812), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n757), .A2(new_n759), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n706), .A2(new_n728), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n760), .B2(new_n830), .ZN(new_n938));
  INV_X1    g752(.A(new_n745), .ZN(new_n939));
  INV_X1    g753(.A(new_n759), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n758), .B1(new_n755), .B2(new_n653), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(KEYINPUT124), .A3(new_n831), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n936), .A2(new_n938), .A3(new_n195), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(G900), .A2(G953), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n932), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n948));
  OR3_X1    g762(.A1(new_n656), .A2(new_n830), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n950));
  OAI22_X1  g764(.A1(new_n656), .A2(new_n830), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n573), .B(new_n721), .C1(new_n592), .C2(new_n821), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n952), .A2(new_n654), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n954), .A2(new_n942), .A3(new_n772), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n955), .A2(G953), .A3(new_n931), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n946), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n944), .A2(new_n945), .ZN(new_n959));
  NAND2_X1  g773(.A1(G227), .A2(G900), .ZN(new_n960));
  AND4_X1   g774(.A1(G953), .A2(new_n959), .A3(new_n960), .A4(new_n931), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n958), .A2(new_n961), .ZN(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT63), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n509), .A2(new_n515), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(new_n483), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n841), .A2(new_n850), .A3(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n964), .B(KEYINPUT125), .ZN(new_n968));
  INV_X1    g782(.A(new_n925), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n955), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n514), .A2(new_n480), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n936), .A2(new_n938), .A3(new_n969), .A4(new_n943), .ZN(new_n974));
  INV_X1    g788(.A(new_n968), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n514), .A2(new_n480), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT126), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n973), .B(new_n899), .C1(new_n976), .C2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(new_n974), .B2(new_n975), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT127), .B1(new_n981), .B2(new_n877), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n972), .B1(new_n980), .B2(new_n982), .ZN(G57));
endmodule


