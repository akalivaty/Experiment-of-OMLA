//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G116), .A2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G50), .B2(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n212), .B(new_n228), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n220), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(new_n206), .A2(G20), .ZN(new_n249));
  INV_X1    g0049(.A(G13), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G50), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n203), .A2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(KEYINPUT8), .B(G58), .Z(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT67), .B1(new_n260), .B2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT67), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(new_n207), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n254), .B1(new_n255), .B2(new_n257), .C1(new_n259), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n208), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n229), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n253), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(G1), .A2(G13), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(new_n208), .B2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n249), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n269), .B1(new_n202), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n229), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(G222), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n280), .B(KEYINPUT66), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G223), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n282), .A2(new_n283), .B1(new_n284), .B2(new_n278), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n277), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT64), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n276), .A2(new_n290), .A3(new_n229), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT64), .B1(new_n270), .B2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(G274), .B(new_n289), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(KEYINPUT65), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT65), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n290), .B1(new_n276), .B2(new_n229), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n270), .A2(KEYINPUT64), .A3(new_n292), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n296), .B1(new_n300), .B2(new_n289), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n289), .B1(new_n298), .B2(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G226), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n286), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n275), .B1(G200), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n305), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G190), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT69), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n273), .A2(new_n274), .B1(new_n309), .B2(KEYINPUT10), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n312), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n294), .A2(KEYINPUT65), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n300), .A2(new_n296), .A3(new_n289), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n303), .A2(G238), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G97), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n220), .A2(G1698), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G226), .B2(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n318), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n277), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n315), .A2(new_n316), .A3(new_n317), .A4(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n327), .A2(KEYINPUT13), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(KEYINPUT13), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT14), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(G179), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n302), .A2(new_n334), .A3(new_n317), .A4(new_n326), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n327), .A2(KEYINPUT13), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT14), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(G169), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n332), .A2(new_n333), .A3(new_n339), .ZN(new_n340));
  OR3_X1    g0140(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT12), .B1(new_n252), .B2(G68), .ZN(new_n342));
  INV_X1    g0142(.A(new_n272), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(G68), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n264), .A2(G77), .B1(G50), .B2(new_n256), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n224), .A2(G20), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n271), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT11), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n347), .A2(new_n348), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n340), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n352), .B1(new_n337), .B2(G200), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n335), .A2(G190), .A3(new_n336), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT70), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(G200), .B1(new_n328), .B2(new_n329), .ZN(new_n357));
  INV_X1    g0157(.A(new_n352), .ZN(new_n358));
  AND4_X1   g0158(.A1(KEYINPUT70), .A2(new_n357), .A3(new_n358), .A4(new_n355), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n313), .A2(new_n314), .A3(new_n353), .A4(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n258), .A2(new_n251), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n272), .B2(new_n258), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT73), .B1(new_n256), .B2(G159), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n256), .A2(KEYINPUT73), .A3(G159), .ZN(new_n366));
  XNOR2_X1  g0166(.A(G58), .B(G68), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n365), .A2(new_n366), .B1(G20), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n278), .B2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n324), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT71), .ZN(new_n374));
  OAI21_X1  g0174(.A(G68), .B1(new_n373), .B2(KEYINPUT71), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI211_X1 g0176(.A(new_n371), .B(G20), .C1(new_n321), .C2(new_n323), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT71), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n224), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT71), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(KEYINPUT72), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n369), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n271), .B1(new_n382), .B2(KEYINPUT16), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n224), .B1(new_n372), .B2(new_n373), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n369), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n363), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G223), .A2(G1698), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n279), .A2(G226), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n324), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n260), .A2(new_n215), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n277), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n303), .A2(G232), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n315), .A2(new_n392), .A3(new_n316), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(G200), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n387), .A2(KEYINPUT17), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n379), .A2(KEYINPUT72), .A3(new_n380), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT72), .B1(new_n379), .B2(new_n380), .ZN(new_n400));
  OAI211_X1 g0200(.A(KEYINPUT16), .B(new_n368), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(new_n386), .A3(new_n268), .ZN(new_n402));
  INV_X1    g0202(.A(new_n363), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n402), .A2(new_n396), .A3(new_n403), .A4(new_n397), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n403), .ZN(new_n407));
  INV_X1    g0207(.A(G179), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n394), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n394), .A2(G169), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT18), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  AOI221_X4 g0213(.A(new_n413), .B1(new_n410), .B2(new_n409), .C1(new_n402), .C2(new_n403), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n398), .B(new_n406), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n324), .A2(G107), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n278), .A2(new_n279), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n416), .B1(new_n417), .B2(new_n220), .C1(new_n225), .C2(new_n282), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n277), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n303), .A2(G244), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n302), .A3(new_n420), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n421), .A2(G179), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n252), .A2(G77), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n272), .A2(new_n284), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n258), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n425));
  XOR2_X1   g0225(.A(KEYINPUT15), .B(G87), .Z(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n425), .B1(new_n265), .B2(new_n427), .ZN(new_n428));
  AOI211_X1 g0228(.A(new_n423), .B(new_n424), .C1(new_n428), .C2(new_n268), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n421), .B2(new_n331), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n421), .A2(G200), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n429), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT68), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n421), .A2(new_n395), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n307), .A2(new_n408), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n305), .A2(new_n331), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n273), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR4_X1   g0241(.A1(new_n361), .A2(new_n415), .A3(new_n437), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT6), .ZN(new_n443));
  AND2_X1   g0243(.A1(G97), .A2(G107), .ZN(new_n444));
  NOR2_X1   g0244(.A1(G97), .A2(G107), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n221), .A2(KEYINPUT6), .A3(G97), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n448), .A2(new_n207), .B1(new_n284), .B2(new_n257), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n221), .B1(new_n372), .B2(new_n373), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n268), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT74), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT7), .B1(new_n324), .B2(new_n207), .ZN(new_n454));
  OAI21_X1  g0254(.A(G107), .B1(new_n454), .B2(new_n377), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n446), .A2(new_n447), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n271), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT74), .ZN(new_n459));
  INV_X1    g0259(.A(G97), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n453), .A2(new_n459), .B1(new_n460), .B2(new_n251), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n321), .A2(new_n323), .A3(G244), .A4(new_n279), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT4), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n279), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n277), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n206), .A2(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n472), .A2(KEYINPUT75), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(KEYINPUT75), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n473), .A2(new_n300), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n472), .A2(new_n474), .B1(new_n298), .B2(new_n299), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G257), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n469), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT76), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT76), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n469), .A2(new_n481), .A3(new_n476), .A4(new_n478), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(G200), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n268), .A2(new_n251), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n206), .A2(G33), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G97), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n469), .A2(new_n478), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(G190), .A3(new_n476), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n461), .A2(new_n483), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT24), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n278), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n221), .A2(G20), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT23), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n495), .A2(KEYINPUT82), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(KEYINPUT82), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g0298(.A1(new_n497), .A2(new_n494), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n493), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n278), .A2(new_n207), .A3(G87), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT22), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n492), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n505), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n507), .A2(new_n501), .A3(KEYINPUT24), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n268), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n486), .A2(new_n221), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n251), .A2(new_n221), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n512), .B(KEYINPUT25), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n509), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n278), .A2(G257), .A3(G1698), .ZN(new_n516));
  INV_X1    g0316(.A(G294), .ZN(new_n517));
  OAI221_X1 g0317(.A(new_n516), .B1(new_n260), .B2(new_n517), .C1(new_n417), .C2(new_n216), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n277), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n477), .A2(G264), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n476), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n331), .ZN(new_n522));
  INV_X1    g0322(.A(new_n521), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n408), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n515), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n251), .A2(new_n460), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n458), .A2(KEYINPUT74), .ZN(new_n527));
  AOI211_X1 g0327(.A(new_n452), .B(new_n271), .C1(new_n455), .C2(new_n457), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n488), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n479), .A2(new_n331), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n489), .A2(new_n408), .A3(new_n476), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n491), .A2(new_n525), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n502), .A2(new_n492), .A3(new_n505), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT24), .B1(new_n507), .B2(new_n501), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n271), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n536), .A2(new_n510), .A3(new_n513), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n523), .A2(G190), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n521), .A2(G200), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT79), .B1(new_n486), .B2(new_n427), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT79), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n484), .A2(new_n542), .A3(new_n426), .A4(new_n485), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT78), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n264), .A2(G97), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT77), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n460), .B1(new_n261), .B2(new_n263), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT77), .B1(new_n550), .B2(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n207), .B1(new_n318), .B2(new_n548), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n445), .A2(new_n215), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n321), .A2(new_n323), .A3(new_n207), .A4(G68), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n549), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n268), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n252), .A2(new_n426), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n545), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  AOI211_X1 g0361(.A(KEYINPUT78), .B(new_n559), .C1(new_n557), .C2(new_n268), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n544), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n278), .B1(G238), .B2(G1698), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n279), .A2(G244), .ZN(new_n565));
  INV_X1    g0365(.A(G116), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n564), .A2(new_n565), .B1(new_n260), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n277), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n298), .A2(new_n299), .B1(new_n216), .B2(new_n471), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(G274), .B2(new_n471), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n331), .ZN(new_n572));
  INV_X1    g0372(.A(new_n571), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n408), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n563), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(G200), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n568), .B2(new_n570), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n573), .B2(G190), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n487), .A2(G87), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n562), .C2(new_n561), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n540), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n278), .A2(G257), .A3(new_n279), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT80), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n278), .A2(KEYINPUT80), .A3(G257), .A4(new_n279), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G303), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n282), .A2(new_n222), .B1(new_n587), .B2(new_n278), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n277), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n477), .A2(G270), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n476), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G200), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT81), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n593), .A2(KEYINPUT20), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n566), .A2(G20), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n466), .B(new_n207), .C1(G33), .C2(new_n460), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n268), .A2(new_n594), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n593), .A3(KEYINPUT20), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n271), .B1(G20), .B2(new_n566), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(KEYINPUT20), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(new_n594), .A4(new_n596), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n251), .A2(new_n566), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n484), .A2(G116), .A3(new_n485), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n598), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n592), .B(new_n605), .C1(new_n395), .C2(new_n591), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n591), .A2(new_n604), .A3(G169), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n591), .A2(new_n408), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n604), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n591), .A2(new_n604), .A3(KEYINPUT21), .A4(G169), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n606), .A2(new_n609), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n442), .A2(new_n533), .A3(new_n581), .A4(new_n614), .ZN(G372));
  NAND2_X1  g0415(.A1(new_n313), .A2(new_n314), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT83), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n414), .B2(new_n412), .ZN(new_n620));
  INV_X1    g0420(.A(new_n411), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n413), .B1(new_n387), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n407), .A2(KEYINPUT18), .A3(new_n411), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(KEYINPUT83), .A3(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n431), .A2(KEYINPUT84), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n431), .A2(KEYINPUT84), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n357), .A2(new_n358), .A3(new_n355), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n629), .A2(new_n630), .B1(new_n352), .B2(new_n340), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n404), .B(KEYINPUT17), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n625), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n441), .B1(new_n618), .B2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n575), .A3(new_n580), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n636), .A2(new_n575), .A3(KEYINPUT26), .A4(new_n580), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n525), .A2(new_n611), .A3(new_n612), .A4(new_n609), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n491), .A2(new_n532), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n581), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n575), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n442), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n635), .A2(new_n646), .ZN(G369));
  OR2_X1    g0447(.A1(new_n613), .A2(KEYINPUT87), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n250), .A2(G20), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n206), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n604), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT86), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n613), .A2(KEYINPUT87), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n648), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n515), .A2(new_n522), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n515), .A2(new_n655), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n660), .A2(new_n524), .B1(new_n540), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n525), .A2(new_n655), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(new_n657), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n659), .A2(new_n664), .A3(G330), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT88), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n540), .A2(new_n661), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n525), .ZN(new_n670));
  INV_X1    g0470(.A(new_n655), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n663), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n210), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G1), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n445), .A2(new_n215), .A3(new_n566), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n678), .A2(new_n679), .B1(new_n231), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n591), .A2(new_n408), .A3(new_n571), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n489), .A3(new_n523), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT89), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n682), .A2(new_n489), .A3(new_n523), .A4(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n591), .A2(new_n479), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n408), .A3(new_n521), .A4(new_n571), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n686), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n655), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT31), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n581), .A2(new_n533), .A3(new_n614), .A4(new_n671), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n575), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n639), .B2(new_n640), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n655), .B1(new_n700), .B2(new_n644), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n698), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n681), .B1(new_n704), .B2(G1), .ZN(G364));
  NAND2_X1  g0505(.A1(new_n659), .A2(new_n666), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n697), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(KEYINPUT90), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n697), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n708), .B(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n678), .B1(G45), .B2(new_n649), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G13), .A2(G33), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n712), .B1(new_n706), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n229), .B1(G20), .B2(new_n331), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n207), .A2(G190), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n408), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n408), .A2(new_n576), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n719), .ZN(new_n723));
  OAI221_X1 g0523(.A(new_n278), .B1(new_n721), .B2(new_n284), .C1(new_n224), .C2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n207), .A2(new_n395), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n576), .A2(G179), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n215), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n722), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n720), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n729), .A2(new_n202), .B1(new_n730), .B2(new_n219), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G179), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n719), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G159), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n728), .B(new_n731), .C1(KEYINPUT32), .C2(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n395), .A2(G179), .A3(G200), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n207), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n736), .B1(KEYINPUT32), .B2(new_n735), .C1(new_n460), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n719), .A2(new_n726), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI211_X1 g0541(.A(new_n724), .B(new_n739), .C1(G107), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n729), .B(KEYINPUT94), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G326), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n734), .A2(G329), .ZN(new_n745));
  INV_X1    g0545(.A(new_n738), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n278), .B1(new_n746), .B2(G294), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G283), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n740), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G322), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n587), .A2(new_n727), .B1(new_n730), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g0552(.A(KEYINPUT33), .B(G317), .Z(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n723), .B1(new_n721), .B2(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n748), .A2(new_n750), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n718), .B1(new_n742), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n716), .A2(new_n718), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT93), .Z(new_n759));
  NAND3_X1  g0559(.A1(new_n210), .A2(G355), .A3(new_n278), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n244), .A2(G45), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT91), .Z(new_n762));
  NOR2_X1   g0562(.A1(new_n675), .A2(new_n278), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G45), .B2(new_n231), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n760), .B1(G116), .B2(new_n210), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT92), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n717), .B(new_n757), .C1(new_n759), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n713), .A2(new_n767), .ZN(G396));
  NAND2_X1  g0568(.A1(new_n645), .A2(new_n671), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n429), .A2(new_n671), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n626), .B2(new_n627), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n437), .B2(new_n770), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n645), .A2(new_n671), .A3(new_n772), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT96), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n693), .A2(new_n695), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G330), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n698), .A2(KEYINPUT96), .B1(new_n774), .B2(new_n775), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n698), .A2(KEYINPUT96), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n712), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n749), .A2(new_n723), .B1(new_n730), .B2(new_n517), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n738), .A2(new_n460), .B1(new_n729), .B2(new_n587), .ZN(new_n785));
  INV_X1    g0585(.A(new_n721), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n784), .B(new_n785), .C1(G116), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n734), .A2(G311), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n324), .B1(new_n727), .B2(new_n221), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT95), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n741), .A2(G87), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n787), .A2(new_n788), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n730), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G143), .A2(new_n793), .B1(new_n786), .B2(G159), .ZN(new_n794));
  INV_X1    g0594(.A(new_n729), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G137), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n794), .B(new_n796), .C1(new_n255), .C2(new_n723), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT34), .Z(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G132), .B2(new_n734), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n741), .A2(G68), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(new_n219), .C2(new_n738), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n278), .B1(new_n727), .B2(new_n202), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n792), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n718), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n718), .A2(new_n714), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n284), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n804), .B(new_n806), .C1(new_n772), .C2(new_n715), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n783), .B1(new_n712), .B2(new_n807), .ZN(G384));
  AOI21_X1  g0608(.A(new_n566), .B1(new_n456), .B2(KEYINPUT35), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n809), .B(new_n230), .C1(KEYINPUT35), .C2(new_n456), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT36), .ZN(new_n811));
  OAI21_X1  g0611(.A(G77), .B1(new_n219), .B2(new_n224), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n812), .A2(new_n231), .B1(G50), .B2(new_n224), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n813), .A2(G1), .A3(new_n250), .ZN(new_n814));
  INV_X1    g0614(.A(new_n653), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n625), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n431), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n671), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n775), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n352), .A2(new_n655), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n360), .B2(new_n353), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n630), .A2(new_n821), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(new_n340), .B2(new_n352), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n822), .A2(KEYINPUT97), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT97), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT70), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n630), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n354), .A2(KEYINPUT70), .A3(new_n355), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n352), .B(new_n655), .C1(new_n830), .C2(new_n340), .ZN(new_n831));
  INV_X1    g0631(.A(new_n824), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n826), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n825), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n820), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n382), .A2(KEYINPUT16), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n363), .B1(new_n836), .B2(new_n383), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n415), .A2(new_n815), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n411), .A2(new_n815), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n404), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT37), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n407), .B1(new_n411), .B2(new_n815), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n404), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n839), .A2(KEYINPUT38), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT38), .B1(new_n839), .B2(new_n846), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n817), .B1(new_n835), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n353), .A2(new_n655), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT39), .B1(new_n847), .B2(new_n848), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT39), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n839), .A2(KEYINPUT38), .A3(new_n846), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n843), .A2(new_n844), .A3(new_n404), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n844), .B1(new_n843), .B2(new_n404), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n620), .A2(new_n624), .A3(new_n632), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n387), .A2(new_n653), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n854), .B(new_n855), .C1(new_n861), .C2(KEYINPUT38), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n852), .B1(new_n853), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT98), .B1(new_n850), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n862), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n839), .A2(new_n846), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n854), .B1(new_n868), .B2(new_n855), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n851), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT97), .B1(new_n822), .B2(new_n824), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n831), .A2(new_n826), .A3(new_n832), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n775), .B2(new_n819), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n868), .A2(new_n855), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n816), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT98), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n870), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n864), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n703), .A2(new_n442), .A3(new_n702), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n635), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n879), .B(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n871), .A2(new_n772), .A3(new_n872), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(new_n696), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT40), .B1(new_n884), .B2(new_n875), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n834), .A2(new_n778), .A3(KEYINPUT40), .A4(new_n772), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n859), .A2(new_n860), .ZN(new_n888));
  INV_X1    g0688(.A(new_n858), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n847), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT99), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n887), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n883), .A2(new_n894), .A3(new_n696), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n855), .B1(new_n861), .B2(KEYINPUT38), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT99), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(G330), .B(new_n886), .C1(new_n893), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n698), .A2(new_n442), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n892), .B1(new_n887), .B2(new_n891), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n895), .A2(KEYINPUT99), .A3(new_n896), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n885), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n442), .A3(new_n778), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n882), .A2(new_n905), .B1(new_n206), .B2(new_n649), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT100), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n882), .A2(new_n905), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n811), .B(new_n814), .C1(new_n907), .C2(new_n908), .ZN(G367));
  INV_X1    g0709(.A(KEYINPUT88), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n667), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n529), .A2(new_n655), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n491), .A2(new_n532), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n532), .B2(new_n671), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n643), .A2(new_n642), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT42), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n664), .A2(new_n917), .A3(new_n918), .A4(new_n672), .ZN(new_n919));
  INV_X1    g0719(.A(new_n663), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n670), .A2(new_n920), .A3(new_n672), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT42), .B1(new_n921), .B2(new_n916), .ZN(new_n922));
  INV_X1    g0722(.A(new_n491), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n532), .B1(new_n923), .B2(new_n525), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n671), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n919), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT43), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n579), .B1(new_n561), .B2(new_n562), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n655), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n575), .A2(new_n580), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n575), .A2(new_n929), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n926), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n932), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n926), .A2(KEYINPUT43), .A3(new_n934), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n915), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT101), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT101), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n915), .B(new_n940), .C1(new_n936), .C2(new_n937), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OR3_X1    g0742(.A1(new_n915), .A2(new_n936), .A3(new_n937), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n676), .B(KEYINPUT41), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT44), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n673), .B2(new_n914), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n665), .A2(new_n671), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n920), .B1(new_n662), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n914), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(KEYINPUT44), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n951), .A3(KEYINPUT102), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT45), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n949), .B2(new_n950), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n914), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT102), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n957), .B(new_n946), .C1(new_n673), .C2(new_n914), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n952), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT103), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n668), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n911), .A2(KEYINPUT103), .A3(new_n959), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n670), .A2(new_n920), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n948), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n921), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT104), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT104), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n964), .A2(new_n967), .A3(new_n921), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n966), .B(new_n968), .C1(new_n697), .C2(new_n706), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n707), .A2(KEYINPUT104), .A3(new_n965), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n961), .A2(new_n704), .A3(new_n962), .A4(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n945), .B1(new_n972), .B2(new_n704), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n206), .B1(new_n649), .B2(G45), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n942), .B(new_n943), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n759), .B1(new_n240), .B2(new_n763), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n675), .A2(new_n426), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n712), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n746), .A2(G107), .ZN(new_n980));
  INV_X1    g0780(.A(new_n727), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(KEYINPUT46), .A3(G116), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT46), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n727), .B2(new_n566), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n980), .A2(new_n982), .A3(new_n324), .A4(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n723), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G294), .A2(new_n986), .B1(new_n786), .B2(G283), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G303), .A2(new_n793), .B1(new_n734), .B2(G317), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n460), .C2(new_n740), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n985), .B(new_n989), .C1(G311), .C2(new_n743), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n734), .A2(G137), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n324), .B1(new_n743), .B2(G143), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n284), .B2(new_n740), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n219), .A2(new_n727), .B1(new_n730), .B2(new_n255), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n746), .A2(G68), .ZN(new_n995));
  INV_X1    g0795(.A(G159), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(new_n202), .B2(new_n721), .C1(new_n996), .C2(new_n723), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n993), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n990), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT47), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n718), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n979), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT105), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n716), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n934), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n976), .A2(new_n1005), .ZN(G387));
  AOI22_X1  g0806(.A1(G311), .A2(new_n986), .B1(new_n793), .B2(G317), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n587), .B2(new_n721), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G322), .B2(new_n743), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT48), .Z(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n749), .B2(new_n738), .C1(new_n517), .C2(new_n727), .ZN(new_n1011));
  XOR2_X1   g0811(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G116), .A2(new_n741), .B1(new_n734), .B2(G326), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n324), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n730), .A2(new_n202), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G77), .A2(new_n981), .B1(new_n734), .B2(G150), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1018), .A2(KEYINPUT107), .B1(G97), .B2(new_n741), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n729), .A2(new_n996), .B1(new_n721), .B2(new_n224), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n324), .B(new_n1020), .C1(new_n258), .C2(new_n986), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT107), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n1017), .A2(new_n1022), .B1(new_n426), .B2(new_n746), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1015), .B1(new_n1016), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n718), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n759), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n763), .B1(new_n237), .B2(new_n288), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n210), .A2(new_n278), .A3(new_n679), .ZN(new_n1029));
  AOI211_X1 g0829(.A(G45), .B(new_n679), .C1(G68), .C2(G77), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n258), .A2(new_n202), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT50), .Z(new_n1032));
  AOI22_X1  g0832(.A1(new_n1028), .A2(new_n1029), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n210), .A2(G107), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1027), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n963), .A2(new_n716), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1026), .A2(new_n711), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n974), .B1(new_n969), .B2(new_n970), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT106), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n704), .A2(new_n971), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT109), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n704), .A2(new_n971), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n676), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1037), .B(new_n1039), .C1(new_n1044), .C2(new_n1045), .ZN(G393));
  OR2_X1    g0846(.A1(new_n911), .A2(new_n959), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n911), .A2(new_n959), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(new_n974), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n950), .A2(new_n716), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G303), .A2(new_n986), .B1(new_n786), .B2(G294), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n566), .B2(new_n738), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT111), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n740), .A2(new_n221), .B1(new_n733), .B2(new_n751), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n278), .B(new_n1055), .C1(G283), .C2(new_n981), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G317), .A2(new_n795), .B1(new_n793), .B2(G311), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  NAND3_X1  g0858(.A1(new_n1054), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n324), .B1(new_n734), .B2(G143), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1060), .B(new_n791), .C1(new_n224), .C2(new_n727), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT110), .Z(new_n1062));
  AOI22_X1  g0862(.A1(new_n986), .A2(G50), .B1(new_n786), .B2(new_n258), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n284), .C2(new_n738), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n729), .A2(new_n255), .B1(new_n730), .B2(new_n996), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT51), .Z(new_n1066));
  OAI21_X1  g0866(.A(new_n1059), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n718), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n763), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1027), .B1(new_n460), .B2(new_n210), .C1(new_n247), .C2(new_n1069), .ZN(new_n1070));
  AND4_X1   g0870(.A1(new_n711), .A2(new_n1051), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1050), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1049), .A2(new_n1043), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n676), .A3(new_n972), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(G390));
  AOI22_X1  g0875(.A1(new_n701), .A2(new_n772), .B1(new_n818), .B2(new_n671), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n873), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n696), .A2(new_n773), .A3(new_n697), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(new_n835), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n880), .A2(new_n635), .A3(new_n899), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1078), .B1(new_n1077), .B2(new_n835), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n896), .B(new_n852), .C1(new_n1076), .C2(new_n873), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n853), .A2(new_n862), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n851), .B1(new_n820), .B2(new_n834), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1078), .A2(new_n834), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(KEYINPUT112), .A3(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n853), .B(new_n862), .C1(new_n874), .C2(new_n851), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(KEYINPUT112), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT112), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1078), .A2(new_n1093), .A3(new_n834), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .A4(new_n1085), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1084), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1083), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n676), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n853), .A2(new_n714), .A3(new_n862), .ZN(new_n1100));
  OR3_X1    g0900(.A1(new_n727), .A2(KEYINPUT53), .A3(new_n255), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n324), .B1(new_n734), .B2(G125), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT54), .B(G143), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n786), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(KEYINPUT53), .B1(new_n727), .B2(new_n255), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n746), .A2(G159), .B1(new_n795), .B2(G128), .ZN(new_n1107));
  INV_X1    g0907(.A(G132), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1107), .B1(new_n202), .B2(new_n740), .C1(new_n1108), .C2(new_n730), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(G137), .C2(new_n986), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n746), .A2(G77), .B1(G294), .B2(new_n734), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1111), .B(new_n800), .C1(new_n749), .C2(new_n729), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n728), .B1(G107), .B2(new_n986), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n324), .C1(new_n460), .C2(new_n721), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1112), .B(new_n1114), .C1(G116), .C2(new_n793), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n718), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n805), .A2(new_n259), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1100), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1097), .A2(new_n975), .B1(new_n711), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1099), .A2(new_n1119), .ZN(G378));
  XNOR2_X1  g0920(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n273), .A2(new_n815), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT55), .Z(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n618), .B2(new_n440), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n616), .A2(new_n617), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT85), .B1(new_n313), .B2(new_n314), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n440), .B(new_n1125), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1122), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n440), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1124), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(new_n1121), .A3(new_n1129), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n898), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n903), .A2(G330), .A3(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1136), .A2(new_n879), .A3(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1136), .A2(new_n1138), .B1(new_n878), .B2(new_n864), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n975), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n714), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n324), .A2(new_n287), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n746), .A2(G68), .B1(new_n793), .B2(G107), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n219), .B2(new_n740), .C1(new_n749), .C2(new_n733), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G97), .B2(new_n986), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n566), .B2(new_n729), .C1(new_n427), .C2(new_n721), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1143), .B(new_n1147), .C1(G77), .C2(new_n981), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT58), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n746), .A2(G150), .B1(new_n795), .B2(G125), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(G132), .A2(new_n986), .B1(new_n786), .B2(G137), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n981), .A2(new_n1103), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n793), .A2(G128), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT59), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(G33), .A2(G41), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT113), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT115), .B(G124), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1158), .B1(new_n996), .B2(new_n740), .C1(new_n733), .C2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1157), .A2(new_n1143), .A3(new_n202), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(KEYINPUT114), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(KEYINPUT114), .B2(new_n1162), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n718), .B1(new_n1149), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n805), .A2(new_n202), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1142), .A2(new_n711), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1141), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1081), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1098), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n677), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1081), .B1(new_n1097), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n864), .A2(new_n878), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n898), .A2(new_n1135), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1137), .B1(new_n903), .B2(G330), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1136), .A2(new_n879), .A3(new_n1138), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1175), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT57), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1168), .B1(new_n1173), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT117), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n974), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1167), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n676), .B1(new_n1181), .B2(KEYINPUT57), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1172), .B(new_n1175), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT117), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1184), .A2(new_n1192), .ZN(G375));
  INV_X1    g0993(.A(new_n1082), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1079), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1081), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1084), .A2(new_n1196), .A3(new_n944), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n834), .A2(new_n715), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n729), .A2(new_n1108), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n324), .B1(new_n986), .B2(new_n1103), .ZN(new_n1200));
  INV_X1    g1000(.A(G128), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1200), .B1(new_n1201), .B2(new_n733), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1199), .B(new_n1202), .C1(G150), .C2(new_n786), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n793), .A2(G137), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n746), .A2(G50), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G159), .A2(new_n981), .B1(new_n741), .B2(G58), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n723), .A2(new_n566), .B1(new_n740), .B2(new_n284), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n278), .B(new_n1208), .C1(G303), .C2(new_n734), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n981), .A2(G97), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n793), .A2(G283), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n427), .A2(new_n738), .B1(new_n517), .B2(new_n729), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G107), .B2(new_n786), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1001), .B1(new_n1207), .B2(new_n1214), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n718), .A2(G68), .A3(new_n714), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1198), .A2(new_n712), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1174), .B2(new_n975), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1197), .A2(new_n1218), .ZN(G381));
  INV_X1    g1019(.A(G378), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1184), .A2(new_n1192), .A3(new_n1220), .ZN(new_n1221));
  OR3_X1    g1021(.A1(new_n1221), .A2(G384), .A3(G381), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n976), .A2(new_n1005), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n704), .A2(new_n971), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n677), .B1(new_n1224), .B2(KEYINPUT109), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n1043), .A3(new_n1042), .ZN(new_n1226));
  INV_X1    g1026(.A(G396), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1223), .A2(new_n1228), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1222), .A2(new_n1229), .ZN(G407));
  OAI221_X1 g1030(.A(G213), .B1(G343), .B2(new_n1221), .C1(new_n1222), .C2(new_n1229), .ZN(G409));
  NAND2_X1  g1031(.A1(G387), .A2(G390), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT122), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1223), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(G393), .A2(G396), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1235), .A2(new_n1228), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1223), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT123), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1235), .A2(new_n1228), .B1(KEYINPUT123), .B2(G390), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1241), .A2(new_n1232), .A3(new_n1233), .A4(new_n1223), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1237), .A2(new_n1239), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT124), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1234), .A2(new_n1236), .B1(new_n1238), .B2(KEYINPUT123), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1246), .A2(KEYINPUT124), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT63), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n944), .B(new_n1170), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT118), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1181), .A2(KEYINPUT118), .A3(new_n944), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1220), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT119), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1141), .A2(KEYINPUT119), .A3(new_n1167), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1254), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1190), .A2(G378), .ZN(new_n1260));
  INV_X1    g1060(.A(G213), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(G343), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1084), .B(new_n676), .C1(new_n1196), .C2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT60), .B1(new_n1195), .B2(new_n1081), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1218), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  XOR2_X1   g1067(.A(G384), .B(KEYINPUT120), .Z(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(G384), .A2(KEYINPUT120), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1218), .B(new_n1270), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1259), .A2(new_n1260), .A3(new_n1263), .A4(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1248), .B1(new_n1249), .B2(new_n1273), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1262), .A2(G2897), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1272), .B(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1263), .B1(new_n1183), .B2(new_n1220), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1252), .A2(new_n1253), .A3(new_n1220), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(KEYINPUT121), .B(new_n1276), .C1(new_n1277), .C2(new_n1280), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1273), .A2(new_n1249), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1276), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT121), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1274), .A2(new_n1281), .A3(new_n1282), .A4(new_n1285), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1273), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT62), .B1(new_n1273), .B2(KEYINPUT126), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1283), .A2(new_n1289), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1246), .A2(new_n1242), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1286), .B1(new_n1291), .B2(new_n1293), .ZN(G405));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1272), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1221), .B2(new_n1260), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1221), .A2(new_n1260), .A3(new_n1296), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1298), .A2(new_n1293), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1293), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(G402));
endmodule


