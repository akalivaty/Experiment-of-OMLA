//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT35), .ZN(new_n203));
  INV_X1    g002(.A(G204gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G197gat), .ZN(new_n205));
  INV_X1    g004(.A(G197gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT69), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n208), .B1(new_n205), .B2(new_n207), .ZN(new_n210));
  NAND2_X1  g009(.A1(G211gat), .A2(G218gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT22), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT70), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n211), .A2(KEYINPUT70), .A3(new_n212), .ZN(new_n214));
  OAI22_X1  g013(.A1(new_n209), .A2(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G211gat), .B(G218gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OAI221_X1 g017(.A(new_n216), .B1(new_n214), .B2(new_n213), .C1(new_n209), .C2(new_n210), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n222), .A2(new_n223), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G183gat), .ZN(new_n231));
  INV_X1    g030(.A(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(KEYINPUT24), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n224), .A2(new_n230), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n224), .A2(new_n230), .A3(new_n235), .A4(KEYINPUT25), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT27), .B(G183gat), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n240), .B(new_n232), .C1(KEYINPUT64), .C2(KEYINPUT28), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n231), .A2(KEYINPUT27), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT27), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G183gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n244), .A3(new_n232), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n226), .A2(new_n227), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n234), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n251), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n238), .A2(new_n239), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT73), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n239), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n248), .A2(new_n253), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT73), .ZN(new_n260));
  INV_X1    g059(.A(new_n255), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n254), .A2(KEYINPUT72), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT29), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n221), .B(new_n263), .C1(new_n267), .C2(new_n261), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n269), .B(new_n255), .C1(new_n254), .C2(KEYINPUT29), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n255), .B1(new_n265), .B2(new_n266), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT29), .B1(new_n257), .B2(new_n258), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT71), .B1(new_n272), .B2(new_n261), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n220), .B(new_n270), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G8gat), .B(G36gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(G64gat), .B(G92gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n268), .A2(new_n274), .A3(new_n278), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(KEYINPUT30), .A3(new_n281), .ZN(new_n282));
  OR3_X1    g081(.A1(new_n275), .A2(KEYINPUT30), .A3(new_n279), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT78), .ZN(new_n285));
  AND2_X1   g084(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n287));
  OAI21_X1  g086(.A(G155gat), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT2), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n290));
  INV_X1    g089(.A(G148gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(new_n291), .B2(G141gat), .ZN(new_n292));
  INV_X1    g091(.A(G141gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n292), .B(new_n294), .C1(new_n293), .C2(G148gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n296));
  INV_X1    g095(.A(G155gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(G162gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G155gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n296), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G155gat), .B(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT75), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n289), .A2(new_n295), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G141gat), .B(G148gat), .ZN(new_n305));
  OAI22_X1  g104(.A1(new_n305), .A2(KEYINPUT2), .B1(new_n298), .B2(new_n300), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT3), .ZN(new_n309));
  XOR2_X1   g108(.A(G113gat), .B(G120gat), .Z(new_n310));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311));
  XNOR2_X1  g110(.A(G127gat), .B(G134gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n311), .ZN(new_n314));
  OR2_X1    g113(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n315), .A2(KEYINPUT66), .A3(G127gat), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n319));
  INV_X1    g118(.A(G134gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(G127gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(new_n316), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n323), .B2(G127gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n313), .B1(new_n318), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n304), .A2(new_n326), .A3(new_n306), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n308), .B1(new_n307), .B2(KEYINPUT3), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n285), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n329), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n327), .A2(new_n325), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT78), .A4(new_n309), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G127gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n322), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n314), .B(new_n317), .C1(new_n336), .C2(new_n321), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n337), .A2(new_n306), .A3(new_n304), .A4(new_n313), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n307), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n337), .A2(new_n313), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n304), .A2(KEYINPUT79), .A3(new_n306), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n340), .B1(new_n345), .B2(new_n339), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(KEYINPUT5), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n334), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT0), .ZN(new_n353));
  XNOR2_X1  g152(.A(G57gat), .B(G85gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n348), .B1(new_n338), .B2(new_n339), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(new_n345), .B2(new_n339), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n334), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n325), .A2(new_n307), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n338), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n348), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT5), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n356), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n358), .B1(new_n330), .B2(new_n333), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n367), .A2(KEYINPUT80), .A3(new_n364), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n351), .B(new_n355), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n360), .A2(new_n356), .A3(new_n365), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT80), .B1(new_n367), .B2(new_n364), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n350), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(new_n355), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n351), .B1(new_n366), .B2(new_n368), .ZN(new_n377));
  INV_X1    g176(.A(new_n355), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(KEYINPUT6), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n284), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G228gat), .A2(G233gat), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n326), .B1(new_n220), .B2(KEYINPUT29), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(new_n307), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n327), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT81), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n327), .A2(new_n388), .A3(new_n385), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n220), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n218), .B2(new_n219), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n304), .A2(KEYINPUT79), .A3(new_n306), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT79), .B1(new_n304), .B2(new_n306), .ZN(new_n393));
  OAI22_X1  g192(.A1(new_n391), .A2(KEYINPUT3), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n386), .A2(new_n220), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n384), .A2(new_n390), .B1(new_n396), .B2(new_n382), .ZN(new_n397));
  INV_X1    g196(.A(G22gat), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n390), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n396), .A2(new_n382), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT31), .B(G50gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n404), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n409), .ZN(new_n411));
  AOI211_X1 g210(.A(KEYINPUT83), .B(new_n411), .C1(new_n402), .C2(new_n405), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n403), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT82), .B1(new_n397), .B2(new_n398), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT83), .B1(new_n414), .B2(new_n411), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n406), .A2(new_n404), .A3(new_n409), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n415), .A2(new_n416), .A3(new_n402), .A4(new_n399), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT67), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n259), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n325), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n259), .A2(new_n343), .A3(new_n419), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT34), .ZN(new_n425));
  NAND2_X1  g224(.A1(G227gat), .A2(G233gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n425), .B1(new_n424), .B2(new_n426), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT68), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n429), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT68), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n427), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n422), .A2(G227gat), .A3(G233gat), .A4(new_n423), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435));
  XOR2_X1   g234(.A(G15gat), .B(G43gat), .Z(new_n436));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n434), .B(KEYINPUT32), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n434), .A2(KEYINPUT32), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n434), .A2(new_n435), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n438), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n430), .A2(new_n433), .A3(new_n440), .A4(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n441), .A2(new_n442), .A3(new_n438), .ZN(new_n446));
  INV_X1    g245(.A(new_n440), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n432), .B(new_n445), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n202), .A2(KEYINPUT35), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n418), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n203), .B1(new_n381), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n450), .ZN(new_n453));
  AOI221_X4 g252(.A(new_n453), .B1(new_n448), .B2(new_n444), .C1(new_n413), .C2(new_n417), .ZN(new_n454));
  INV_X1    g253(.A(new_n284), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n377), .A2(new_n378), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n370), .A3(new_n369), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n457), .B2(new_n379), .ZN(new_n458));
  INV_X1    g257(.A(new_n203), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT38), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n279), .A2(KEYINPUT37), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n280), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n275), .A2(KEYINPUT37), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n279), .B1(new_n275), .B2(KEYINPUT37), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n221), .B(new_n270), .C1(new_n271), .C2(new_n273), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n220), .B(new_n263), .C1(new_n267), .C2(new_n261), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT37), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n461), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n281), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n472), .A3(new_n379), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n361), .A2(new_n347), .A3(new_n338), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT39), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT85), .ZN(new_n478));
  INV_X1    g277(.A(new_n340), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n392), .A2(new_n393), .A3(new_n325), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(KEYINPUT4), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n330), .B2(new_n333), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n478), .B1(new_n482), .B2(new_n347), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n334), .A2(new_n346), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT84), .B(KEYINPUT39), .Z(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n348), .A3(new_n485), .ZN(new_n486));
  AND4_X1   g285(.A1(new_n475), .A2(new_n483), .A3(new_n486), .A4(new_n355), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT86), .B(KEYINPUT40), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n347), .B1(new_n334), .B2(new_n346), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n378), .B1(new_n490), .B2(new_n485), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n489), .B1(new_n491), .B2(new_n483), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n283), .B(new_n282), .C1(new_n374), .C2(new_n355), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n474), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n483), .A2(new_n486), .A3(new_n355), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n488), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n491), .A2(new_n475), .A3(new_n483), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n499), .A2(new_n455), .A3(KEYINPUT87), .A4(new_n456), .ZN(new_n500));
  AND4_X1   g299(.A1(new_n473), .A2(new_n495), .A3(new_n500), .A4(new_n418), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n448), .A2(KEYINPUT36), .A3(new_n444), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT36), .B1(new_n444), .B2(new_n448), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n458), .B2(new_n418), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n452), .B(new_n460), .C1(new_n501), .C2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT14), .B(G29gat), .ZN(new_n507));
  INV_X1    g306(.A(G36gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G29gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT90), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n512), .A2(new_n514), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n512), .A2(new_n515), .A3(new_n519), .A4(new_n514), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n522), .A2(G1gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT91), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT16), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n522), .B1(new_n525), .B2(G1gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n527), .A3(G8gat), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n523), .B(new_n526), .C1(KEYINPUT91), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT93), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n521), .A2(KEYINPUT93), .A3(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n521), .A2(new_n531), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT13), .Z(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(KEYINPUT94), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n537), .B1(new_n534), .B2(new_n535), .ZN(new_n544));
  INV_X1    g343(.A(new_n541), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT18), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n521), .B(KEYINPUT17), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n531), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n536), .ZN(new_n553));
  INV_X1    g352(.A(new_n540), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n549), .A2(new_n551), .B1(new_n534), .B2(new_n535), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(KEYINPUT18), .A3(new_n540), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n547), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G113gat), .B(G141gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT89), .B(G197gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT11), .B(G169gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT12), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n558), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n547), .A2(new_n555), .A3(new_n557), .A4(new_n564), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n506), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT41), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n570), .B(new_n573), .Z(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OAI22_X1  g376(.A1(new_n577), .A2(KEYINPUT105), .B1(new_n572), .B2(new_n571), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT100), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT7), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n581), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n579), .B2(new_n580), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT102), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(KEYINPUT102), .A3(new_n589), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n584), .A2(new_n588), .A3(new_n586), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n584), .A2(KEYINPUT101), .A3(new_n588), .A4(new_n586), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n592), .A2(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n597), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT102), .B1(new_n587), .B2(new_n589), .ZN(new_n602));
  AOI211_X1 g401(.A(new_n591), .B(new_n588), .C1(new_n584), .C2(new_n586), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT103), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n578), .B1(new_n606), .B2(new_n521), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n600), .A2(new_n605), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT104), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n609), .A3(new_n549), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n609), .B1(new_n608), .B2(new_n549), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n607), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n577), .A2(KEYINPUT105), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n612), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n610), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n614), .B1(new_n618), .B2(new_n607), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n575), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n613), .A2(new_n615), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n614), .A3(new_n607), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(new_n622), .A3(new_n574), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(G183gat), .B(G211gat), .Z(new_n625));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626));
  NOR2_X1   g425(.A1(G71gat), .A2(G78gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G57gat), .B(G64gat), .Z(new_n631));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT9), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n631), .A2(new_n632), .B1(new_n633), .B2(new_n628), .ZN(new_n634));
  XNOR2_X1  g433(.A(G57gat), .B(G64gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT96), .ZN(new_n636));
  AOI211_X1 g435(.A(new_n627), .B(new_n630), .C1(new_n634), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n627), .A2(KEYINPUT9), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n635), .B1(new_n628), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n626), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n634), .A2(new_n636), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n630), .A2(new_n627), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT97), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n645), .A2(KEYINPUT21), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n645), .B2(KEYINPUT21), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n335), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n335), .B1(new_n647), .B2(new_n648), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n625), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n651), .ZN(new_n653));
  INV_X1    g452(.A(new_n625), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n654), .A3(new_n649), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT98), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G155gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n645), .A2(KEYINPUT21), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n530), .A3(new_n528), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT99), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n661), .A2(KEYINPUT99), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  INV_X1    g465(.A(new_n659), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n656), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n652), .A2(new_n655), .A3(new_n668), .A4(new_n665), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT10), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n640), .B2(new_n644), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n600), .A2(new_n605), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n601), .A2(new_n643), .A3(new_n590), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n676), .B(new_n673), .C1(new_n645), .C2(new_n598), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G230gat), .A2(G233gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n676), .B1(new_n645), .B2(new_n598), .ZN(new_n681));
  INV_X1    g480(.A(new_n679), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(G120gat), .B(G148gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(G176gat), .B(G204gat), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n684), .B(new_n685), .Z(new_n686));
  NAND3_X1  g485(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n686), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n682), .B1(new_n675), .B2(new_n677), .ZN(new_n689));
  INV_X1    g488(.A(new_n683), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n624), .A2(new_n672), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT106), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n569), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n376), .A2(new_n380), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G1gat), .ZN(G1324gat));
  AND3_X1   g498(.A1(new_n569), .A2(new_n455), .A3(new_n695), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT16), .B(G8gat), .Z(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n529), .B2(new_n700), .ZN(new_n703));
  MUX2_X1   g502(.A(new_n702), .B(new_n703), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g503(.A(G15gat), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n696), .A2(new_n705), .A3(new_n449), .ZN(new_n706));
  INV_X1    g505(.A(new_n504), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n696), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n708), .B2(new_n705), .ZN(G1326gat));
  INV_X1    g508(.A(new_n418), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n696), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  INV_X1    g512(.A(new_n672), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n693), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n624), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n569), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n510), .A3(new_n697), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n620), .A2(new_n623), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n506), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n506), .A2(KEYINPUT44), .A3(new_n721), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n568), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n715), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n697), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n720), .A2(new_n731), .ZN(G1328gat));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n508), .A3(new_n455), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT46), .Z(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n729), .B2(new_n284), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1329gat));
  NAND4_X1  g535(.A1(new_n724), .A2(new_n707), .A3(new_n725), .A4(new_n728), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G43gat), .ZN(new_n738));
  INV_X1    g537(.A(G43gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n717), .A2(new_n739), .A3(new_n449), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n741), .A2(KEYINPUT108), .A3(KEYINPUT47), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT47), .B1(new_n741), .B2(KEYINPUT108), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(G1330gat));
  NAND3_X1  g543(.A1(new_n726), .A2(new_n710), .A3(new_n728), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n418), .A2(G50gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n569), .A2(new_n716), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(KEYINPUT48), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(KEYINPUT110), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(G50gat), .B2(new_n745), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(G1331gat));
  NOR4_X1   g552(.A1(new_n721), .A2(new_n714), .A3(new_n568), .A4(new_n693), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n506), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n697), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g556(.A(new_n284), .B(KEYINPUT111), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT112), .Z(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1333gat));
  NAND2_X1  g562(.A1(new_n755), .A2(new_n449), .ZN(new_n764));
  AOI21_X1  g563(.A(G71gat), .B1(new_n764), .B2(KEYINPUT113), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(KEYINPUT113), .B2(new_n764), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n755), .A2(G71gat), .A3(new_n707), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT50), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n766), .A2(new_n770), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1334gat));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n710), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g573(.A1(new_n672), .A2(new_n568), .A3(new_n693), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n726), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n730), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n501), .A2(new_n505), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n452), .A2(new_n460), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n778), .B(new_n721), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n672), .A2(new_n568), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n778), .B1(new_n506), .B2(new_n721), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT51), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n692), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n722), .A2(KEYINPUT114), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n787), .A2(new_n788), .A3(new_n782), .A4(new_n781), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n697), .A2(new_n579), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n777), .B1(new_n790), .B2(new_n791), .ZN(G1336gat));
  OAI21_X1  g591(.A(G92gat), .B1(new_n776), .B2(new_n758), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n758), .A2(G92gat), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n785), .A2(new_n789), .A3(new_n692), .A4(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n724), .A2(new_n455), .A3(new_n725), .A4(new_n775), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G92gat), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n797), .B1(new_n794), .B2(new_n800), .ZN(G1337gat));
  INV_X1    g600(.A(G99gat), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n776), .A2(new_n802), .A3(new_n504), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n449), .A3(new_n789), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n802), .ZN(G1338gat));
  NOR2_X1   g604(.A1(new_n418), .A2(G106gat), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n785), .A2(new_n789), .A3(new_n692), .A4(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n724), .A2(new_n710), .A3(new_n725), .A4(new_n775), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT53), .B1(new_n809), .B2(KEYINPUT115), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n807), .B(new_n809), .C1(KEYINPUT115), .C2(KEYINPUT53), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(G1339gat));
  NAND3_X1  g613(.A1(new_n675), .A2(new_n677), .A3(new_n682), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n680), .A2(KEYINPUT54), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n686), .B1(new_n689), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n687), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT116), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n822), .A3(new_n687), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT55), .B1(new_n816), .B2(new_n818), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n821), .A2(new_n568), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n556), .A2(new_n540), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n539), .A2(new_n541), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n563), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n567), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n692), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n721), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n824), .B1(new_n820), .B2(KEYINPUT116), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n823), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n620), .A2(new_n830), .A3(new_n623), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n714), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n694), .A2(new_n568), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n730), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n449), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n710), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n758), .ZN(new_n844));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n568), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n710), .B1(new_n837), .B2(new_n839), .ZN(new_n846));
  AND4_X1   g645(.A1(new_n697), .A2(new_n846), .A3(new_n449), .A4(new_n758), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n568), .A2(G113gat), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(G1340gat));
  INV_X1    g648(.A(G120gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n844), .A2(new_n850), .A3(new_n692), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n692), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(G120gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT117), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n851), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(G1341gat));
  NAND3_X1  g657(.A1(new_n844), .A2(new_n335), .A3(new_n672), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n847), .A2(new_n672), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n335), .B2(new_n860), .ZN(G1342gat));
  NAND2_X1  g660(.A1(new_n721), .A2(new_n284), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n322), .B(new_n862), .C1(new_n863), .C2(KEYINPUT56), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n843), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n847), .A2(new_n721), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(G134gat), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(G1343gat));
  NOR2_X1   g671(.A1(new_n707), .A2(new_n418), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT121), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n727), .A2(G141gat), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n840), .A2(new_n758), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(KEYINPUT122), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n758), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n730), .A2(new_n707), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n418), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n557), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT18), .B1(new_n556), .B2(new_n540), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n564), .B1(new_n886), .B2(new_n547), .ZN(new_n887));
  INV_X1    g686(.A(new_n567), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n825), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n831), .B1(new_n889), .B2(new_n820), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n624), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n721), .A2(new_n830), .A3(new_n823), .A4(new_n833), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n672), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n838), .B1(new_n893), .B2(KEYINPUT120), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n824), .B1(new_n566), .B2(new_n567), .ZN(new_n895));
  INV_X1    g694(.A(new_n820), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n895), .A2(new_n896), .B1(new_n692), .B2(new_n830), .ZN(new_n897));
  OAI22_X1  g696(.A1(new_n897), .A2(new_n721), .B1(new_n834), .B2(new_n835), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n714), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n883), .B1(new_n894), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n837), .A2(new_n839), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT57), .B1(new_n903), .B2(new_n710), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n568), .B(new_n880), .C1(new_n902), .C2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n878), .B1(new_n905), .B2(G141gat), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n877), .A2(KEYINPUT122), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n906), .B(new_n907), .ZN(G1344gat));
  NAND2_X1  g707(.A1(new_n880), .A2(new_n692), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n672), .B1(new_n898), .B2(KEYINPUT124), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n891), .A2(new_n911), .A3(new_n892), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n910), .A2(new_n912), .B1(new_n695), .B2(new_n727), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n881), .B1(new_n913), .B2(new_n418), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n903), .A2(new_n882), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n909), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT59), .B1(new_n916), .B2(new_n291), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n692), .B(new_n880), .C1(new_n902), .C2(new_n904), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n291), .A2(KEYINPUT59), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n840), .A2(new_n874), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n879), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n291), .A3(new_n692), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n923), .A2(new_n926), .ZN(G1345gat));
  OAI21_X1  g726(.A(new_n880), .B1(new_n902), .B2(new_n904), .ZN(new_n928));
  OAI21_X1  g727(.A(G155gat), .B1(new_n928), .B2(new_n714), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n297), .A3(new_n672), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1346gat));
  OR2_X1    g730(.A1(new_n286), .A2(new_n287), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(new_n928), .B2(new_n624), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n862), .A2(new_n932), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n924), .B2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n697), .A2(new_n284), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n449), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT125), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n846), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n846), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(new_n226), .A3(new_n727), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n697), .B1(new_n837), .B2(new_n839), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(new_n842), .A3(new_n879), .ZN(new_n946));
  AOI21_X1  g745(.A(G169gat), .B1(new_n946), .B2(new_n568), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n944), .A2(new_n947), .ZN(G1348gat));
  OAI21_X1  g747(.A(G176gat), .B1(new_n943), .B2(new_n693), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n227), .A3(new_n692), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1349gat));
  NAND3_X1  g750(.A1(new_n946), .A2(new_n240), .A3(new_n672), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n940), .A2(new_n672), .A3(new_n942), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n231), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT60), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT60), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n952), .B(new_n956), .C1(new_n953), .C2(new_n231), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n946), .A2(new_n232), .A3(new_n721), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n940), .A2(new_n721), .A3(new_n942), .ZN(new_n960));
  XNOR2_X1  g759(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n960), .A2(G190gat), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n960), .B2(G190gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1351gat));
  AND4_X1   g763(.A1(new_n730), .A2(new_n903), .A3(new_n879), .A4(new_n873), .ZN(new_n965));
  AOI21_X1  g764(.A(G197gat), .B1(new_n965), .B2(new_n568), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n910), .A2(new_n912), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n695), .A2(new_n727), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT57), .B1(new_n969), .B2(new_n710), .ZN(new_n970));
  INV_X1    g769(.A(new_n915), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n936), .A2(new_n504), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n727), .A2(new_n206), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n966), .B1(new_n974), .B2(new_n975), .ZN(G1352gat));
  NAND3_X1  g775(.A1(new_n965), .A2(new_n204), .A3(new_n692), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT62), .Z(new_n978));
  NOR3_X1   g777(.A1(new_n972), .A2(new_n693), .A3(new_n973), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n979), .B2(new_n204), .ZN(G1353gat));
  INV_X1    g779(.A(G211gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n981), .A3(new_n672), .ZN(new_n982));
  INV_X1    g781(.A(new_n973), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n672), .B(new_n983), .C1(new_n970), .C2(new_n971), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(G1354gat));
  INV_X1    g786(.A(G218gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n965), .A2(new_n988), .A3(new_n721), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n972), .A2(new_n624), .A3(new_n973), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n990), .B2(new_n988), .ZN(G1355gat));
endmodule


