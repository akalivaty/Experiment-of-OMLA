

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775;

  BUF_X1 U371 ( .A(n694), .Z(n704) );
  AND2_X1 U372 ( .A1(n375), .A2(n580), .ZN(n378) );
  AND2_X1 U373 ( .A1(n557), .A2(n556), .ZN(n403) );
  XNOR2_X1 U374 ( .A(n394), .B(KEYINPUT39), .ZN(n420) );
  INV_X1 U375 ( .A(n615), .ZN(n717) );
  XNOR2_X1 U376 ( .A(n485), .B(n484), .ZN(n542) );
  XNOR2_X1 U377 ( .A(n434), .B(n433), .ZN(n465) );
  XNOR2_X1 U378 ( .A(n429), .B(KEYINPUT3), .ZN(n434) );
  XNOR2_X2 U379 ( .A(n401), .B(n356), .ZN(n648) );
  XNOR2_X2 U380 ( .A(n350), .B(n454), .ZN(n568) );
  NAND2_X1 U381 ( .A1(n611), .A2(n452), .ZN(n350) );
  NAND2_X1 U382 ( .A1(n685), .A2(n364), .ZN(n607) );
  XNOR2_X2 U383 ( .A(n417), .B(KEYINPUT40), .ZN(n685) );
  XNOR2_X2 U384 ( .A(n351), .B(KEYINPUT96), .ZN(n598) );
  NAND2_X1 U385 ( .A1(n726), .A2(n594), .ZN(n351) );
  NOR2_X1 U386 ( .A1(G953), .A2(G237), .ZN(n514) );
  INV_X2 U387 ( .A(G953), .ZN(n771) );
  NOR2_X2 U388 ( .A1(n648), .A2(n640), .ZN(n353) );
  OR2_X2 U389 ( .A1(n707), .A2(G902), .ZN(n503) );
  XNOR2_X2 U390 ( .A(G119), .B(KEYINPUT92), .ZN(n429) );
  XNOR2_X2 U391 ( .A(n424), .B(n355), .ZN(n401) );
  NAND2_X1 U392 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U393 ( .A1(n374), .A2(n555), .ZN(n377) );
  NAND2_X1 U394 ( .A1(n420), .A2(n717), .ZN(n417) );
  NAND2_X1 U395 ( .A1(n404), .A2(n590), .ZN(n379) );
  XNOR2_X1 U396 ( .A(n609), .B(KEYINPUT110), .ZN(n682) );
  NAND2_X1 U397 ( .A1(n407), .A2(n406), .ZN(n394) );
  AND2_X1 U398 ( .A1(n370), .A2(n430), .ZN(n368) );
  OR2_X1 U399 ( .A1(n561), .A2(n562), .ZN(n615) );
  XNOR2_X1 U400 ( .A(n418), .B(G140), .ZN(n491) );
  XNOR2_X2 U401 ( .A(n353), .B(n443), .ZN(n352) );
  INV_X1 U402 ( .A(n352), .ZN(n614) );
  XNOR2_X1 U403 ( .A(n594), .B(KEYINPUT1), .ZN(n727) );
  BUF_X1 U404 ( .A(n415), .Z(n354) );
  XNOR2_X2 U405 ( .A(n426), .B(n425), .ZN(n694) );
  XNOR2_X2 U406 ( .A(n605), .B(KEYINPUT75), .ZN(n407) );
  XNOR2_X1 U407 ( .A(n465), .B(n435), .ZN(n424) );
  XNOR2_X1 U408 ( .A(n619), .B(KEYINPUT108), .ZN(n634) );
  AND2_X1 U409 ( .A1(n724), .A2(n644), .ZN(n382) );
  INV_X1 U410 ( .A(G137), .ZN(n418) );
  XNOR2_X1 U411 ( .A(G146), .B(G101), .ZN(n497) );
  NAND2_X1 U412 ( .A1(n431), .A2(KEYINPUT36), .ZN(n390) );
  XNOR2_X1 U413 ( .A(n550), .B(KEYINPUT65), .ZN(n404) );
  NOR2_X1 U414 ( .A1(n725), .A2(n393), .ZN(n398) );
  INV_X1 U415 ( .A(n395), .ZN(n393) );
  NAND2_X1 U416 ( .A1(n372), .A2(KEYINPUT34), .ZN(n366) );
  INV_X1 U417 ( .A(KEYINPUT46), .ZN(n606) );
  XNOR2_X1 U418 ( .A(G137), .B(G113), .ZN(n459) );
  XOR2_X1 U419 ( .A(G116), .B(G146), .Z(n456) );
  XNOR2_X1 U420 ( .A(G101), .B(KEYINPUT70), .ZN(n433) );
  XNOR2_X1 U421 ( .A(G122), .B(G113), .ZN(n436) );
  XNOR2_X1 U422 ( .A(n471), .B(n470), .ZN(n525) );
  XNOR2_X1 U423 ( .A(KEYINPUT82), .B(KEYINPUT8), .ZN(n470) );
  AND2_X1 U424 ( .A1(n771), .A2(G234), .ZN(n471) );
  XNOR2_X1 U425 ( .A(G116), .B(G107), .ZN(n526) );
  XNOR2_X1 U426 ( .A(KEYINPUT100), .B(KEYINPUT11), .ZN(n508) );
  XOR2_X1 U427 ( .A(G140), .B(KEYINPUT99), .Z(n509) );
  NAND2_X1 U428 ( .A1(n395), .A2(n382), .ZN(n381) );
  INV_X1 U429 ( .A(KEYINPUT64), .ZN(n425) );
  XNOR2_X1 U430 ( .A(G146), .B(G125), .ZN(n476) );
  NAND2_X1 U431 ( .A1(n670), .A2(n642), .ZN(n724) );
  XNOR2_X1 U432 ( .A(n352), .B(n365), .ZN(n406) );
  INV_X1 U433 ( .A(KEYINPUT38), .ZN(n365) );
  INV_X1 U434 ( .A(KEYINPUT95), .ZN(n414) );
  XNOR2_X1 U435 ( .A(G128), .B(G119), .ZN(n472) );
  XNOR2_X1 U436 ( .A(n476), .B(KEYINPUT10), .ZN(n671) );
  XNOR2_X1 U437 ( .A(G134), .B(G122), .ZN(n530) );
  NAND2_X1 U438 ( .A1(n410), .A2(n408), .ZN(n758) );
  NAND2_X1 U439 ( .A1(n409), .A2(n412), .ZN(n408) );
  AND2_X1 U440 ( .A1(n411), .A2(n413), .ZN(n410) );
  OR2_X1 U441 ( .A1(n548), .A2(n731), .ZN(n543) );
  XNOR2_X1 U442 ( .A(n446), .B(KEYINPUT19), .ZN(n611) );
  NAND2_X1 U443 ( .A1(n352), .A2(n445), .ZN(n446) );
  INV_X1 U444 ( .A(KEYINPUT22), .ZN(n428) );
  XNOR2_X1 U445 ( .A(n672), .B(n500), .ZN(n707) );
  XNOR2_X1 U446 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U447 ( .A(n416), .B(KEYINPUT42), .ZN(n364) );
  NAND2_X1 U448 ( .A1(n758), .A2(n610), .ZN(n416) );
  OR2_X1 U449 ( .A1(n431), .A2(KEYINPUT36), .ZN(n392) );
  NAND2_X1 U450 ( .A1(n396), .A2(n762), .ZN(n763) );
  INV_X1 U451 ( .A(G140), .ZN(n721) );
  INV_X1 U452 ( .A(G122), .ZN(n400) );
  INV_X1 U453 ( .A(G110), .ZN(n380) );
  XOR2_X1 U454 ( .A(n513), .B(n494), .Z(n355) );
  XOR2_X1 U455 ( .A(n464), .B(n440), .Z(n356) );
  XNOR2_X1 U456 ( .A(n582), .B(KEYINPUT112), .ZN(n742) );
  NOR2_X1 U457 ( .A1(n598), .A2(n560), .ZN(n357) );
  NOR2_X1 U458 ( .A1(n544), .A2(n618), .ZN(n358) );
  AND2_X1 U459 ( .A1(n352), .A2(n608), .ZN(n359) );
  XNOR2_X1 U460 ( .A(n583), .B(KEYINPUT41), .ZN(n360) );
  BUF_X1 U461 ( .A(n542), .Z(n731) );
  XOR2_X1 U462 ( .A(KEYINPUT85), .B(KEYINPUT35), .Z(n361) );
  INV_X1 U463 ( .A(n665), .ZN(n419) );
  AND2_X1 U464 ( .A1(n640), .A2(KEYINPUT2), .ZN(n362) );
  OR2_X1 U465 ( .A1(n406), .A2(n445), .ZN(n747) );
  NAND2_X1 U466 ( .A1(n406), .A2(n445), .ZN(n582) );
  XNOR2_X1 U467 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X2 U468 ( .A(n426), .B(n425), .ZN(n363) );
  NAND2_X2 U469 ( .A1(n423), .A2(n405), .ZN(n426) );
  NAND2_X1 U470 ( .A1(n647), .A2(n642), .ZN(n395) );
  XNOR2_X1 U471 ( .A(n364), .B(G137), .ZN(G39) );
  NAND2_X2 U472 ( .A1(n367), .A2(n366), .ZN(n373) );
  AND2_X2 U473 ( .A1(n369), .A2(n368), .ZN(n367) );
  NAND2_X1 U474 ( .A1(n371), .A2(n506), .ZN(n369) );
  OR2_X1 U475 ( .A1(n757), .A2(n507), .ZN(n370) );
  AND2_X1 U476 ( .A1(n757), .A2(n507), .ZN(n371) );
  INV_X1 U477 ( .A(n506), .ZN(n372) );
  XNOR2_X2 U478 ( .A(n373), .B(n361), .ZN(n538) );
  NAND2_X1 U479 ( .A1(n553), .A2(n554), .ZN(n374) );
  NAND2_X1 U480 ( .A1(n558), .A2(n399), .ZN(n375) );
  XNOR2_X2 U481 ( .A(n376), .B(n581), .ZN(n647) );
  NAND2_X1 U482 ( .A1(n403), .A2(n379), .ZN(n402) );
  INV_X1 U483 ( .A(n379), .ZN(n551) );
  XNOR2_X1 U484 ( .A(n551), .B(n380), .ZN(G12) );
  NAND2_X1 U485 ( .A1(n383), .A2(n381), .ZN(n423) );
  NAND2_X1 U486 ( .A1(n384), .A2(KEYINPUT67), .ZN(n383) );
  NAND2_X1 U487 ( .A1(n385), .A2(n362), .ZN(n384) );
  INV_X1 U488 ( .A(n641), .ZN(n385) );
  XNOR2_X1 U489 ( .A(n492), .B(n386), .ZN(n687) );
  XNOR2_X2 U490 ( .A(n464), .B(n463), .ZN(n492) );
  XNOR2_X2 U491 ( .A(n527), .B(KEYINPUT4), .ZN(n464) );
  XNOR2_X1 U492 ( .A(n465), .B(n466), .ZN(n386) );
  NAND2_X1 U493 ( .A1(n387), .A2(n392), .ZN(n620) );
  NAND2_X1 U494 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U495 ( .A1(n634), .A2(KEYINPUT36), .ZN(n388) );
  NAND2_X1 U496 ( .A1(n391), .A2(n390), .ZN(n389) );
  INV_X1 U497 ( .A(n634), .ZN(n391) );
  NAND2_X1 U498 ( .A1(n397), .A2(n405), .ZN(n396) );
  XNOR2_X1 U499 ( .A(n398), .B(KEYINPUT80), .ZN(n397) );
  INV_X1 U500 ( .A(n538), .ZN(n399) );
  XNOR2_X1 U501 ( .A(n538), .B(n400), .ZN(G24) );
  XNOR2_X1 U502 ( .A(n401), .B(KEYINPUT127), .ZN(n773) );
  NAND2_X1 U503 ( .A1(n402), .A2(KEYINPUT88), .ZN(n558) );
  XNOR2_X2 U504 ( .A(n547), .B(n546), .ZN(n557) );
  NAND2_X1 U505 ( .A1(n422), .A2(n421), .ZN(n405) );
  NAND2_X1 U506 ( .A1(n407), .A2(n359), .ZN(n609) );
  XNOR2_X1 U507 ( .A(n646), .B(n427), .ZN(n422) );
  NAND2_X2 U508 ( .A1(n639), .A2(n638), .ZN(n670) );
  INV_X1 U509 ( .A(n742), .ZN(n409) );
  NAND2_X1 U510 ( .A1(n742), .A2(n360), .ZN(n411) );
  NOR2_X1 U511 ( .A1(n745), .A2(n360), .ZN(n412) );
  NAND2_X1 U512 ( .A1(n745), .A2(n360), .ZN(n413) );
  NAND2_X1 U513 ( .A1(n506), .A2(n357), .ZN(n565) );
  XNOR2_X1 U514 ( .A(n568), .B(n414), .ZN(n506) );
  NAND2_X1 U515 ( .A1(n358), .A2(n415), .ZN(n547) );
  NAND2_X1 U516 ( .A1(n415), .A2(n549), .ZN(n550) );
  NAND2_X1 U517 ( .A1(n354), .A2(n567), .ZN(n669) );
  XNOR2_X2 U518 ( .A(n541), .B(n428), .ZN(n415) );
  NAND2_X1 U519 ( .A1(n420), .A2(n419), .ZN(n681) );
  XNOR2_X2 U520 ( .A(n492), .B(n491), .ZN(n672) );
  INV_X1 U521 ( .A(n766), .ZN(n421) );
  INV_X1 U522 ( .A(KEYINPUT84), .ZN(n427) );
  BUF_X1 U523 ( .A(n647), .Z(n766) );
  XNOR2_X2 U524 ( .A(n469), .B(n468), .ZN(n734) );
  XOR2_X1 U525 ( .A(n537), .B(KEYINPUT78), .Z(n430) );
  NOR2_X1 U526 ( .A1(n614), .A2(n633), .ZN(n431) );
  XOR2_X1 U527 ( .A(n540), .B(KEYINPUT105), .Z(n432) );
  NAND2_X1 U528 ( .A1(n538), .A2(KEYINPUT88), .ZN(n554) );
  INV_X1 U529 ( .A(KEYINPUT68), .ZN(n626) );
  INV_X1 U530 ( .A(KEYINPUT5), .ZN(n458) );
  XNOR2_X1 U531 ( .A(n459), .B(n458), .ZN(n460) );
  AND2_X2 U532 ( .A1(n542), .A2(n730), .ZN(n726) );
  XNOR2_X1 U533 ( .A(n461), .B(n460), .ZN(n466) );
  INV_X1 U534 ( .A(KEYINPUT34), .ZN(n507) );
  INV_X1 U535 ( .A(KEYINPUT60), .ZN(n663) );
  XNOR2_X1 U536 ( .A(n526), .B(KEYINPUT16), .ZN(n435) );
  XNOR2_X1 U537 ( .A(n436), .B(G104), .ZN(n513) );
  XNOR2_X1 U538 ( .A(KEYINPUT74), .B(G110), .ZN(n494) );
  XNOR2_X2 U539 ( .A(G143), .B(G128), .ZN(n527) );
  XNOR2_X1 U540 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n438) );
  NAND2_X1 U541 ( .A1(n771), .A2(G224), .ZN(n437) );
  XNOR2_X1 U542 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U543 ( .A(n476), .B(n439), .ZN(n440) );
  XNOR2_X1 U544 ( .A(G902), .B(KEYINPUT15), .ZN(n643) );
  INV_X1 U545 ( .A(n643), .ZN(n640) );
  NOR2_X1 U546 ( .A1(G902), .A2(G237), .ZN(n441) );
  XNOR2_X1 U547 ( .A(n441), .B(KEYINPUT73), .ZN(n444) );
  AND2_X1 U548 ( .A1(n444), .A2(G210), .ZN(n442) );
  XNOR2_X1 U549 ( .A(n442), .B(KEYINPUT93), .ZN(n443) );
  AND2_X1 U550 ( .A1(n444), .A2(G214), .ZN(n744) );
  INV_X1 U551 ( .A(n744), .ZN(n445) );
  NAND2_X1 U552 ( .A1(G234), .A2(G237), .ZN(n447) );
  XNOR2_X1 U553 ( .A(n447), .B(KEYINPUT94), .ZN(n448) );
  XNOR2_X1 U554 ( .A(KEYINPUT14), .B(n448), .ZN(n450) );
  AND2_X1 U555 ( .A1(n450), .A2(G953), .ZN(n449) );
  NAND2_X1 U556 ( .A1(G902), .A2(n449), .ZN(n584) );
  OR2_X1 U557 ( .A1(n584), .A2(G898), .ZN(n451) );
  NAND2_X1 U558 ( .A1(G952), .A2(n450), .ZN(n755) );
  OR2_X1 U559 ( .A1(n755), .A2(G953), .ZN(n586) );
  NAND2_X1 U560 ( .A1(n451), .A2(n586), .ZN(n452) );
  INV_X1 U561 ( .A(KEYINPUT90), .ZN(n453) );
  XNOR2_X1 U562 ( .A(n453), .B(KEYINPUT0), .ZN(n454) );
  NAND2_X1 U563 ( .A1(n514), .A2(G210), .ZN(n457) );
  XNOR2_X1 U564 ( .A(n457), .B(n456), .ZN(n461) );
  INV_X1 U565 ( .A(G134), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n462), .B(G131), .ZN(n463) );
  INV_X1 U567 ( .A(G902), .ZN(n520) );
  NAND2_X1 U568 ( .A1(n687), .A2(n520), .ZN(n469) );
  INV_X1 U569 ( .A(KEYINPUT72), .ZN(n467) );
  XNOR2_X1 U570 ( .A(n467), .B(G472), .ZN(n468) );
  XNOR2_X1 U571 ( .A(n734), .B(KEYINPUT6), .ZN(n618) );
  NAND2_X1 U572 ( .A1(n525), .A2(G221), .ZN(n475) );
  XNOR2_X1 U573 ( .A(n472), .B(KEYINPUT76), .ZN(n473) );
  XNOR2_X1 U574 ( .A(n473), .B(n491), .ZN(n474) );
  XNOR2_X1 U575 ( .A(n475), .B(n474), .ZN(n481) );
  XNOR2_X1 U576 ( .A(G110), .B(KEYINPUT23), .ZN(n478) );
  XNOR2_X1 U577 ( .A(KEYINPUT24), .B(KEYINPUT71), .ZN(n477) );
  XNOR2_X1 U578 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U579 ( .A(n671), .B(n479), .ZN(n480) );
  XNOR2_X1 U580 ( .A(n481), .B(n480), .ZN(n695) );
  OR2_X2 U581 ( .A1(n695), .A2(G902), .ZN(n485) );
  NAND2_X1 U582 ( .A1(n643), .A2(G234), .ZN(n482) );
  XNOR2_X1 U583 ( .A(n482), .B(KEYINPUT20), .ZN(n486) );
  AND2_X1 U584 ( .A1(n486), .A2(G217), .ZN(n483) );
  XNOR2_X1 U585 ( .A(n483), .B(KEYINPUT25), .ZN(n484) );
  INV_X1 U586 ( .A(n486), .ZN(n488) );
  INV_X1 U587 ( .A(G221), .ZN(n487) );
  OR2_X1 U588 ( .A1(n488), .A2(n487), .ZN(n490) );
  INV_X1 U589 ( .A(KEYINPUT21), .ZN(n489) );
  XNOR2_X1 U590 ( .A(n490), .B(n489), .ZN(n730) );
  AND2_X1 U591 ( .A1(n618), .A2(n726), .ZN(n504) );
  NAND2_X1 U592 ( .A1(n771), .A2(G227), .ZN(n493) );
  XNOR2_X1 U593 ( .A(n493), .B(KEYINPUT77), .ZN(n495) );
  XNOR2_X1 U594 ( .A(n495), .B(n494), .ZN(n499) );
  XNOR2_X1 U595 ( .A(G107), .B(G104), .ZN(n496) );
  XNOR2_X1 U596 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U597 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U598 ( .A(KEYINPUT69), .ZN(n501) );
  XNOR2_X1 U599 ( .A(n501), .B(G469), .ZN(n502) );
  XNOR2_X2 U600 ( .A(n503), .B(n502), .ZN(n594) );
  NAND2_X1 U601 ( .A1(n504), .A2(n727), .ZN(n505) );
  XNOR2_X1 U602 ( .A(n505), .B(KEYINPUT33), .ZN(n757) );
  XNOR2_X1 U603 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U604 ( .A(n510), .B(KEYINPUT12), .Z(n512) );
  XNOR2_X1 U605 ( .A(G143), .B(G131), .ZN(n511) );
  XNOR2_X1 U606 ( .A(n512), .B(n511), .ZN(n519) );
  INV_X1 U607 ( .A(n513), .ZN(n516) );
  NAND2_X1 U608 ( .A1(G214), .A2(n514), .ZN(n515) );
  XNOR2_X1 U609 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U610 ( .A(n517), .B(n671), .ZN(n518) );
  XNOR2_X1 U611 ( .A(n519), .B(n518), .ZN(n659) );
  NAND2_X1 U612 ( .A1(n659), .A2(n520), .ZN(n524) );
  XOR2_X1 U613 ( .A(KEYINPUT102), .B(KEYINPUT13), .Z(n522) );
  XNOR2_X1 U614 ( .A(KEYINPUT101), .B(G475), .ZN(n521) );
  XNOR2_X1 U615 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U616 ( .A(n524), .B(n523), .ZN(n561) );
  INV_X1 U617 ( .A(n561), .ZN(n564) );
  NAND2_X1 U618 ( .A1(n525), .A2(G217), .ZN(n529) );
  XNOR2_X1 U619 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U620 ( .A(n529), .B(n528), .ZN(n534) );
  XOR2_X1 U621 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n532) );
  XNOR2_X1 U622 ( .A(n530), .B(KEYINPUT9), .ZN(n531) );
  XNOR2_X1 U623 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U624 ( .A(n534), .B(n533), .ZN(n700) );
  OR2_X1 U625 ( .A1(n700), .A2(G902), .ZN(n536) );
  XNOR2_X1 U626 ( .A(KEYINPUT104), .B(G478), .ZN(n535) );
  XNOR2_X1 U627 ( .A(n536), .B(n535), .ZN(n562) );
  AND2_X1 U628 ( .A1(n564), .A2(n562), .ZN(n608) );
  INV_X1 U629 ( .A(n608), .ZN(n537) );
  OR2_X1 U630 ( .A1(n564), .A2(n562), .ZN(n745) );
  INV_X1 U631 ( .A(n730), .ZN(n539) );
  NOR2_X1 U632 ( .A1(n745), .A2(n539), .ZN(n540) );
  NAND2_X1 U633 ( .A1(n568), .A2(n432), .ZN(n541) );
  INV_X1 U634 ( .A(n727), .ZN(n548) );
  XNOR2_X1 U635 ( .A(n543), .B(KEYINPUT106), .ZN(n544) );
  INV_X1 U636 ( .A(KEYINPUT79), .ZN(n545) );
  XNOR2_X1 U637 ( .A(n545), .B(KEYINPUT32), .ZN(n546) );
  NAND2_X1 U638 ( .A1(n557), .A2(KEYINPUT44), .ZN(n552) );
  AND2_X1 U639 ( .A1(n548), .A2(n734), .ZN(n549) );
  NOR2_X1 U640 ( .A1(n552), .A2(n551), .ZN(n553) );
  INV_X1 U641 ( .A(KEYINPUT44), .ZN(n556) );
  NAND2_X1 U642 ( .A1(n556), .A2(KEYINPUT88), .ZN(n555) );
  INV_X1 U643 ( .A(n734), .ZN(n560) );
  OR2_X1 U644 ( .A1(n565), .A2(n615), .ZN(n712) );
  INV_X1 U645 ( .A(n562), .ZN(n563) );
  OR2_X1 U646 ( .A1(n564), .A2(n563), .ZN(n665) );
  OR2_X1 U647 ( .A1(n565), .A2(n665), .ZN(n713) );
  NAND2_X1 U648 ( .A1(n712), .A2(n713), .ZN(n579) );
  INV_X1 U649 ( .A(n731), .ZN(n590) );
  OR2_X1 U650 ( .A1(n618), .A2(n590), .ZN(n566) );
  NOR2_X1 U651 ( .A1(n566), .A2(n727), .ZN(n567) );
  INV_X1 U652 ( .A(n568), .ZN(n572) );
  INV_X1 U653 ( .A(n726), .ZN(n569) );
  NOR2_X1 U654 ( .A1(n734), .A2(n569), .ZN(n570) );
  AND2_X1 U655 ( .A1(n727), .A2(n570), .ZN(n738) );
  INV_X1 U656 ( .A(n738), .ZN(n571) );
  OR2_X1 U657 ( .A1(n572), .A2(n571), .ZN(n576) );
  XNOR2_X1 U658 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n574) );
  INV_X1 U659 ( .A(KEYINPUT97), .ZN(n573) );
  XNOR2_X1 U660 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U661 ( .A(n576), .B(n575), .ZN(n679) );
  NAND2_X1 U662 ( .A1(n615), .A2(n665), .ZN(n743) );
  NAND2_X1 U663 ( .A1(n679), .A2(n743), .ZN(n577) );
  NAND2_X1 U664 ( .A1(n669), .A2(n577), .ZN(n578) );
  NOR2_X1 U665 ( .A1(n579), .A2(n578), .ZN(n580) );
  INV_X1 U666 ( .A(KEYINPUT45), .ZN(n581) );
  INV_X1 U667 ( .A(KEYINPUT113), .ZN(n583) );
  NOR2_X1 U668 ( .A1(G900), .A2(n584), .ZN(n585) );
  XOR2_X1 U669 ( .A(KEYINPUT107), .B(n585), .Z(n588) );
  INV_X1 U670 ( .A(n586), .ZN(n587) );
  NOR2_X1 U671 ( .A1(n588), .A2(n587), .ZN(n601) );
  INV_X1 U672 ( .A(n601), .ZN(n589) );
  AND2_X1 U673 ( .A1(n589), .A2(n730), .ZN(n591) );
  NAND2_X1 U674 ( .A1(n591), .A2(n590), .ZN(n616) );
  OR2_X1 U675 ( .A1(n734), .A2(n616), .ZN(n593) );
  INV_X1 U676 ( .A(KEYINPUT28), .ZN(n592) );
  XNOR2_X1 U677 ( .A(n593), .B(n592), .ZN(n597) );
  INV_X1 U678 ( .A(n594), .ZN(n595) );
  XNOR2_X1 U679 ( .A(n595), .B(KEYINPUT111), .ZN(n596) );
  AND2_X1 U680 ( .A1(n597), .A2(n596), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n598), .B(KEYINPUT109), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n734), .A2(n744), .ZN(n600) );
  INV_X1 U683 ( .A(KEYINPUT30), .ZN(n599) );
  XNOR2_X1 U684 ( .A(n600), .B(n599), .ZN(n602) );
  NOR2_X1 U685 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U687 ( .A(n607), .B(n606), .ZN(n629) );
  AND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n718) );
  NAND2_X1 U689 ( .A1(n718), .A2(n743), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n621), .A2(KEYINPUT47), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n682), .A2(n612), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n613), .B(KEYINPUT81), .ZN(n625) );
  NAND2_X1 U693 ( .A1(n717), .A2(n445), .ZN(n633) );
  INV_X1 U694 ( .A(n616), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n620), .A2(n727), .ZN(n684) );
  XNOR2_X1 U697 ( .A(n684), .B(KEYINPUT87), .ZN(n623) );
  NOR2_X1 U698 ( .A1(n621), .A2(KEYINPUT47), .ZN(n622) );
  NOR2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n632) );
  INV_X1 U703 ( .A(KEYINPUT86), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n630), .B(KEYINPUT48), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n632), .B(n631), .ZN(n639) );
  OR2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n635) );
  OR2_X1 U707 ( .A1(n635), .A2(n727), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n636), .B(KEYINPUT43), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n637), .A2(n614), .ZN(n722) );
  AND2_X1 U710 ( .A1(n681), .A2(n722), .ZN(n638) );
  NOR2_X1 U711 ( .A1(n647), .A2(n670), .ZN(n641) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n642) );
  NOR2_X1 U713 ( .A1(n643), .A2(KEYINPUT67), .ZN(n644) );
  INV_X1 U714 ( .A(n670), .ZN(n645) );
  NAND2_X1 U715 ( .A1(n645), .A2(KEYINPUT2), .ZN(n646) );
  NAND2_X1 U716 ( .A1(n363), .A2(G210), .ZN(n652) );
  BUF_X1 U717 ( .A(n648), .Z(n650) );
  XNOR2_X1 U718 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n652), .B(n651), .ZN(n654) );
  INV_X1 U720 ( .A(G952), .ZN(n653) );
  NAND2_X1 U721 ( .A1(n653), .A2(G953), .ZN(n698) );
  NAND2_X1 U722 ( .A1(n654), .A2(n698), .ZN(n656) );
  INV_X1 U723 ( .A(KEYINPUT56), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(G51) );
  NAND2_X1 U725 ( .A1(n363), .A2(G475), .ZN(n661) );
  XNOR2_X1 U726 ( .A(KEYINPUT66), .B(KEYINPUT124), .ZN(n657) );
  XOR2_X1 U727 ( .A(n657), .B(KEYINPUT59), .Z(n658) );
  XNOR2_X1 U728 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U729 ( .A1(n662), .A2(n698), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n664), .B(n663), .ZN(G60) );
  NAND2_X1 U731 ( .A1(n718), .A2(n419), .ZN(n667) );
  XOR2_X1 U732 ( .A(G128), .B(KEYINPUT29), .Z(n666) );
  XNOR2_X1 U733 ( .A(n667), .B(n666), .ZN(G30) );
  NAND2_X1 U734 ( .A1(n679), .A2(n717), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n668), .B(G113), .ZN(G15) );
  XNOR2_X1 U736 ( .A(n669), .B(G101), .ZN(G3) );
  XOR2_X1 U737 ( .A(n672), .B(n671), .Z(n674) );
  XNOR2_X1 U738 ( .A(n670), .B(n674), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n673), .A2(n771), .ZN(n678) );
  XNOR2_X1 U740 ( .A(n674), .B(G227), .ZN(n675) );
  NAND2_X1 U741 ( .A1(n675), .A2(G900), .ZN(n676) );
  NAND2_X1 U742 ( .A1(n676), .A2(G953), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n678), .A2(n677), .ZN(G72) );
  NAND2_X1 U744 ( .A1(n679), .A2(n419), .ZN(n680) );
  XNOR2_X1 U745 ( .A(n680), .B(G116), .ZN(G18) );
  XNOR2_X1 U746 ( .A(n681), .B(G134), .ZN(G36) );
  XNOR2_X1 U747 ( .A(n682), .B(G143), .ZN(G45) );
  XOR2_X1 U748 ( .A(G125), .B(KEYINPUT37), .Z(n683) );
  XNOR2_X1 U749 ( .A(n684), .B(n683), .ZN(G27) );
  XNOR2_X1 U750 ( .A(n557), .B(G119), .ZN(G21) );
  XNOR2_X1 U751 ( .A(n685), .B(G131), .ZN(G33) );
  NAND2_X1 U752 ( .A1(n694), .A2(G472), .ZN(n689) );
  XOR2_X1 U753 ( .A(KEYINPUT91), .B(KEYINPUT62), .Z(n686) );
  XNOR2_X1 U754 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U755 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U756 ( .A1(n690), .A2(n698), .ZN(n693) );
  XOR2_X1 U757 ( .A(KEYINPUT114), .B(KEYINPUT63), .Z(n691) );
  XNOR2_X1 U758 ( .A(n691), .B(KEYINPUT89), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n693), .B(n692), .ZN(G57) );
  NAND2_X1 U760 ( .A1(n704), .A2(G217), .ZN(n697) );
  XNOR2_X1 U761 ( .A(n695), .B(KEYINPUT126), .ZN(n696) );
  XNOR2_X1 U762 ( .A(n697), .B(n696), .ZN(n699) );
  INV_X1 U763 ( .A(n698), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n699), .A2(n710), .ZN(G66) );
  NAND2_X1 U765 ( .A1(n704), .A2(G478), .ZN(n702) );
  XOR2_X1 U766 ( .A(KEYINPUT125), .B(n700), .Z(n701) );
  XNOR2_X1 U767 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U768 ( .A1(n703), .A2(n710), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n704), .A2(G469), .ZN(n709) );
  XNOR2_X1 U770 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n705) );
  XNOR2_X1 U771 ( .A(n705), .B(KEYINPUT57), .ZN(n706) );
  XNOR2_X1 U772 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U773 ( .A(n709), .B(n708), .ZN(n711) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(G54) );
  XNOR2_X1 U775 ( .A(G104), .B(n712), .ZN(G6) );
  XOR2_X1 U776 ( .A(KEYINPUT115), .B(KEYINPUT26), .Z(n714) );
  XNOR2_X1 U777 ( .A(n714), .B(n713), .ZN(n716) );
  XOR2_X1 U778 ( .A(G107), .B(KEYINPUT27), .Z(n715) );
  XNOR2_X1 U779 ( .A(n716), .B(n715), .ZN(G9) );
  NAND2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U781 ( .A(n719), .B(KEYINPUT116), .ZN(n720) );
  XNOR2_X1 U782 ( .A(G146), .B(n720), .ZN(G48) );
  XNOR2_X1 U783 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U784 ( .A(n723), .B(KEYINPUT117), .ZN(G42) );
  XNOR2_X1 U785 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n765) );
  XNOR2_X1 U786 ( .A(n724), .B(KEYINPUT83), .ZN(n725) );
  NOR2_X1 U787 ( .A1(n727), .A2(n726), .ZN(n729) );
  XNOR2_X1 U788 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n728) );
  XNOR2_X1 U789 ( .A(n729), .B(n728), .ZN(n736) );
  NOR2_X1 U790 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U791 ( .A(n732), .B(KEYINPUT49), .ZN(n733) );
  NAND2_X1 U792 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U793 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U794 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U795 ( .A(n739), .B(KEYINPUT51), .Z(n740) );
  XNOR2_X1 U796 ( .A(KEYINPUT119), .B(n740), .ZN(n741) );
  NAND2_X1 U797 ( .A1(n741), .A2(n758), .ZN(n752) );
  NAND2_X1 U798 ( .A1(n409), .A2(n743), .ZN(n749) );
  INV_X1 U799 ( .A(n745), .ZN(n746) );
  NAND2_X1 U800 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U801 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U802 ( .A1(n750), .A2(n757), .ZN(n751) );
  NAND2_X1 U803 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U804 ( .A(KEYINPUT52), .B(n753), .Z(n754) );
  NOR2_X1 U805 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U806 ( .A(n756), .B(KEYINPUT120), .ZN(n761) );
  NAND2_X1 U807 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U808 ( .A1(n759), .A2(n771), .ZN(n760) );
  NOR2_X1 U809 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U810 ( .A(n763), .B(KEYINPUT53), .ZN(n764) );
  XNOR2_X1 U811 ( .A(n765), .B(n764), .ZN(G75) );
  NAND2_X1 U812 ( .A1(n421), .A2(n771), .ZN(n770) );
  NAND2_X1 U813 ( .A1(G953), .A2(G224), .ZN(n767) );
  XNOR2_X1 U814 ( .A(KEYINPUT61), .B(n767), .ZN(n768) );
  NAND2_X1 U815 ( .A1(n768), .A2(G898), .ZN(n769) );
  NAND2_X1 U816 ( .A1(n770), .A2(n769), .ZN(n775) );
  NOR2_X1 U817 ( .A1(n771), .A2(G898), .ZN(n772) );
  NOR2_X1 U818 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U819 ( .A(n775), .B(n774), .ZN(G69) );
endmodule

