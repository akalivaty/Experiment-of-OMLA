//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT2), .A2(G113), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT66), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT2), .A3(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G116), .B(G119), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n194), .B2(new_n197), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n192), .B1(KEYINPUT2), .B2(G113), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n190), .A2(KEYINPUT66), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n197), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n198), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n191), .A2(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n198), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT68), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G137), .ZN(new_n213));
  AOI21_X1  g027(.A(G131), .B1(new_n212), .B2(G137), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT11), .A3(G134), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT64), .A4(new_n216), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n213), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n219), .A2(new_n220), .B1(G131), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G143), .B(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G146), .ZN(new_n230));
  OR2_X1    g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n228), .A2(new_n230), .B1(new_n231), .B2(new_n225), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  OAI22_X1  g047(.A1(new_n202), .A2(new_n210), .B1(new_n223), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n228), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n224), .B1(new_n237), .B2(G128), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n230), .A3(G128), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT67), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G131), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n215), .A2(G134), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(new_n221), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n219), .B2(new_n220), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n235), .A2(new_n236), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n224), .A3(G128), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n240), .B2(new_n228), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n247), .B(new_n249), .C1(new_n251), .C2(new_n224), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n242), .A2(new_n246), .A3(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(new_n234), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n219), .A2(new_n220), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n222), .A2(G131), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n224), .A2(new_n225), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n231), .A2(new_n225), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n224), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n242), .A2(new_n246), .A3(new_n252), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n201), .B1(new_n199), .B2(new_n200), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n207), .A2(KEYINPUT68), .A3(new_n209), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n261), .A2(new_n262), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n207), .A2(new_n209), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n249), .B1(new_n251), .B2(new_n224), .ZN(new_n269));
  INV_X1    g083(.A(new_n245), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n269), .A2(new_n255), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n233), .B1(new_n255), .B2(new_n256), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n254), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT28), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n234), .A2(new_n253), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(KEYINPUT28), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(G237), .A2(G953), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G210), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT27), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT26), .B(G101), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n254), .A2(new_n267), .A3(new_n284), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n271), .B2(new_n272), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT30), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(new_n268), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(KEYINPUT31), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT31), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n254), .A2(new_n267), .A3(new_n284), .ZN(new_n294));
  INV_X1    g108(.A(new_n291), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n189), .B1(new_n286), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n187), .B1(new_n298), .B2(KEYINPUT32), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n291), .A2(new_n254), .A3(new_n267), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n285), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n275), .A2(new_n284), .A3(new_n278), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n300), .A2(KEYINPUT71), .A3(new_n285), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n264), .B(new_n263), .C1(new_n253), .C2(new_n272), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n254), .A2(new_n308), .A3(new_n267), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n277), .B1(new_n309), .B2(KEYINPUT28), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n285), .A2(new_n305), .ZN(new_n311));
  AOI21_X1  g125(.A(G902), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G472), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n298), .A2(KEYINPUT32), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT32), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n285), .A2(new_n279), .B1(new_n292), .B2(new_n296), .ZN(new_n317));
  OAI211_X1 g131(.A(KEYINPUT70), .B(new_n316), .C1(new_n317), .C2(new_n189), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n299), .A2(new_n314), .A3(new_n315), .A4(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G221), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT9), .B(G234), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G902), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT77), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G140), .ZN(new_n326));
  INV_X1    g140(.A(G953), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n327), .A2(G227), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n326), .B(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G107), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G104), .ZN(new_n332));
  INV_X1    g146(.A(G104), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G107), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n335), .A2(G101), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT3), .B1(new_n333), .B2(G107), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n331), .A3(G104), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n331), .A2(G104), .ZN(new_n341));
  AND2_X1   g155(.A1(KEYINPUT78), .A2(G101), .ZN(new_n342));
  NOR2_X1   g156(.A1(KEYINPUT78), .A2(G101), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n344), .A3(KEYINPUT79), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n337), .A2(new_n339), .ZN(new_n347));
  OR2_X1    g161(.A1(KEYINPUT78), .A2(G101), .ZN(new_n348));
  NAND2_X1  g162(.A1(KEYINPUT78), .A2(G101), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n334), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n346), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n336), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n224), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n354), .B(KEYINPUT1), .C1(new_n229), .C2(G146), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G128), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n354), .B1(new_n228), .B2(KEYINPUT1), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n249), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n345), .A2(new_n351), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n337), .A2(new_n339), .A3(new_n334), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(G101), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n363), .A3(G101), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n260), .A2(new_n367), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n360), .A2(new_n361), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n242), .A2(new_n252), .ZN(new_n371));
  AOI211_X1 g185(.A(new_n361), .B(new_n336), .C1(new_n345), .C2(new_n351), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n336), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n362), .A2(KEYINPUT10), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n242), .A2(new_n252), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT81), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n223), .B(new_n369), .C1(new_n373), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT79), .B1(new_n340), .B2(new_n344), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n347), .A2(new_n350), .A3(new_n346), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n374), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n269), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n223), .B1(new_n383), .B2(new_n360), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT12), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(KEYINPUT12), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n362), .A2(new_n359), .A3(new_n374), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n269), .B1(new_n362), .B2(new_n374), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n257), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT12), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(KEYINPUT82), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n387), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n330), .B(new_n378), .C1(new_n386), .C2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n387), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n384), .B2(new_n392), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n390), .A2(KEYINPUT82), .A3(new_n391), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n401), .A2(KEYINPUT83), .A3(new_n330), .A4(new_n378), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n371), .A2(new_n370), .A3(new_n372), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT81), .B1(new_n375), .B2(new_n376), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n405), .A2(new_n223), .A3(new_n369), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n223), .B1(new_n405), .B2(new_n369), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n329), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n397), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G469), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n323), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n323), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n330), .B1(new_n406), .B2(new_n407), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n401), .A2(new_n329), .A3(new_n378), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n412), .B1(new_n415), .B2(G469), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n325), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n364), .A2(G101), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n363), .A2(new_n419), .B1(new_n207), .B2(new_n209), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n421));
  INV_X1    g235(.A(G116), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n422), .A2(KEYINPUT5), .A3(G119), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(new_n196), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n421), .A2(new_n424), .B1(new_n208), .B2(new_n198), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n420), .A2(new_n366), .B1(new_n352), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G122), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n418), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n427), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n352), .A2(new_n425), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n362), .A2(new_n365), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n268), .A2(new_n367), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n430), .B(new_n432), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n428), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n233), .A2(KEYINPUT85), .A3(G125), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n269), .A2(G125), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  INV_X1    g254(.A(G125), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n260), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n438), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT86), .B(G224), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n327), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n445), .B(KEYINPUT87), .Z(new_n446));
  XNOR2_X1  g260(.A(new_n443), .B(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT84), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n449), .A2(new_n418), .A3(new_n435), .A4(new_n429), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n437), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(KEYINPUT7), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n443), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n432), .B(new_n427), .C1(new_n433), .C2(new_n434), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n438), .B(new_n452), .C1(new_n439), .C2(new_n442), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(KEYINPUT88), .B(KEYINPUT8), .Z(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(new_n427), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT90), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n352), .B2(new_n425), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n421), .A2(KEYINPUT89), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n424), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n421), .A2(KEYINPUT89), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n209), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n461), .B1(new_n465), .B2(new_n381), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n352), .A2(new_n460), .A3(new_n425), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(G902), .B1(new_n457), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n451), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G210), .B1(G237), .B2(G902), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(KEYINPUT91), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n472), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n451), .A2(new_n474), .A3(new_n469), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G214), .B1(G237), .B2(G902), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT94), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n229), .A2(G128), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n229), .A2(G128), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT13), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n479), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n250), .A2(G143), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n250), .A2(G143), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(KEYINPUT13), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT94), .B1(new_n480), .B2(new_n482), .ZN(new_n487));
  OAI211_X1 g301(.A(G134), .B(new_n483), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT95), .ZN(new_n489));
  INV_X1    g303(.A(G122), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G116), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n422), .A2(G122), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT93), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n491), .B2(new_n492), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n331), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n492), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT93), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(G107), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n479), .B1(new_n484), .B2(KEYINPUT13), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT95), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n504), .A2(new_n505), .A3(G134), .A4(new_n483), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n484), .A2(new_n481), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n212), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n489), .A2(new_n501), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n507), .B(new_n212), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n491), .B1(new_n492), .B2(KEYINPUT14), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n492), .A2(KEYINPUT14), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n492), .A2(KEYINPUT96), .A3(KEYINPUT14), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n510), .B(new_n496), .C1(new_n331), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G217), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n321), .A2(new_n518), .A3(G953), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n509), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT97), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT97), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n509), .A2(new_n522), .A3(new_n517), .A4(new_n519), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n519), .B1(new_n509), .B2(new_n517), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT98), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT99), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n323), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G478), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G475), .ZN(new_n536));
  XNOR2_X1  g350(.A(G113), .B(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n333), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n280), .A2(G143), .A3(G214), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(G143), .B1(new_n280), .B2(G214), .ZN(new_n541));
  OAI21_X1  g355(.A(G131), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n543));
  INV_X1    g357(.A(G237), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n327), .A3(G214), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n229), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n243), .A3(new_n539), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n542), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G140), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G125), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n441), .A2(G140), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT75), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .A4(KEYINPUT16), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT16), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT75), .B1(new_n550), .B2(KEYINPUT16), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G146), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n227), .B(new_n553), .C1(new_n554), .C2(new_n555), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n546), .A2(new_n539), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(KEYINPUT17), .A3(G131), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n548), .A2(new_n557), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n550), .A2(new_n551), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n562), .B1(new_n563), .B2(G146), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT76), .A4(new_n227), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(G146), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(KEYINPUT18), .A2(G131), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n546), .A2(new_n539), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n559), .A2(KEYINPUT18), .A3(G131), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n538), .B1(new_n561), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n561), .A2(new_n538), .A3(new_n572), .ZN(new_n575));
  AOI21_X1  g389(.A(G902), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n536), .B1(new_n576), .B2(KEYINPUT92), .ZN(new_n577));
  INV_X1    g391(.A(new_n575), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n323), .B1(new_n578), .B2(new_n573), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT92), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n542), .A2(new_n547), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n563), .B(KEYINPUT19), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n557), .B(new_n582), .C1(new_n583), .C2(G146), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n538), .B1(new_n584), .B2(new_n572), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(G475), .A2(G902), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT20), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT20), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n590), .B(new_n587), .C1(new_n578), .C2(new_n585), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n577), .A2(new_n581), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n529), .A2(new_n530), .A3(new_n323), .A4(new_n533), .ZN(new_n593));
  INV_X1    g407(.A(G952), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(G953), .ZN(new_n595));
  INV_X1    g409(.A(G234), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n595), .B1(new_n596), .B2(new_n544), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI211_X1 g412(.A(new_n323), .B(new_n327), .C1(G234), .C2(G237), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT21), .B(G898), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n535), .A2(new_n592), .A3(new_n593), .A4(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n478), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n518), .B1(G234), .B2(new_n323), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT24), .B(G110), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n250), .A2(G119), .ZN(new_n607));
  INV_X1    g421(.A(G119), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G128), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n607), .A2(new_n609), .A3(KEYINPUT72), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT72), .B1(new_n607), .B2(new_n609), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G110), .ZN(new_n613));
  NAND2_X1  g427(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n614), .ZN(new_n616));
  NOR2_X1   g430(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(G119), .B(G128), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n613), .B(new_n615), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n557), .A2(new_n621), .A3(new_n566), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT22), .B(G137), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n327), .A2(G221), .A3(G234), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OR3_X1    g439(.A1(new_n610), .A2(new_n611), .A3(new_n606), .ZN(new_n626));
  INV_X1    g440(.A(new_n558), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT16), .ZN(new_n628));
  OR3_X1    g442(.A1(new_n441), .A2(KEYINPUT16), .A3(G140), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(KEYINPUT75), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n227), .B1(new_n630), .B2(new_n553), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n626), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n607), .A2(new_n609), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT73), .B(KEYINPUT23), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n633), .A2(new_n634), .B1(new_n607), .B2(new_n614), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n635), .A2(KEYINPUT74), .A3(new_n613), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT74), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n638), .B2(G110), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n622), .B(new_n625), .C1(new_n632), .C2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n557), .A2(new_n558), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT74), .B1(new_n635), .B2(new_n613), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n638), .A2(new_n637), .A3(G110), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n643), .A2(new_n646), .A3(new_n626), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n625), .B1(new_n647), .B2(new_n622), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT25), .B1(new_n649), .B2(new_n323), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT25), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n642), .A2(new_n648), .A3(new_n651), .A4(G902), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n605), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n605), .A2(G902), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n649), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n319), .A2(new_n417), .A3(new_n604), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n348), .A2(new_n349), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G3));
  AOI21_X1  g473(.A(G902), .B1(new_n286), .B2(new_n297), .ZN(new_n660));
  INV_X1    g474(.A(G472), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT100), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n298), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n664), .B(G472), .C1(new_n317), .C2(G902), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n417), .A3(new_n656), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n323), .A2(G478), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n520), .B1(new_n525), .B2(KEYINPUT102), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n509), .A2(new_n670), .A3(new_n517), .A4(new_n519), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT33), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT33), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n524), .A2(new_n527), .A3(new_n674), .A4(new_n528), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n668), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(G478), .B1(new_n529), .B2(new_n323), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n577), .A2(new_n581), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n589), .A2(new_n591), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n471), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(KEYINPUT101), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n451), .B2(new_n469), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n471), .B(KEYINPUT101), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n451), .A2(new_n469), .A3(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n687), .A2(new_n477), .A3(new_n602), .A4(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n667), .A2(new_n682), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT34), .B(G104), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G6));
  NAND2_X1  g507(.A1(new_n679), .A2(KEYINPUT103), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n577), .A2(new_n695), .A3(new_n581), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n694), .A2(new_n696), .B1(new_n589), .B2(new_n591), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n535), .A2(new_n593), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n667), .A2(new_n690), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT35), .B(G107), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G9));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n647), .A2(new_n703), .A3(new_n622), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n703), .B1(new_n647), .B2(new_n622), .ZN(new_n706));
  INV_X1    g520(.A(new_n625), .ZN(new_n707));
  OAI22_X1  g521(.A1(new_n705), .A2(new_n706), .B1(KEYINPUT36), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n647), .A2(new_n622), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT104), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n707), .A2(KEYINPUT36), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n704), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n708), .A2(new_n655), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT105), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n708), .A2(new_n712), .A3(new_n715), .A4(new_n655), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n653), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT106), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n653), .A2(new_n714), .A3(new_n719), .A4(new_n716), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n666), .A2(new_n417), .A3(new_n604), .A4(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT37), .B(G110), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G12));
  AND3_X1   g538(.A1(new_n451), .A2(new_n469), .A3(new_n688), .ZN(new_n725));
  INV_X1    g539(.A(new_n477), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n725), .A2(new_n686), .A3(new_n726), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n718), .A2(new_n727), .A3(new_n720), .ZN(new_n728));
  INV_X1    g542(.A(G900), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n599), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n597), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n697), .A2(new_n698), .A3(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n319), .A2(new_n728), .A3(new_n732), .A4(new_n417), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G128), .ZN(G30));
  XNOR2_X1  g548(.A(new_n731), .B(KEYINPUT39), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n417), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT40), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT38), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n476), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT38), .B1(new_n473), .B2(new_n475), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n717), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n592), .B1(new_n535), .B2(new_n593), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n477), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n309), .A2(new_n284), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(G902), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n300), .A2(new_n284), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n661), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n298), .B2(KEYINPUT32), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n299), .A2(new_n752), .A3(new_n318), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n747), .A2(KEYINPUT107), .A3(new_n753), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n739), .A2(new_n740), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G143), .ZN(G45));
  OAI211_X1 g573(.A(new_n681), .B(new_n731), .C1(new_n676), .C2(new_n677), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n319), .A2(new_n728), .A3(new_n417), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G146), .ZN(G48));
  AND3_X1   g577(.A1(new_n409), .A2(new_n410), .A3(new_n323), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n410), .B1(new_n409), .B2(new_n323), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n764), .A2(new_n765), .A3(new_n324), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n682), .A2(new_n690), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n319), .A2(new_n766), .A3(new_n656), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT41), .B(G113), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G15));
  NOR2_X1   g584(.A1(new_n699), .A2(new_n690), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n319), .A3(new_n766), .A4(new_n656), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G116), .ZN(G18));
  NAND3_X1  g587(.A1(new_n718), .A2(new_n727), .A3(new_n720), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n603), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n319), .A3(new_n766), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT109), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(new_n778), .A3(new_n319), .A4(new_n766), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G119), .ZN(G21));
  OAI21_X1  g595(.A(G472), .B1(new_n317), .B2(G902), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT31), .B1(new_n287), .B2(new_n291), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n294), .A2(new_n295), .A3(new_n293), .ZN(new_n784));
  OAI22_X1  g598(.A1(new_n783), .A2(new_n784), .B1(new_n310), .B2(new_n284), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n188), .B(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n656), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n727), .A2(new_n602), .A3(new_n746), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n766), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G122), .ZN(G24));
  OAI211_X1 g605(.A(new_n787), .B(new_n717), .C1(new_n660), .C2(new_n661), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n760), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n766), .A3(new_n727), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G125), .ZN(G27));
  INV_X1    g609(.A(new_n324), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n473), .A2(new_n796), .A3(new_n477), .A4(new_n475), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n411), .B2(new_n416), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n761), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n316), .B1(new_n317), .B2(new_n189), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n314), .A2(new_n315), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n656), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT42), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n760), .A2(KEYINPUT42), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n319), .A2(new_n798), .A3(new_n656), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(KEYINPUT111), .B(G131), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G33));
  NAND4_X1  g622(.A1(new_n319), .A2(new_n732), .A3(new_n656), .A4(new_n798), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G134), .ZN(G36));
  NOR2_X1   g624(.A1(new_n666), .A2(new_n745), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n592), .B(KEYINPUT43), .C1(new_n676), .C2(new_n677), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n592), .B1(new_n676), .B2(new_n677), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT43), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n816), .A2(KEYINPUT112), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT112), .B1(new_n816), .B2(new_n817), .ZN(new_n819));
  OAI22_X1  g633(.A1(new_n814), .A2(new_n815), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT44), .B1(new_n811), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n410), .B1(new_n415), .B2(KEYINPUT45), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT45), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n413), .A2(new_n414), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n412), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n411), .B1(new_n825), .B2(KEYINPUT46), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT46), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n827), .B(new_n412), .C1(new_n822), .C2(new_n824), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n796), .B(new_n735), .C1(new_n826), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n821), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n811), .A2(KEYINPUT44), .A3(new_n820), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n473), .A2(new_n477), .A3(new_n475), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(KEYINPUT114), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT114), .B1(new_n831), .B2(new_n833), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(new_n215), .ZN(G39));
  OAI21_X1  g652(.A(new_n796), .B1(new_n826), .B2(new_n828), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT47), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(KEYINPUT47), .B(new_n796), .C1(new_n826), .C2(new_n828), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n319), .A2(new_n656), .A3(new_n760), .A4(new_n832), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(G140), .ZN(G42));
  NOR4_X1   g660(.A1(new_n744), .A2(new_n325), .A3(new_n726), .A4(new_n816), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n764), .A2(new_n765), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(KEYINPUT49), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n299), .A2(new_n752), .A3(new_n656), .A4(new_n318), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(KEYINPUT49), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n847), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n299), .A2(new_n752), .A3(new_n318), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n411), .A2(new_n416), .ZN(new_n857));
  INV_X1    g671(.A(new_n731), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n324), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n653), .A2(new_n714), .A3(new_n716), .A4(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n857), .A2(new_n727), .A3(new_n746), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n855), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n727), .A2(new_n860), .A3(new_n746), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n753), .A2(new_n863), .A3(KEYINPUT115), .A4(new_n857), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n774), .A2(new_n699), .A3(new_n858), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n774), .A2(new_n760), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n319), .B(new_n417), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(KEYINPUT52), .A2(new_n865), .A3(new_n794), .A4(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n733), .A2(new_n762), .A3(new_n794), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT52), .B1(new_n870), .B2(new_n865), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n696), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n695), .B1(new_n577), .B2(new_n581), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n680), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n535), .A2(new_n593), .A3(new_n731), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n875), .A2(new_n832), .A3(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n319), .A2(new_n417), .A3(new_n877), .A4(new_n721), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n793), .A2(new_n798), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n809), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n806), .A2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n772), .A2(new_n768), .A3(new_n790), .ZN(new_n882));
  INV_X1    g696(.A(new_n475), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n474), .B1(new_n451), .B2(new_n469), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n477), .B(new_n602), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n698), .A2(new_n592), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n682), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n666), .A2(new_n887), .A3(new_n417), .A4(new_n656), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n888), .A2(new_n722), .A3(new_n657), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n881), .A2(new_n780), .A3(new_n882), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n854), .B1(new_n872), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n809), .A2(new_n878), .A3(new_n879), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n889), .A2(new_n893), .A3(new_n803), .A4(new_n805), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n780), .A2(new_n882), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT52), .ZN(new_n897));
  INV_X1    g711(.A(new_n865), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n733), .A2(new_n762), .A3(new_n794), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n870), .A2(KEYINPUT52), .A3(new_n865), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n896), .A2(new_n902), .A3(KEYINPUT53), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n891), .A2(new_n892), .A3(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(KEYINPUT116), .B(new_n854), .C1(new_n872), .C2(new_n890), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(KEYINPUT54), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n891), .A2(new_n907), .A3(new_n903), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT51), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n818), .A2(new_n819), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n812), .B(KEYINPUT113), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n598), .B(new_n788), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n832), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n848), .A2(new_n325), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT117), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n843), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT117), .B1(new_n841), .B2(new_n842), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT118), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n920), .B(new_n913), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT50), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n726), .B1(new_n742), .B2(new_n743), .ZN(new_n924));
  INV_X1    g738(.A(new_n765), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n796), .A3(new_n411), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n923), .B1(new_n912), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n816), .A2(new_n817), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT112), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n816), .A2(KEYINPUT112), .A3(new_n817), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n812), .B(new_n813), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n597), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n924), .A2(new_n926), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n935), .A2(KEYINPUT50), .A3(new_n936), .A4(new_n788), .ZN(new_n937));
  NOR4_X1   g751(.A1(new_n764), .A2(new_n765), .A3(new_n832), .A4(new_n324), .ZN(new_n938));
  INV_X1    g752(.A(new_n792), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n820), .A2(new_n598), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT119), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n935), .A2(KEYINPUT119), .A3(new_n939), .A4(new_n938), .ZN(new_n943));
  AOI22_X1  g757(.A1(new_n928), .A2(new_n937), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n678), .A2(new_n681), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n851), .A2(new_n938), .A3(new_n598), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT120), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n926), .A2(new_n597), .A3(new_n832), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n949), .A3(new_n851), .A4(new_n945), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT121), .B1(new_n944), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n928), .A2(new_n937), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n942), .A2(new_n943), .ZN(new_n954));
  AND4_X1   g768(.A1(KEYINPUT121), .A2(new_n953), .A3(new_n951), .A4(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n909), .B1(new_n922), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n935), .A2(new_n938), .ZN(new_n958));
  INV_X1    g772(.A(new_n802), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT48), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT48), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n958), .A2(new_n962), .A3(new_n959), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n935), .A2(new_n727), .A3(new_n766), .A4(new_n788), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n948), .A2(new_n681), .A3(new_n678), .A4(new_n851), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n964), .A2(new_n595), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n841), .A2(new_n842), .A3(new_n914), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n909), .B1(new_n968), .B2(new_n913), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n944), .A2(new_n951), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT122), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n944), .A2(new_n969), .A3(KEYINPUT122), .A4(new_n951), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n906), .A2(new_n908), .A3(new_n957), .A4(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT123), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n594), .A2(new_n327), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n975), .B2(new_n976), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n853), .B1(new_n977), .B2(new_n979), .ZN(G75));
  NOR2_X1   g794(.A1(new_n327), .A2(G952), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT56), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n891), .A2(new_n903), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(G902), .ZN(new_n985));
  INV_X1    g799(.A(G210), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n437), .A2(new_n450), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n447), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT55), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n982), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n987), .A2(new_n991), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT124), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n987), .A2(KEYINPUT124), .A3(new_n991), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G51));
  XNOR2_X1  g811(.A(new_n412), .B(KEYINPUT57), .ZN(new_n998));
  INV_X1    g812(.A(new_n908), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n907), .B1(new_n891), .B2(new_n903), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n409), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n984), .A2(G902), .A3(new_n824), .A4(new_n822), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n981), .B1(new_n1002), .B2(new_n1003), .ZN(G54));
  NAND2_X1  g818(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n586), .B1(new_n985), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n982), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n985), .A2(new_n586), .A3(new_n1005), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(G60));
  AND2_X1   g823(.A1(new_n673), .A2(new_n675), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G478), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT59), .Z(new_n1012));
  NOR2_X1   g826(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n999), .B2(new_n1000), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n982), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n906), .A2(new_n908), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1012), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1015), .B1(new_n1010), .B2(new_n1018), .ZN(G63));
  NAND2_X1  g833(.A1(G217), .A2(G902), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT125), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT60), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n984), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n649), .B(KEYINPUT126), .Z(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n708), .A2(new_n712), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n1025), .B(new_n982), .C1(new_n1026), .C2(new_n1023), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT61), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(G66));
  INV_X1    g843(.A(new_n600), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n327), .B1(new_n1030), .B2(new_n444), .ZN(new_n1031));
  INV_X1    g845(.A(new_n895), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(new_n889), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1031), .B1(new_n1033), .B2(new_n327), .ZN(new_n1034));
  INV_X1    g848(.A(G898), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n988), .B1(new_n1035), .B2(G953), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1034), .B(new_n1036), .ZN(G69));
  AOI21_X1  g851(.A(new_n837), .B1(new_n843), .B2(new_n844), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n959), .A2(new_n727), .A3(new_n746), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n870), .B1(new_n829), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n809), .ZN(new_n1041));
  NOR3_X1   g855(.A1(new_n1040), .A2(new_n806), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1038), .A2(new_n327), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n289), .A2(new_n290), .ZN(new_n1044));
  XNOR2_X1  g858(.A(new_n1044), .B(new_n583), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n1043), .B(new_n1045), .C1(new_n729), .C2(new_n327), .ZN(new_n1046));
  INV_X1    g860(.A(new_n736), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n832), .B1(new_n682), .B2(new_n886), .ZN(new_n1048));
  NAND4_X1  g862(.A1(new_n1047), .A2(new_n319), .A3(new_n656), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1038), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n758), .A2(new_n870), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT62), .ZN(new_n1053));
  XNOR2_X1  g867(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  AOI21_X1  g868(.A(G953), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1046), .B1(new_n1055), .B2(new_n1045), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n327), .B1(G227), .B2(G900), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1057), .ZN(new_n1059));
  OAI211_X1 g873(.A(new_n1046), .B(new_n1059), .C1(new_n1055), .C2(new_n1045), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1058), .A2(new_n1060), .ZN(G72));
  INV_X1    g875(.A(new_n750), .ZN(new_n1062));
  XNOR2_X1  g876(.A(new_n1052), .B(KEYINPUT62), .ZN(new_n1063));
  NOR3_X1   g877(.A1(new_n1063), .A2(new_n1050), .A3(new_n1033), .ZN(new_n1064));
  NAND2_X1  g878(.A1(G472), .A2(G902), .ZN(new_n1065));
  XOR2_X1   g879(.A(new_n1065), .B(KEYINPUT63), .Z(new_n1066));
  INV_X1    g880(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g881(.A(new_n1062), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g882(.A(new_n1033), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n1038), .A2(new_n1069), .A3(new_n1042), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1070), .A2(new_n1066), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1071), .A2(KEYINPUT127), .ZN(new_n1072));
  INV_X1    g886(.A(KEYINPUT127), .ZN(new_n1073));
  NAND3_X1  g887(.A1(new_n1070), .A2(new_n1073), .A3(new_n1066), .ZN(new_n1074));
  NOR2_X1   g888(.A1(new_n300), .A2(new_n284), .ZN(new_n1075));
  NAND3_X1  g889(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g890(.A1(new_n303), .A2(new_n306), .ZN(new_n1077));
  NOR2_X1   g891(.A1(new_n294), .A2(new_n295), .ZN(new_n1078));
  OR2_X1    g892(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g893(.A1(new_n904), .A2(new_n905), .A3(new_n1066), .A4(new_n1079), .ZN(new_n1080));
  AND4_X1   g894(.A1(new_n982), .A2(new_n1068), .A3(new_n1076), .A4(new_n1080), .ZN(G57));
endmodule


