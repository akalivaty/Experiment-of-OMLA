//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940;
  OAI21_X1  g000(.A(KEYINPUT91), .B1(G71gat), .B2(G78gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G71gat), .B(G78gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n207), .B(KEYINPUT92), .Z(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(new_n208), .ZN(new_n211));
  XNOR2_X1  g010(.A(G15gat), .B(G22gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT90), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G1gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT16), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n218), .B1(new_n215), .B2(new_n214), .ZN(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  MUX2_X1   g020(.A(new_n211), .B(new_n209), .S(new_n221), .Z(new_n222));
  NAND2_X1  g021(.A1(G231gat), .A2(G233gat), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(G211gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n222), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G127gat), .B(G155gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n230), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G232gat), .A2(G233gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(KEYINPUT41), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT93), .ZN(new_n237));
  XNOR2_X1  g036(.A(G134gat), .B(G162gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT14), .ZN(new_n241));
  INV_X1    g040(.A(G29gat), .ZN(new_n242));
  INV_X1    g041(.A(G36gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n244), .A2(new_n245), .B1(G29gat), .B2(G36gat), .ZN(new_n246));
  AND2_X1   g045(.A1(G43gat), .A2(G50gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(G43gat), .A2(G50gat), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT15), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT88), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n247), .A2(KEYINPUT15), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT89), .B(G50gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(G43gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n246), .A3(new_n249), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT17), .ZN(new_n257));
  NAND2_X1  g056(.A1(G99gat), .A2(G106gat), .ZN(new_n258));
  INV_X1    g057(.A(G85gat), .ZN(new_n259));
  INV_X1    g058(.A(G92gat), .ZN(new_n260));
  AOI22_X1  g059(.A1(KEYINPUT8), .A2(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT96), .ZN(new_n262));
  NAND2_X1  g061(.A1(G85gat), .A2(G92gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(KEYINPUT95), .B2(KEYINPUT7), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT94), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT7), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT95), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n264), .A2(new_n268), .B1(new_n263), .B2(new_n266), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G99gat), .B(G106gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT97), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G190gat), .B(G218gat), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n276), .B(KEYINPUT98), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n272), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n279), .A2(new_n256), .B1(KEYINPUT41), .B2(new_n235), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n275), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n278), .B1(new_n275), .B2(new_n280), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n240), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n280), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n277), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n275), .A2(new_n278), .A3(new_n280), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n239), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n233), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT99), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G113gat), .B(G141gat), .ZN(new_n292));
  INV_X1    g091(.A(G197gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT11), .B(G169gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT12), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n219), .B(G8gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n257), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G229gat), .A2(G233gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n221), .A2(new_n256), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT18), .ZN(new_n303));
  INV_X1    g102(.A(new_n256), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n300), .B(KEYINPUT13), .Z(new_n307));
  AOI22_X1  g106(.A1(new_n302), .A2(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n299), .A2(new_n301), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(KEYINPUT18), .A3(new_n300), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n297), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n310), .A3(new_n297), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G230gat), .ZN(new_n315));
  INV_X1    g114(.A(G233gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n262), .A2(new_n271), .A3(new_n269), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT100), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n207), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n272), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT10), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n210), .A2(new_n272), .A3(new_n322), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n317), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n317), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT101), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G120gat), .B(G148gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G176gat), .B(G204gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  OR3_X1    g131(.A1(new_n321), .A2(KEYINPUT101), .A3(new_n327), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n329), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n332), .B1(new_n329), .B2(new_n333), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n291), .A2(new_n314), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT32), .ZN(new_n338));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  INV_X1    g138(.A(G169gat), .ZN(new_n340));
  INV_X1    g139(.A(G176gat), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT26), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT26), .B1(new_n340), .B2(new_n341), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n345));
  NOR2_X1   g144(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT27), .B(G183gat), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n345), .ZN(new_n354));
  NAND2_X1  g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n344), .A2(new_n350), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n224), .A2(new_n349), .A3(KEYINPUT65), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT65), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(G183gat), .B2(G190gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n362));
  AND4_X1   g161(.A1(new_n358), .A2(new_n359), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT23), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(G169gat), .B2(G176gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n366), .A3(new_n339), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT25), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n224), .A2(new_n349), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n358), .A2(new_n362), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT64), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n364), .A2(new_n366), .A3(new_n339), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n358), .A2(new_n369), .A3(KEYINPUT64), .A4(new_n362), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n356), .A2(new_n368), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G134gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G127gat), .ZN(new_n379));
  INV_X1    g178(.A(G127gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G134gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G113gat), .B(G120gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT67), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n384), .A2(KEYINPUT1), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G120gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G113gat), .ZN(new_n388));
  INV_X1    g187(.A(G113gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G120gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G127gat), .B(G134gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n384), .A2(KEYINPUT1), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n377), .B(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n338), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(G15gat), .B(G43gat), .Z(new_n399));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT33), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT68), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n396), .A2(new_n397), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n405), .B(KEYINPUT34), .Z(new_n406));
  INV_X1    g205(.A(new_n398), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n396), .A2(new_n397), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n410), .A3(new_n401), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n404), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n403), .A2(KEYINPUT68), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT68), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n414), .B1(new_n398), .B2(new_n402), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n411), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n405), .B(KEYINPUT34), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT84), .ZN(new_n420));
  AND2_X1   g219(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n422));
  OAI21_X1  g221(.A(G148gat), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G141gat), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT76), .B1(new_n424), .B2(G148gat), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT76), .ZN(new_n426));
  INV_X1    g225(.A(G148gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(G141gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G155gat), .A2(G162gat), .ZN(new_n430));
  INV_X1    g229(.A(G155gat), .ZN(new_n431));
  INV_X1    g230(.A(G162gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n430), .B1(new_n433), .B2(KEYINPUT2), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n433), .A2(new_n430), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT2), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n424), .A2(G148gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n427), .A2(G141gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n429), .A2(new_n434), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G197gat), .B(G204gat), .ZN(new_n441));
  INV_X1    g240(.A(G211gat), .ZN(new_n442));
  INV_X1    g241(.A(G218gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n441), .B1(KEYINPUT22), .B2(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(G211gat), .B(G218gat), .Z(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(KEYINPUT77), .B(KEYINPUT3), .Z(new_n450));
  AOI21_X1  g249(.A(new_n440), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OR2_X1    g250(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n427), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n425), .A2(new_n428), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n434), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n435), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n450), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n447), .B1(new_n448), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n420), .B1(new_n451), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT3), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n456), .B2(new_n457), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(new_n419), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT29), .B1(new_n440), .B2(new_n450), .ZN(new_n464));
  OAI221_X1 g263(.A(new_n463), .B1(new_n464), .B2(new_n447), .C1(new_n440), .C2(new_n449), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(G78gat), .B(G106gat), .Z(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT83), .B(G50gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G22gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n466), .A2(new_n471), .ZN(new_n476));
  INV_X1    g275(.A(G22gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n472), .B2(new_n473), .ZN(new_n480));
  AOI211_X1 g279(.A(KEYINPUT85), .B(G22gat), .C1(new_n466), .C2(new_n471), .ZN(new_n481));
  OAI22_X1  g280(.A1(new_n480), .A2(new_n481), .B1(new_n471), .B2(new_n466), .ZN(new_n482));
  AND4_X1   g281(.A1(new_n412), .A2(new_n418), .A3(new_n479), .A4(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G225gat), .A2(G233gat), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n386), .A2(new_n394), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n440), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n440), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT78), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n486), .B1(new_n440), .B2(new_n450), .ZN(new_n493));
  INV_X1    g292(.A(new_n462), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n458), .A2(new_n395), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n496), .A2(KEYINPUT78), .A3(new_n462), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n485), .B(new_n491), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G1gat), .B(G29gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(new_n259), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT0), .B(G57gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n502), .B(new_n503), .Z(new_n504));
  NAND3_X1  g303(.A1(new_n493), .A2(new_n492), .A3(new_n494), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT78), .B1(new_n496), .B2(new_n462), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n507), .A2(KEYINPUT5), .A3(new_n485), .A4(new_n491), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n487), .A2(KEYINPUT79), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n456), .A2(new_n457), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n395), .ZN(new_n511));
  INV_X1    g310(.A(new_n485), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n395), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n487), .A2(new_n513), .A3(KEYINPUT79), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n500), .A2(new_n504), .A3(new_n508), .A4(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n509), .B(new_n513), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n498), .A2(new_n499), .B1(new_n520), .B2(new_n512), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n504), .B1(new_n521), .B2(new_n508), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n516), .A2(new_n518), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n484), .A2(KEYINPUT35), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n527));
  NAND2_X1  g326(.A1(G226gat), .A2(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT69), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n377), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n377), .A2(KEYINPUT71), .A3(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT70), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n377), .A2(new_n448), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(new_n528), .ZN(new_n538));
  INV_X1    g337(.A(new_n528), .ZN(new_n539));
  AOI211_X1 g338(.A(KEYINPUT70), .B(new_n539), .C1(new_n377), .C2(new_n448), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n535), .B(new_n447), .C1(new_n538), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT72), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n539), .B1(new_n377), .B2(new_n448), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(new_n536), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n447), .A4(new_n535), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n537), .A2(new_n529), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n377), .A2(new_n539), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n447), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n542), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G8gat), .B(G36gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G64gat), .B(G92gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n549), .B1(new_n541), .B2(KEYINPUT72), .ZN(new_n556));
  INV_X1    g355(.A(new_n554), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n556), .A2(KEYINPUT30), .A3(new_n546), .A4(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n527), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n558), .A2(new_n527), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n551), .A2(new_n554), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(KEYINPUT30), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n526), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n524), .B1(new_n523), .B2(KEYINPUT81), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT81), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n519), .B2(new_n522), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n563), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  AND4_X1   g370(.A1(KEYINPUT30), .A2(new_n556), .A3(new_n546), .A4(new_n557), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n557), .B1(new_n556), .B2(new_n546), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT73), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n527), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT74), .B1(new_n559), .B2(new_n560), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n571), .A2(new_n577), .A3(new_n483), .A4(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT87), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT35), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n579), .B2(KEYINPUT35), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n567), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n479), .A2(new_n482), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT86), .Z(new_n585));
  AND2_X1   g384(.A1(new_n571), .A2(new_n577), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n585), .B1(new_n586), .B2(new_n578), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n412), .A2(new_n418), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT36), .Z(new_n589));
  OR2_X1    g388(.A1(new_n520), .A2(new_n512), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n507), .A2(new_n491), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n590), .B(KEYINPUT39), .C1(new_n485), .C2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n504), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n591), .A2(KEYINPUT39), .A3(new_n485), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT40), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n516), .ZN(new_n599));
  AOI211_X1 g398(.A(new_n597), .B(new_n599), .C1(new_n561), .C2(new_n564), .ZN(new_n600));
  INV_X1    g399(.A(new_n584), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT37), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n556), .A2(new_n602), .A3(new_n546), .ZN(new_n603));
  INV_X1    g402(.A(new_n447), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n544), .A2(new_n604), .A3(new_n535), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n547), .A2(new_n548), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n602), .B1(new_n606), .B2(new_n447), .ZN(new_n607));
  AOI211_X1 g406(.A(KEYINPUT38), .B(new_n557), .C1(new_n605), .C2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n562), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n525), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n603), .A2(new_n554), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n551), .A2(KEYINPUT37), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n601), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n589), .B1(new_n600), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n587), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n337), .B1(new_n583), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n568), .A2(new_n570), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g422(.A(KEYINPUT16), .B(G8gat), .Z(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n565), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(KEYINPUT42), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT42), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n619), .A2(new_n565), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n628), .B2(G8gat), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n626), .B1(new_n625), .B2(new_n629), .ZN(G1325gat));
  INV_X1    g429(.A(new_n588), .ZN(new_n631));
  AOI21_X1  g430(.A(G15gat), .B1(new_n619), .B2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n589), .B(KEYINPUT102), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n634), .A2(G15gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n619), .B2(new_n635), .ZN(G1326gat));
  INV_X1    g435(.A(new_n585), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n619), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT43), .B(G22gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(G1327gat));
  INV_X1    g439(.A(new_n288), .ZN(new_n641));
  NOR4_X1   g440(.A1(new_n484), .A2(new_n565), .A3(KEYINPUT35), .A4(new_n525), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n579), .A2(KEYINPUT35), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT87), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT35), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n641), .B1(new_n646), .B2(new_n617), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n336), .ZN(new_n649));
  INV_X1    g448(.A(new_n314), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n649), .A2(new_n650), .A3(new_n233), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n652), .A2(G29gat), .A3(new_n620), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT45), .Z(new_n654));
  NAND2_X1  g453(.A1(new_n647), .A2(KEYINPUT44), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n583), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(KEYINPUT105), .B(new_n567), .C1(new_n581), .C2(new_n582), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n617), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n283), .A2(new_n287), .A3(KEYINPUT106), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT106), .B1(new_n283), .B2(new_n287), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n655), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n233), .B(KEYINPUT104), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n312), .A2(new_n667), .A3(new_n313), .ZN(new_n668));
  INV_X1    g467(.A(new_n313), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT103), .B1(new_n669), .B2(new_n311), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n666), .A2(new_n649), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G29gat), .B1(new_n673), .B2(new_n620), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n654), .A2(new_n674), .ZN(G1328gat));
  NOR3_X1   g474(.A1(new_n652), .A2(G36gat), .A3(new_n566), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT46), .ZN(new_n677));
  OAI21_X1  g476(.A(G36gat), .B1(new_n673), .B2(new_n566), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1329gat));
  NOR2_X1   g478(.A1(new_n588), .A2(G43gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n648), .A2(new_n651), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT108), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT47), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G43gat), .B1(new_n673), .B2(new_n589), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n664), .A2(new_n634), .A3(new_n672), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n687), .A2(new_n688), .A3(G43gat), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n687), .B2(G43gat), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n689), .A2(new_n690), .A3(new_n682), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n686), .B1(new_n691), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g491(.A1(new_n652), .A2(new_n585), .A3(new_n253), .ZN(new_n693));
  INV_X1    g492(.A(new_n673), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n637), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n695), .B2(new_n253), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n697));
  INV_X1    g496(.A(new_n253), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n694), .B2(new_n584), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT48), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  OAI22_X1  g500(.A1(new_n696), .A2(new_n697), .B1(new_n699), .B2(new_n701), .ZN(G1331gat));
  NAND3_X1  g501(.A1(new_n291), .A2(new_n649), .A3(new_n671), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n659), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n621), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g505(.A1(new_n659), .A2(new_n566), .A3(new_n703), .ZN(new_n707));
  NOR2_X1   g506(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n708));
  AND2_X1   g507(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(new_n707), .B2(new_n708), .ZN(G1333gat));
  NAND2_X1  g510(.A1(new_n704), .A2(new_n634), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n588), .A2(G71gat), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n712), .A2(G71gat), .B1(new_n704), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g514(.A1(new_n704), .A2(new_n637), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT110), .B(G78gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1335gat));
  NAND2_X1  g517(.A1(new_n668), .A2(new_n670), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n719), .A2(new_n336), .A3(new_n233), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n664), .A2(KEYINPUT111), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT111), .B1(new_n664), .B2(new_n720), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT112), .B1(new_n723), .B2(new_n621), .ZN(new_n724));
  OAI211_X1 g523(.A(KEYINPUT112), .B(new_n621), .C1(new_n721), .C2(new_n722), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G85gat), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n719), .A2(new_n233), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n641), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n659), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(KEYINPUT51), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n659), .A2(new_n731), .A3(new_n728), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n649), .A2(new_n259), .A3(new_n621), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT113), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n724), .A2(new_n726), .B1(new_n733), .B2(new_n735), .ZN(G1336gat));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n566), .A2(new_n336), .A3(G92gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n664), .A2(new_n720), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n740), .A2(new_n565), .ZN(new_n741));
  OAI221_X1 g540(.A(new_n737), .B1(new_n733), .B2(new_n739), .C1(new_n741), .C2(new_n260), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n646), .A2(KEYINPUT105), .ZN(new_n743));
  INV_X1    g542(.A(new_n658), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n618), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n728), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(KEYINPUT114), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n659), .B2(new_n728), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n749), .A3(new_n731), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT115), .ZN(new_n751));
  INV_X1    g550(.A(new_n732), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n747), .A2(new_n749), .A3(new_n753), .A4(new_n731), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n565), .B1(new_n721), .B2(new_n722), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n755), .A2(new_n738), .B1(new_n756), .B2(G92gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n742), .B1(new_n757), .B2(new_n737), .ZN(G1337gat));
  AND2_X1   g557(.A1(new_n723), .A2(new_n634), .ZN(new_n759));
  INV_X1    g558(.A(G99gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n649), .A2(new_n760), .A3(new_n631), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n759), .A2(new_n760), .B1(new_n733), .B2(new_n761), .ZN(G1338gat));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n637), .B1(new_n721), .B2(new_n722), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(G106gat), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n336), .A2(G106gat), .A3(new_n601), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n755), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n730), .B2(new_n732), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT116), .B1(new_n740), .B2(new_n584), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n664), .A2(KEYINPUT116), .A3(new_n584), .A4(new_n720), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G106gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n765), .A2(new_n767), .B1(new_n772), .B2(new_n763), .ZN(G1339gat));
  NOR2_X1   g572(.A1(new_n309), .A2(new_n300), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n306), .A2(new_n307), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n296), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n776), .A2(new_n313), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n334), .B2(new_n335), .ZN(new_n778));
  INV_X1    g577(.A(new_n326), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n323), .A2(new_n317), .A3(new_n325), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(KEYINPUT54), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n332), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n326), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT117), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  INV_X1    g587(.A(new_n335), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n781), .A2(new_n790), .A3(new_n784), .A4(KEYINPUT55), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n787), .A2(new_n788), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n778), .B1(new_n792), .B2(new_n671), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n662), .ZN(new_n794));
  INV_X1    g593(.A(new_n792), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n288), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n283), .A2(new_n287), .A3(KEYINPUT106), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n795), .A2(new_n799), .A3(new_n777), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n794), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n335), .B1(new_n786), .B2(new_n785), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n719), .A2(new_n803), .A3(new_n791), .A4(new_n787), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n799), .B1(new_n804), .B2(new_n778), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n803), .A2(new_n791), .A3(new_n787), .A4(new_n777), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n662), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT118), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n802), .A2(new_n808), .A3(new_n665), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n291), .A2(new_n336), .A3(new_n671), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n621), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n565), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n637), .A2(new_n588), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G113gat), .B1(new_n815), .B2(new_n650), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n812), .A2(new_n484), .A3(new_n565), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n389), .A3(new_n719), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1340gat));
  OAI21_X1  g618(.A(G120gat), .B1(new_n815), .B2(new_n336), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n649), .A2(new_n387), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT119), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(G1341gat));
  NOR3_X1   g623(.A1(new_n815), .A2(new_n380), .A3(new_n665), .ZN(new_n825));
  AOI21_X1  g624(.A(G127gat), .B1(new_n817), .B2(new_n233), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(G1342gat));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n484), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n288), .A2(new_n565), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n378), .A3(new_n829), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n830), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(KEYINPUT56), .ZN(new_n832));
  OAI21_X1  g631(.A(G134gat), .B1(new_n815), .B2(new_n288), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT120), .B1(new_n830), .B2(KEYINPUT56), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n834), .ZN(G1343gat));
  NAND2_X1  g634(.A1(new_n633), .A2(new_n584), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT121), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n813), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n650), .A2(G141gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n589), .A2(new_n621), .A3(new_n566), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n795), .A2(new_n314), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n641), .B1(new_n841), .B2(new_n778), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n233), .B1(new_n843), .B2(new_n800), .ZN(new_n844));
  INV_X1    g643(.A(new_n810), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n637), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n840), .B1(new_n846), .B2(KEYINPUT57), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n601), .B1(new_n809), .B2(new_n810), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n719), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n421), .A2(new_n422), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n838), .A2(new_n839), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854));
  INV_X1    g653(.A(new_n852), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n847), .A2(new_n850), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n314), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n813), .A2(new_n837), .A3(new_n839), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n854), .ZN(new_n859));
  OAI22_X1  g658(.A1(new_n853), .A2(new_n854), .B1(new_n857), .B2(new_n859), .ZN(G1344gat));
  NAND2_X1  g659(.A1(new_n427), .A2(KEYINPUT59), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n838), .B2(new_n649), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n649), .A3(new_n850), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n811), .A2(new_n584), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT57), .ZN(new_n867));
  INV_X1    g666(.A(new_n233), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n806), .A2(new_n288), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n842), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n291), .A2(new_n650), .A3(new_n336), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n585), .A2(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n840), .A2(new_n864), .A3(new_n336), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n867), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n865), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n862), .B1(new_n877), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g677(.A(G155gat), .B1(new_n838), .B2(new_n233), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n665), .A2(new_n431), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n856), .B2(new_n880), .ZN(G1346gat));
  AND2_X1   g680(.A1(new_n856), .A2(new_n799), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n837), .A2(new_n432), .A3(new_n829), .ZN(new_n883));
  OAI22_X1  g682(.A1(new_n882), .A2(new_n432), .B1(new_n812), .B2(new_n883), .ZN(G1347gat));
  NOR2_X1   g683(.A1(new_n566), .A2(new_n621), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n811), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n814), .ZN(new_n887));
  OAI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n650), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n811), .A2(new_n483), .A3(new_n885), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n340), .A3(new_n719), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1348gat));
  NAND4_X1  g690(.A1(new_n886), .A2(G176gat), .A3(new_n649), .A4(new_n814), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  AOI21_X1  g694(.A(G176gat), .B1(new_n889), .B2(new_n649), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G1349gat));
  OAI21_X1  g696(.A(G183gat), .B1(new_n887), .B2(new_n665), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n889), .A2(new_n348), .A3(new_n233), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT60), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(KEYINPUT60), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n898), .A2(new_n903), .A3(new_n899), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1350gat));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n349), .A3(new_n799), .ZN(new_n906));
  OAI21_X1  g705(.A(G190gat), .B1(new_n887), .B2(new_n288), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(G1351gat));
  AND2_X1   g709(.A1(new_n633), .A2(new_n885), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n848), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(new_n293), .A3(new_n719), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT124), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n874), .B(new_n911), .C1(new_n848), .C2(new_n849), .ZN(new_n915));
  OAI21_X1  g714(.A(G197gat), .B1(new_n915), .B2(new_n650), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1352gat));
  INV_X1    g716(.A(G204gat), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n915), .A2(new_n336), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(KEYINPUT125), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(KEYINPUT125), .B2(new_n919), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n912), .A2(new_n918), .A3(new_n649), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(G1353gat));
  OAI211_X1 g724(.A(KEYINPUT63), .B(G211gat), .C1(new_n915), .C2(new_n868), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n867), .A2(new_n233), .A3(new_n874), .A4(new_n911), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n929), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n930));
  OAI21_X1  g729(.A(G211gat), .B1(new_n915), .B2(new_n868), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n928), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n912), .A2(new_n442), .A3(new_n233), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT126), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1354gat));
  AND2_X1   g736(.A1(new_n912), .A2(new_n799), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n641), .A2(G218gat), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n938), .A2(G218gat), .B1(new_n915), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(G1355gat));
endmodule


