//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n588, new_n589,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n638, new_n641, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1209,
    new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(G2104), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR3_X1   g040(.A1(new_n465), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n467), .B2(G101), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(new_n466), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  NOR3_X1   g045(.A1(new_n469), .A2(KEYINPUT68), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G137), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n478), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n463), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n472), .A2(new_n480), .ZN(G160));
  AOI21_X1  g056(.A(new_n463), .B1(new_n474), .B2(new_n475), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT69), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n476), .A2(G136), .ZN(new_n488));
  NOR3_X1   g063(.A1(new_n484), .A2(new_n487), .A3(new_n488), .ZN(G162));
  AND2_X1   g064(.A1(KEYINPUT70), .A2(G114), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT70), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n482), .A2(G126), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n476), .B2(G138), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n496), .A2(new_n463), .A3(G138), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n478), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT71), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(KEYINPUT71), .A2(KEYINPUT6), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n503), .A2(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n507), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n504), .B2(new_n506), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT73), .A3(new_n512), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(G88), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n521), .B1(new_n520), .B2(new_n523), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(G75), .A2(G543), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n505), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT72), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n513), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G62), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(KEYINPUT75), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  NOR3_X1   g112(.A1(new_n524), .A2(new_n525), .A3(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT76), .B(G51), .Z(new_n542));
  NAND2_X1  g117(.A1(new_n522), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n516), .A2(G89), .A3(new_n519), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  AND3_X1   g123(.A1(new_n518), .A2(KEYINPUT73), .A3(new_n512), .ZN(new_n549));
  AOI21_X1  g124(.A(KEYINPUT73), .B1(new_n518), .B2(new_n512), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  NOR3_X1   g126(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n522), .A2(G52), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n554), .B2(new_n528), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(G171));
  NAND3_X1  g131(.A1(new_n516), .A2(G81), .A3(new_n519), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n518), .B2(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n558), .B1(new_n561), .B2(new_n528), .ZN(new_n562));
  OAI211_X1 g137(.A(G56), .B(new_n513), .C1(new_n531), .C2(new_n532), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(new_n559), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n564), .A2(KEYINPUT77), .A3(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n522), .A2(G43), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n557), .A2(new_n562), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  OAI211_X1 g148(.A(G65), .B(new_n513), .C1(new_n531), .C2(new_n532), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n522), .A2(new_n577), .A3(G53), .ZN(new_n578));
  AND3_X1   g153(.A1(KEYINPUT71), .A2(KEYINPUT6), .A3(G651), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT6), .B1(KEYINPUT71), .B2(G651), .ZN(new_n580));
  OAI211_X1 g155(.A(G53), .B(G543), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT9), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n576), .A2(G651), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n516), .A2(G91), .A3(new_n519), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  NAND2_X1  g162(.A1(new_n520), .A2(new_n523), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n529), .A2(new_n536), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G303));
  OAI21_X1  g167(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g170(.A(KEYINPUT78), .B(G651), .C1(new_n518), .C2(G74), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n516), .A2(G87), .A3(new_n519), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n522), .A2(G49), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G288));
  NOR2_X1   g175(.A1(new_n549), .A2(new_n550), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G86), .B1(G48), .B2(new_n522), .ZN(new_n602));
  OAI211_X1 g177(.A(G61), .B(new_n513), .C1(new_n531), .C2(new_n532), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(KEYINPUT79), .B1(G73), .B2(G543), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT79), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n518), .A2(new_n605), .A3(G61), .ZN(new_n606));
  AOI211_X1 g181(.A(KEYINPUT80), .B(new_n528), .C1(new_n604), .C2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(KEYINPUT79), .ZN(new_n609));
  NAND2_X1  g184(.A1(G73), .A2(G543), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n608), .B1(new_n611), .B2(G651), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n602), .B1(new_n607), .B2(new_n612), .ZN(G305));
  NAND2_X1  g188(.A1(G72), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G60), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n533), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G47), .B2(new_n522), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n516), .A2(G85), .A3(new_n519), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT81), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n516), .A2(G92), .A3(new_n519), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n516), .A2(KEYINPUT10), .A3(G92), .A4(new_n519), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT82), .B(G66), .Z(new_n627));
  AOI22_X1  g202(.A1(new_n518), .A2(new_n627), .B1(G79), .B2(G543), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n528), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n518), .A2(new_n627), .ZN(new_n631));
  AND2_X1   g206(.A1(G79), .A2(G543), .ZN(new_n632));
  OAI21_X1  g207(.A(KEYINPUT83), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n630), .A2(new_n633), .B1(G54), .B2(new_n522), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n621), .B1(G868), .B2(new_n635), .ZN(G284));
  OAI21_X1  g211(.A(new_n621), .B1(G868), .B2(new_n635), .ZN(G321));
  NAND2_X1  g212(.A1(G286), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n585), .B2(G868), .ZN(G297));
  OAI21_X1  g214(.A(new_n638), .B1(new_n585), .B2(G868), .ZN(G280));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n635), .B1(new_n641), .B2(G860), .ZN(G148));
  NAND2_X1  g217(.A1(new_n635), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G868), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g221(.A1(new_n467), .A2(new_n478), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT13), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n476), .A2(G135), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n482), .A2(G123), .ZN(new_n653));
  OR2_X1    g228(.A1(G99), .A2(G2105), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n654), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n656), .A2(G2096), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(G2096), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n657), .A3(new_n658), .ZN(G156));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n665), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  AND3_X1   g248(.A1(new_n672), .A2(new_n673), .A3(G14), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT85), .Z(G401));
  XNOR2_X1  g250(.A(G2084), .B(G2090), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2072), .B(G2078), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n679), .B(KEYINPUT17), .Z(new_n685));
  AOI21_X1  g260(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n684), .B1(new_n677), .B2(new_n685), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n678), .ZN(new_n688));
  XOR2_X1   g263(.A(G2096), .B(G2100), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT19), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT20), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n694), .A2(new_n695), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n693), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n693), .B2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1991), .B(G1996), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  NAND2_X1  g284(.A1(new_n478), .A2(G127), .ZN(new_n710));
  INV_X1    g285(.A(G115), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n465), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT94), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n463), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n713), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n718), .A2(new_n719), .B1(new_n476), .B2(G139), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n723), .B2(G33), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(G2072), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(G2072), .ZN(new_n728));
  NAND2_X1  g303(.A1(G160), .A2(G29), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G34), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n729), .B1(G29), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G2084), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT31), .B(G11), .Z(new_n735));
  NOR2_X1   g310(.A1(new_n656), .A2(new_n723), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT98), .B(G28), .Z(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT30), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n737), .B2(KEYINPUT30), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n735), .B(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n727), .A2(new_n728), .A3(new_n734), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n723), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n723), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT29), .ZN(new_n744));
  INV_X1    g319(.A(G16), .ZN(new_n745));
  NOR2_X1   g320(.A1(G286), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT97), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT97), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G16), .B2(G21), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n747), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n744), .A2(G2090), .B1(G1966), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G27), .A2(G29), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G164), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT100), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G2078), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n751), .B(new_n755), .C1(G2090), .C2(new_n744), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n723), .A2(G26), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT28), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n476), .A2(G140), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n482), .A2(G128), .ZN(new_n760));
  OR2_X1    g335(.A1(G104), .A2(G2105), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n758), .B1(new_n763), .B2(G29), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT92), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G2067), .Z(new_n766));
  AND2_X1   g341(.A1(new_n723), .A2(G32), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n476), .A2(G141), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n467), .A2(G105), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n482), .A2(G129), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AND4_X1   g348(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT96), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(KEYINPUT96), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n767), .B1(new_n777), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT27), .B(G1996), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G1961), .ZN(new_n781));
  NOR2_X1   g356(.A1(G171), .A2(new_n745), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G5), .B2(new_n745), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n766), .B(new_n780), .C1(new_n781), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n750), .A2(G1966), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n741), .A2(new_n756), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n732), .A2(new_n733), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n778), .B2(new_n779), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n781), .B2(new_n783), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT99), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n745), .A2(G4), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n635), .B2(new_n745), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT91), .B(G1348), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n745), .A2(G20), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT23), .Z(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G299), .B2(G16), .ZN(new_n797));
  INV_X1    g372(.A(G1956), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n568), .A2(new_n745), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n745), .B2(G19), .ZN(new_n801));
  INV_X1    g376(.A(G1341), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n801), .A2(new_n802), .B1(new_n754), .B2(G2078), .ZN(new_n803));
  AOI211_X1 g378(.A(new_n799), .B(new_n803), .C1(new_n802), .C2(new_n801), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n786), .A2(new_n790), .A3(new_n794), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n723), .A2(G25), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n476), .A2(G131), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n482), .A2(G119), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n463), .A2(G107), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT88), .Z(new_n812));
  OAI21_X1  g387(.A(new_n806), .B1(new_n812), .B2(new_n723), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n745), .A2(G24), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G290), .B2(G16), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(G1986), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n813), .A2(new_n815), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(G1986), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n816), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n745), .A2(G23), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(new_n745), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT33), .Z(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(G1976), .ZN(new_n828));
  NOR2_X1   g403(.A1(G16), .A2(G22), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G166), .B2(G16), .ZN(new_n830));
  INV_X1    g405(.A(G1971), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n827), .A2(G1976), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n828), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n745), .A2(G6), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n522), .A2(G48), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n516), .A2(new_n519), .ZN(new_n837));
  INV_X1    g412(.A(G86), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n611), .A2(G651), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT80), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n528), .B1(new_n604), .B2(new_n606), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n608), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n839), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n835), .B1(new_n844), .B2(new_n745), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT32), .B(G1981), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT90), .B1(new_n834), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G1976), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n827), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT90), .ZN(new_n851));
  INV_X1    g426(.A(new_n847), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n832), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n823), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n855), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n848), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT36), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n856), .A2(new_n861), .A3(new_n858), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n805), .B1(new_n860), .B2(new_n862), .ZN(G311));
  INV_X1    g438(.A(new_n805), .ZN(new_n864));
  INV_X1    g439(.A(new_n862), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n861), .B1(new_n856), .B2(new_n858), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(G150));
  NAND2_X1  g442(.A1(new_n635), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g444(.A1(G80), .A2(G543), .ZN(new_n870));
  INV_X1    g445(.A(G67), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n533), .B2(new_n871), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n872), .A2(G651), .B1(G55), .B2(new_n522), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n516), .A2(G93), .A3(new_n519), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n567), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n567), .A2(new_n875), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n869), .B(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n880), .A2(new_n881), .A3(G860), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n875), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n884));
  XOR2_X1   g459(.A(new_n883), .B(new_n884), .Z(new_n885));
  OR2_X1    g460(.A1(new_n882), .A2(new_n885), .ZN(G145));
  INV_X1    g461(.A(new_n763), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n775), .A2(new_n776), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n775), .B2(new_n776), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n649), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  INV_X1    g467(.A(new_n649), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n893), .A3(new_n888), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n500), .B(KEYINPUT102), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n896), .A2(new_n721), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n721), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n476), .A2(G142), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n482), .A2(G130), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n463), .A2(G118), .ZN(new_n901));
  OAI21_X1  g476(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n899), .B(new_n900), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n811), .B(new_n903), .Z(new_n904));
  AND3_X1   g479(.A1(new_n897), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n897), .B2(new_n898), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n895), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n891), .A2(new_n894), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n905), .B2(new_n906), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(G160), .B(new_n656), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(G162), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(KEYINPUT103), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n911), .A2(new_n913), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(G37), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g497(.A(new_n643), .B(new_n878), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n626), .A2(new_n585), .A3(new_n634), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n585), .B1(new_n626), .B2(new_n634), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n626), .A2(new_n634), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G299), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n626), .A2(new_n634), .A3(new_n585), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n923), .A2(new_n928), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n932), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n936), .B2(new_n923), .ZN(new_n937));
  XOR2_X1   g512(.A(new_n937), .B(KEYINPUT42), .Z(new_n938));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n617), .A2(new_n939), .A3(new_n618), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n617), .B2(new_n618), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n825), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(G290), .A2(KEYINPUT105), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n617), .A2(new_n939), .A3(new_n618), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(G288), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(G166), .A2(new_n844), .ZN(new_n947));
  NOR2_X1   g522(.A1(G303), .A2(G305), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G166), .A2(new_n844), .ZN(new_n950));
  NAND2_X1  g525(.A1(G303), .A2(G305), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n942), .A4(new_n945), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(KEYINPUT106), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n938), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n938), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n875), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(G868), .B2(new_n958), .ZN(G295));
  OAI21_X1  g534(.A(new_n957), .B1(G868), .B2(new_n958), .ZN(G331));
  NAND2_X1  g535(.A1(new_n928), .A2(new_n933), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n516), .A2(G90), .A3(new_n519), .ZN(new_n962));
  NAND2_X1  g537(.A1(G77), .A2(G543), .ZN(new_n963));
  INV_X1    g538(.A(G64), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n533), .B2(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n965), .A2(G651), .B1(G52), .B2(new_n522), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n516), .A2(G89), .A3(new_n519), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n962), .B(new_n966), .C1(new_n967), .C2(new_n544), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n546), .B(new_n545), .C1(new_n552), .C2(new_n555), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n876), .B2(new_n877), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n557), .A2(new_n562), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n565), .A2(new_n566), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n874), .A4(new_n873), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n567), .A2(new_n875), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n968), .A4(new_n969), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n961), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n971), .A2(new_n976), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n936), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n953), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G37), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n953), .B1(new_n978), .B2(new_n980), .ZN(new_n984));
  OR3_X1    g559(.A1(new_n983), .A2(KEYINPUT43), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n935), .B1(new_n976), .B2(new_n971), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT41), .B1(new_n926), .B2(new_n927), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n930), .A2(new_n932), .A3(new_n924), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n988), .B1(new_n977), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(new_n992), .B2(new_n953), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n977), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n980), .ZN(new_n995));
  INV_X1    g570(.A(new_n953), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(KEYINPUT109), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n983), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n985), .B(KEYINPUT44), .C1(new_n986), .C2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT43), .B1(new_n983), .B2(new_n984), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT108), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(KEYINPUT43), .C1(new_n983), .C2(new_n984), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n998), .A2(new_n1005), .A3(new_n986), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n981), .A2(new_n982), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n992), .A2(new_n987), .A3(new_n953), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT109), .B1(new_n995), .B2(new_n996), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n986), .B(new_n1007), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT110), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1004), .A2(new_n1006), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n1014));
  OAI21_X1  g589(.A(new_n999), .B1(new_n1013), .B2(new_n1014), .ZN(G397));
  INV_X1    g590(.A(G40), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n472), .A2(new_n1016), .A3(new_n480), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  INV_X1    g593(.A(G1384), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n500), .A2(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1996), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT111), .Z(new_n1024));
  INV_X1    g599(.A(new_n1021), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n763), .B(G2067), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n777), .B2(G1996), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1024), .A2(new_n777), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n811), .B(new_n815), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n1021), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(G290), .B(G1986), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n1021), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n585), .B(KEYINPUT57), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1020), .A2(new_n1018), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n1019), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n1017), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT56), .B(G2072), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1040));
  NOR2_X1   g615(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n500), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT114), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n500), .A2(new_n1044), .A3(new_n1041), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1040), .A2(new_n1043), .A3(new_n1017), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1046), .A2(new_n1047), .A3(new_n798), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1046), .B2(new_n798), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1039), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1034), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1039), .B(new_n1034), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1040), .A2(new_n1017), .A3(new_n1042), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n793), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1020), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1017), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(G2067), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1054), .A2(new_n635), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1034), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1050), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT61), .B1(new_n1063), .B2(new_n1054), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g641(.A(KEYINPUT121), .B(KEYINPUT61), .C1(new_n1063), .C2(new_n1054), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1059), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT60), .A3(new_n635), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n635), .A2(KEYINPUT60), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n635), .A2(KEYINPUT60), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1071), .B1(new_n1059), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1035), .A2(new_n1017), .A3(new_n1022), .A4(new_n1036), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(new_n802), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1075), .A2(new_n1076), .B1(new_n1058), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1037), .A2(KEYINPUT119), .A3(new_n1022), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n567), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1074), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1054), .A2(KEYINPUT61), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n1053), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1061), .B1(new_n1068), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1035), .A2(new_n1036), .A3(new_n1017), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT124), .B1(new_n1089), .B2(G2078), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT53), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  OAI211_X1 g667(.A(KEYINPUT124), .B(new_n1092), .C1(new_n1089), .C2(G2078), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1055), .A2(new_n781), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G171), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1091), .A2(G301), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(KEYINPUT54), .A3(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT125), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G303), .A2(G8), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT55), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1089), .A2(new_n831), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1055), .A2(G2090), .ZN(new_n1105));
  OAI21_X1  g680(.A(G8), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1100), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G8), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1105), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(new_n1103), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT55), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1101), .B(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1112), .A3(KEYINPUT112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1103), .B1(G2090), .B2(new_n1046), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G8), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1102), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1108), .B1(new_n1017), .B2(new_n1057), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n849), .B2(G288), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT52), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT52), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n825), .B2(G1976), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1981), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n844), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(G1981), .B1(new_n839), .B2(new_n842), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT49), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT49), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1132), .A3(new_n1129), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1126), .B1(new_n1134), .B2(new_n1121), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1114), .A2(new_n1120), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G1966), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1089), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1040), .A2(new_n1017), .A3(new_n733), .A4(new_n1042), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1108), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(G286), .A2(G8), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT122), .Z(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT51), .B1(new_n1140), .B2(KEYINPUT123), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1141), .A2(KEYINPUT123), .A3(KEYINPUT51), .A4(new_n1143), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1149), .A2(new_n1143), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1146), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1136), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1153), .A2(KEYINPUT54), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1099), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1088), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1135), .A2(new_n1107), .A3(new_n1113), .ZN(new_n1157));
  AND4_X1   g732(.A1(new_n849), .A2(new_n1131), .A3(new_n825), .A4(new_n1133), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1128), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1121), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT113), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1157), .A2(new_n1160), .A3(KEYINPUT113), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1141), .A2(G286), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1114), .A2(new_n1120), .A3(new_n1135), .A4(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1140), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1114), .A2(new_n1135), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT116), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT116), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1114), .A2(new_n1174), .A3(new_n1171), .A4(new_n1135), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1169), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1136), .A2(new_n1096), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1146), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT62), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1146), .A2(new_n1147), .A3(new_n1180), .A4(new_n1150), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1177), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1165), .A2(new_n1176), .A3(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1033), .B1(new_n1156), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1024), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1185), .A2(KEYINPUT46), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(KEYINPUT46), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1021), .B1(new_n777), .B2(new_n1026), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT126), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT47), .ZN(new_n1191));
  INV_X1    g766(.A(new_n812), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1028), .A2(new_n1192), .A3(new_n815), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n763), .A2(G2067), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1021), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1025), .A2(G1986), .A3(G290), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT48), .Z(new_n1197));
  NAND2_X1  g772(.A1(new_n1030), .A2(new_n1197), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1191), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1184), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n1202));
  NOR3_X1   g776(.A1(new_n674), .A2(new_n459), .A3(G227), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n708), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n1204), .B1(new_n918), .B2(new_n920), .ZN(new_n1205));
  AND3_X1   g779(.A1(new_n1012), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g780(.A(new_n1202), .B1(new_n1012), .B2(new_n1205), .ZN(new_n1207));
  NOR2_X1   g781(.A1(new_n1206), .A2(new_n1207), .ZN(G308));
  NAND2_X1  g782(.A1(new_n1012), .A2(new_n1205), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n1209), .A2(KEYINPUT127), .ZN(new_n1210));
  NAND3_X1  g784(.A1(new_n1012), .A2(new_n1205), .A3(new_n1202), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n1211), .ZN(G225));
endmodule


