

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U554 ( .A(KEYINPUT97), .B(n704), .ZN(n803) );
  NOR2_X1 U555 ( .A1(n711), .A2(n710), .ZN(n713) );
  BUF_X1 U556 ( .A(n554), .Z(n534) );
  BUF_X1 U557 ( .A(n551), .Z(n525) );
  XNOR2_X1 U558 ( .A(n731), .B(n730), .ZN(n736) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n730) );
  NOR2_X1 U560 ( .A1(n745), .A2(n744), .ZN(n748) );
  NAND2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XOR2_X1 U562 ( .A(KEYINPUT23), .B(n549), .Z(n521) );
  AND2_X1 U563 ( .A1(n753), .A2(G8), .ZN(n522) );
  AND2_X1 U564 ( .A1(n835), .A2(n828), .ZN(n523) );
  INV_X1 U565 ( .A(KEYINPUT110), .ZN(n746) );
  XNOR2_X1 U566 ( .A(n746), .B(KEYINPUT31), .ZN(n747) );
  AND2_X1 U567 ( .A1(n766), .A2(n765), .ZN(n767) );
  INV_X1 U568 ( .A(KEYINPUT17), .ZN(n531) );
  INV_X1 U569 ( .A(KEYINPUT13), .ZN(n580) );
  XNOR2_X1 U570 ( .A(n531), .B(KEYINPUT68), .ZN(n532) );
  XNOR2_X1 U571 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U572 ( .A(n533), .B(n532), .ZN(n554) );
  NOR2_X2 U573 ( .A1(G651), .A2(G543), .ZN(n655) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n529), .ZN(n892) );
  NAND2_X1 U575 ( .A1(n523), .A2(n825), .ZN(n826) );
  OR2_X1 U576 ( .A1(n827), .A2(n826), .ZN(n842) );
  NOR2_X1 U577 ( .A1(G651), .A2(n671), .ZN(n665) );
  INV_X1 U578 ( .A(G2105), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n892), .A2(G126), .ZN(n527) );
  XOR2_X1 U580 ( .A(KEYINPUT66), .B(n524), .Z(n551) );
  NAND2_X1 U581 ( .A1(G114), .A2(n525), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U583 ( .A(KEYINPUT96), .B(n528), .ZN(n538) );
  NAND2_X1 U584 ( .A1(n529), .A2(G2104), .ZN(n530) );
  XNOR2_X1 U585 ( .A(n530), .B(KEYINPUT65), .ZN(n548) );
  BUF_X1 U586 ( .A(n548), .Z(n889) );
  NAND2_X1 U587 ( .A1(n889), .A2(G102), .ZN(n536) );
  NOR2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  NAND2_X1 U589 ( .A1(G138), .A2(n534), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U592 ( .A1(G91), .A2(n655), .ZN(n540) );
  XOR2_X1 U593 ( .A(G543), .B(KEYINPUT0), .Z(n671) );
  INV_X1 U594 ( .A(G651), .ZN(n541) );
  NOR2_X1 U595 ( .A1(n671), .A2(n541), .ZN(n657) );
  NAND2_X1 U596 ( .A1(G78), .A2(n657), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n546) );
  NOR2_X1 U598 ( .A1(G543), .A2(n541), .ZN(n542) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n542), .Z(n669) );
  NAND2_X1 U600 ( .A1(G65), .A2(n669), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G53), .A2(n665), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U604 ( .A(KEYINPUT72), .B(n547), .ZN(n725) );
  INV_X1 U605 ( .A(n725), .ZN(G299) );
  NAND2_X1 U606 ( .A1(G125), .A2(n892), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G101), .A2(n548), .ZN(n549) );
  AND2_X1 U608 ( .A1(n550), .A2(n521), .ZN(n559) );
  NAND2_X1 U609 ( .A1(G113), .A2(n551), .ZN(n553) );
  INV_X1 U610 ( .A(KEYINPUT67), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n553), .B(n552), .ZN(n556) );
  NAND2_X1 U612 ( .A1(G137), .A2(n554), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U614 ( .A(n557), .B(KEYINPUT69), .ZN(n558) );
  AND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U616 ( .A(n560), .B(KEYINPUT64), .ZN(n703) );
  BUF_X1 U617 ( .A(n703), .Z(G160) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G108), .ZN(G238) );
  INV_X1 U620 ( .A(G120), .ZN(G236) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  NAND2_X1 U624 ( .A1(G89), .A2(n655), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(KEYINPUT4), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT78), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G76), .A2(n657), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U629 ( .A(KEYINPUT5), .B(n565), .ZN(n571) );
  XNOR2_X1 U630 ( .A(KEYINPUT79), .B(KEYINPUT6), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G63), .A2(n669), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G51), .A2(n665), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT7), .B(n572), .ZN(G168) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n573) );
  XOR2_X1 U639 ( .A(n573), .B(KEYINPUT10), .Z(n844) );
  INV_X1 U640 ( .A(n844), .ZN(G223) );
  INV_X1 U641 ( .A(G567), .ZN(n697) );
  NOR2_X1 U642 ( .A1(n697), .A2(G223), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n574), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U644 ( .A1(n669), .A2(G56), .ZN(n575) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n575), .Z(n583) );
  NAND2_X1 U646 ( .A1(G81), .A2(n655), .ZN(n576) );
  XOR2_X1 U647 ( .A(KEYINPUT12), .B(n576), .Z(n577) );
  XNOR2_X1 U648 ( .A(n577), .B(KEYINPUT73), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G68), .A2(n657), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n581) );
  NOR2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n584), .B(KEYINPUT74), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G43), .A2(n665), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X2 U655 ( .A(KEYINPUT75), .B(n587), .ZN(n949) );
  XNOR2_X1 U656 ( .A(G860), .B(KEYINPUT76), .ZN(n608) );
  NAND2_X1 U657 ( .A1(n949), .A2(n608), .ZN(G153) );
  NAND2_X1 U658 ( .A1(G90), .A2(n655), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G77), .A2(n657), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n591) );
  XOR2_X1 U661 ( .A(KEYINPUT9), .B(KEYINPUT71), .Z(n590) );
  XNOR2_X1 U662 ( .A(n591), .B(n590), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G64), .A2(n669), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G52), .A2(n665), .ZN(n592) );
  AND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(G301) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n605) );
  NAND2_X1 U668 ( .A1(G79), .A2(n657), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G54), .A2(n665), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G92), .A2(n655), .ZN(n599) );
  NAND2_X1 U672 ( .A1(G66), .A2(n669), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U674 ( .A(KEYINPUT77), .B(n600), .Z(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U676 ( .A(KEYINPUT15), .B(n603), .Z(n940) );
  OR2_X1 U677 ( .A1(n940), .A2(G868), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(G284) );
  INV_X1 U679 ( .A(G868), .ZN(n683) );
  NOR2_X1 U680 ( .A1(G286), .A2(n683), .ZN(n607) );
  NOR2_X1 U681 ( .A1(G299), .A2(G868), .ZN(n606) );
  NOR2_X1 U682 ( .A1(n607), .A2(n606), .ZN(G297) );
  XOR2_X1 U683 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n613) );
  INV_X1 U684 ( .A(G559), .ZN(n609) );
  NOR2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U686 ( .A(KEYINPUT80), .B(n610), .Z(n611) );
  NAND2_X1 U687 ( .A1(n611), .A2(n940), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n613), .B(n612), .ZN(G148) );
  NAND2_X1 U689 ( .A1(n940), .A2(G868), .ZN(n614) );
  XOR2_X1 U690 ( .A(KEYINPUT83), .B(n614), .Z(n615) );
  NOR2_X1 U691 ( .A1(G559), .A2(n615), .ZN(n618) );
  INV_X1 U692 ( .A(n949), .ZN(n711) );
  NOR2_X1 U693 ( .A1(G868), .A2(n711), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n616), .B(KEYINPUT82), .ZN(n617) );
  NOR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(G282) );
  XOR2_X1 U696 ( .A(G2100), .B(KEYINPUT84), .Z(n627) );
  NAND2_X1 U697 ( .A1(G123), .A2(n892), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n619), .B(KEYINPUT18), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G111), .A2(n525), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n889), .A2(G99), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G135), .A2(n534), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n986) );
  XNOR2_X1 U705 ( .A(G2096), .B(n986), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(G156) );
  NAND2_X1 U707 ( .A1(G67), .A2(n669), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G55), .A2(n665), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U710 ( .A(KEYINPUT86), .B(n630), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G93), .A2(n655), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G80), .A2(n657), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  OR2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n682) );
  NAND2_X1 U715 ( .A1(G559), .A2(n940), .ZN(n635) );
  XOR2_X1 U716 ( .A(n949), .B(n635), .Z(n680) );
  NOR2_X1 U717 ( .A1(G860), .A2(n680), .ZN(n637) );
  XNOR2_X1 U718 ( .A(KEYINPUT85), .B(KEYINPUT87), .ZN(n636) );
  XNOR2_X1 U719 ( .A(n637), .B(n636), .ZN(n638) );
  XOR2_X1 U720 ( .A(n682), .B(n638), .Z(G145) );
  NAND2_X1 U721 ( .A1(G86), .A2(n655), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G61), .A2(n669), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n657), .A2(G73), .ZN(n641) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n641), .Z(n642) );
  NOR2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n665), .A2(G48), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U729 ( .A1(G85), .A2(n655), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G72), .A2(n657), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U732 ( .A(KEYINPUT70), .B(n648), .Z(n652) );
  NAND2_X1 U733 ( .A1(G60), .A2(n669), .ZN(n650) );
  NAND2_X1 U734 ( .A1(G47), .A2(n665), .ZN(n649) );
  AND2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U736 ( .A1(n652), .A2(n651), .ZN(G290) );
  NAND2_X1 U737 ( .A1(G62), .A2(n669), .ZN(n654) );
  NAND2_X1 U738 ( .A1(G50), .A2(n665), .ZN(n653) );
  NAND2_X1 U739 ( .A1(n654), .A2(n653), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n655), .A2(G88), .ZN(n656) );
  XNOR2_X1 U741 ( .A(KEYINPUT89), .B(n656), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n657), .A2(G75), .ZN(n658) );
  XOR2_X1 U743 ( .A(KEYINPUT90), .B(n658), .Z(n659) );
  NOR2_X1 U744 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U745 ( .A(n661), .B(KEYINPUT91), .ZN(n662) );
  NOR2_X1 U746 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U747 ( .A(KEYINPUT92), .B(n664), .ZN(G166) );
  NAND2_X1 U748 ( .A1(G49), .A2(n665), .ZN(n667) );
  NAND2_X1 U749 ( .A1(G74), .A2(G651), .ZN(n666) );
  NAND2_X1 U750 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U751 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n670), .B(KEYINPUT88), .ZN(n673) );
  NAND2_X1 U753 ( .A1(G87), .A2(n671), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n673), .A2(n672), .ZN(G288) );
  XOR2_X1 U755 ( .A(KEYINPUT93), .B(KEYINPUT19), .Z(n674) );
  XNOR2_X1 U756 ( .A(G305), .B(n674), .ZN(n675) );
  XOR2_X1 U757 ( .A(n682), .B(n675), .Z(n677) );
  XOR2_X1 U758 ( .A(G290), .B(G166), .Z(n676) );
  XNOR2_X1 U759 ( .A(n677), .B(n676), .ZN(n678) );
  XOR2_X1 U760 ( .A(n678), .B(G299), .Z(n679) );
  XNOR2_X1 U761 ( .A(n679), .B(G288), .ZN(n907) );
  XOR2_X1 U762 ( .A(n680), .B(n907), .Z(n681) );
  NAND2_X1 U763 ( .A1(n681), .A2(G868), .ZN(n685) );
  NAND2_X1 U764 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n685), .A2(n684), .ZN(G295) );
  NAND2_X1 U766 ( .A1(G2084), .A2(G2078), .ZN(n686) );
  XOR2_X1 U767 ( .A(KEYINPUT20), .B(n686), .Z(n687) );
  NAND2_X1 U768 ( .A1(G2090), .A2(n687), .ZN(n688) );
  XNOR2_X1 U769 ( .A(KEYINPUT21), .B(n688), .ZN(n689) );
  NAND2_X1 U770 ( .A1(n689), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U771 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n690) );
  XNOR2_X1 U773 ( .A(KEYINPUT22), .B(n690), .ZN(n691) );
  NAND2_X1 U774 ( .A1(n691), .A2(G96), .ZN(n692) );
  NOR2_X1 U775 ( .A1(G218), .A2(n692), .ZN(n693) );
  XOR2_X1 U776 ( .A(KEYINPUT94), .B(n693), .Z(n929) );
  NAND2_X1 U777 ( .A1(n929), .A2(G2106), .ZN(n694) );
  XNOR2_X1 U778 ( .A(n694), .B(KEYINPUT95), .ZN(n699) );
  NOR2_X1 U779 ( .A1(G236), .A2(G238), .ZN(n695) );
  NAND2_X1 U780 ( .A1(G69), .A2(n695), .ZN(n696) );
  NOR2_X1 U781 ( .A1(G237), .A2(n696), .ZN(n928) );
  NOR2_X1 U782 ( .A1(n697), .A2(n928), .ZN(n698) );
  NOR2_X1 U783 ( .A1(n699), .A2(n698), .ZN(G319) );
  INV_X1 U784 ( .A(G319), .ZN(n701) );
  NAND2_X1 U785 ( .A1(G483), .A2(G661), .ZN(n700) );
  NOR2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n846) );
  NAND2_X1 U787 ( .A1(n846), .A2(G36), .ZN(G176) );
  INV_X1 U788 ( .A(G166), .ZN(G303) );
  INV_X1 U789 ( .A(G301), .ZN(G171) );
  NOR2_X1 U790 ( .A1(G1976), .A2(G288), .ZN(n939) );
  NOR2_X1 U791 ( .A1(G303), .A2(G1971), .ZN(n702) );
  NOR2_X1 U792 ( .A1(n939), .A2(n702), .ZN(n770) );
  NOR2_X1 U793 ( .A1(G164), .A2(G1384), .ZN(n802) );
  INV_X1 U794 ( .A(n802), .ZN(n705) );
  AND2_X1 U795 ( .A1(n703), .A2(G40), .ZN(n704) );
  NOR2_X4 U796 ( .A1(n705), .A2(n803), .ZN(n737) );
  AND2_X1 U797 ( .A1(n737), .A2(G1996), .ZN(n707) );
  XOR2_X1 U798 ( .A(KEYINPUT26), .B(KEYINPUT108), .Z(n706) );
  XNOR2_X1 U799 ( .A(n707), .B(n706), .ZN(n709) );
  INV_X1 U800 ( .A(n737), .ZN(n759) );
  NAND2_X1 U801 ( .A1(n759), .A2(G1341), .ZN(n708) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U803 ( .A1(n713), .A2(n940), .ZN(n712) );
  XNOR2_X1 U804 ( .A(n712), .B(KEYINPUT109), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n713), .A2(n940), .ZN(n717) );
  NOR2_X1 U806 ( .A1(G2067), .A2(n759), .ZN(n715) );
  NOR2_X1 U807 ( .A1(n737), .A2(G1348), .ZN(n714) );
  NOR2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n724) );
  NAND2_X1 U811 ( .A1(n737), .A2(G2072), .ZN(n720) );
  XNOR2_X1 U812 ( .A(n720), .B(KEYINPUT27), .ZN(n722) );
  XNOR2_X1 U813 ( .A(G1956), .B(KEYINPUT107), .ZN(n959) );
  NOR2_X1 U814 ( .A1(n959), .A2(n737), .ZN(n721) );
  NOR2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n726), .A2(n725), .ZN(n723) );
  NAND2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U819 ( .A(n727), .B(KEYINPUT28), .Z(n728) );
  NAND2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n731) );
  NOR2_X1 U821 ( .A1(n737), .A2(G1961), .ZN(n732) );
  XOR2_X1 U822 ( .A(KEYINPUT106), .B(n732), .Z(n734) );
  XNOR2_X1 U823 ( .A(G2078), .B(KEYINPUT25), .ZN(n1014) );
  NAND2_X1 U824 ( .A1(n737), .A2(n1014), .ZN(n733) );
  NAND2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n743) );
  NAND2_X1 U826 ( .A1(n743), .A2(G171), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n750) );
  NAND2_X1 U828 ( .A1(G8), .A2(n759), .ZN(n787) );
  NOR2_X1 U829 ( .A1(G1966), .A2(n787), .ZN(n751) );
  INV_X1 U830 ( .A(n751), .ZN(n740) );
  INV_X1 U831 ( .A(G2084), .ZN(n738) );
  AND2_X1 U832 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U833 ( .A(n739), .B(KEYINPUT105), .ZN(n753) );
  NAND2_X1 U834 ( .A1(n740), .A2(n522), .ZN(n741) );
  XNOR2_X1 U835 ( .A(n741), .B(KEYINPUT30), .ZN(n742) );
  NOR2_X1 U836 ( .A1(G168), .A2(n742), .ZN(n745) );
  NOR2_X1 U837 ( .A1(G171), .A2(n743), .ZN(n744) );
  XNOR2_X1 U838 ( .A(n748), .B(n747), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n758) );
  XNOR2_X1 U840 ( .A(KEYINPUT111), .B(n758), .ZN(n752) );
  NOR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n756) );
  INV_X1 U842 ( .A(n753), .ZN(n754) );
  NAND2_X1 U843 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n769) );
  AND2_X1 U845 ( .A1(G286), .A2(G8), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n766) );
  INV_X1 U847 ( .A(G8), .ZN(n764) );
  NOR2_X1 U848 ( .A1(G1971), .A2(n787), .ZN(n761) );
  NOR2_X1 U849 ( .A1(G2090), .A2(n759), .ZN(n760) );
  NOR2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n762), .A2(G303), .ZN(n763) );
  OR2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U853 ( .A(n767), .B(KEYINPUT32), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n769), .A2(n768), .ZN(n781) );
  AND2_X1 U855 ( .A1(n770), .A2(n781), .ZN(n773) );
  NAND2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n935) );
  INV_X1 U857 ( .A(n787), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n935), .A2(n771), .ZN(n772) );
  NOR2_X2 U859 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U860 ( .A1(KEYINPUT33), .A2(n774), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n939), .A2(KEYINPUT33), .ZN(n775) );
  NOR2_X1 U862 ( .A1(n775), .A2(n787), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U864 ( .A(G1981), .B(G305), .Z(n932) );
  AND2_X1 U865 ( .A1(n778), .A2(n932), .ZN(n791) );
  NOR2_X1 U866 ( .A1(G303), .A2(G2090), .ZN(n779) );
  XNOR2_X1 U867 ( .A(n779), .B(KEYINPUT112), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n780), .A2(G8), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n783), .A2(n787), .ZN(n789) );
  NOR2_X1 U871 ( .A1(G1981), .A2(G305), .ZN(n784) );
  XOR2_X1 U872 ( .A(n784), .B(KEYINPUT24), .Z(n785) );
  XNOR2_X1 U873 ( .A(KEYINPUT104), .B(n785), .ZN(n786) );
  OR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U876 ( .A1(n791), .A2(n790), .ZN(n827) );
  XNOR2_X1 U877 ( .A(KEYINPUT37), .B(G2067), .ZN(n837) );
  NAND2_X1 U878 ( .A1(n889), .A2(G104), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G140), .A2(n534), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n795) );
  XOR2_X1 U881 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n794) );
  XNOR2_X1 U882 ( .A(n795), .B(n794), .ZN(n800) );
  NAND2_X1 U883 ( .A1(n892), .A2(G128), .ZN(n797) );
  NAND2_X1 U884 ( .A1(G116), .A2(n525), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U886 ( .A(KEYINPUT35), .B(n798), .Z(n799) );
  NOR2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U888 ( .A(KEYINPUT36), .B(n801), .ZN(n885) );
  NOR2_X1 U889 ( .A1(n837), .A2(n885), .ZN(n995) );
  NOR2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U891 ( .A(n804), .B(KEYINPUT98), .ZN(n839) );
  NAND2_X1 U892 ( .A1(n995), .A2(n839), .ZN(n805) );
  XNOR2_X1 U893 ( .A(n805), .B(KEYINPUT100), .ZN(n835) );
  NAND2_X1 U894 ( .A1(n889), .A2(G95), .ZN(n812) );
  NAND2_X1 U895 ( .A1(G119), .A2(n892), .ZN(n807) );
  NAND2_X1 U896 ( .A1(G131), .A2(n534), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G107), .A2(n525), .ZN(n808) );
  XNOR2_X1 U899 ( .A(KEYINPUT101), .B(n808), .ZN(n809) );
  NOR2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U902 ( .A(KEYINPUT102), .B(n813), .ZN(n883) );
  AND2_X1 U903 ( .A1(n883), .A2(G1991), .ZN(n823) );
  NAND2_X1 U904 ( .A1(G129), .A2(n892), .ZN(n815) );
  NAND2_X1 U905 ( .A1(G141), .A2(n534), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n815), .A2(n814), .ZN(n819) );
  NAND2_X1 U907 ( .A1(G105), .A2(n889), .ZN(n816) );
  XNOR2_X1 U908 ( .A(n816), .B(KEYINPUT103), .ZN(n817) );
  XNOR2_X1 U909 ( .A(n817), .B(KEYINPUT38), .ZN(n818) );
  NOR2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U911 ( .A1(G117), .A2(n525), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n899) );
  AND2_X1 U913 ( .A1(n899), .A2(G1996), .ZN(n822) );
  NOR2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n989) );
  INV_X1 U915 ( .A(n989), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n839), .A2(n824), .ZN(n828) );
  XNOR2_X1 U917 ( .A(G1986), .B(G290), .ZN(n938) );
  NAND2_X1 U918 ( .A1(n938), .A2(n839), .ZN(n825) );
  NOR2_X1 U919 ( .A1(G1996), .A2(n899), .ZN(n984) );
  INV_X1 U920 ( .A(n828), .ZN(n832) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n829) );
  NOR2_X1 U922 ( .A1(n883), .A2(G1991), .ZN(n987) );
  NOR2_X1 U923 ( .A1(n829), .A2(n987), .ZN(n830) );
  XOR2_X1 U924 ( .A(KEYINPUT113), .B(n830), .Z(n831) );
  NOR2_X1 U925 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U926 ( .A1(n984), .A2(n833), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n834), .B(KEYINPUT39), .ZN(n836) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(n838) );
  NAND2_X1 U929 ( .A1(n837), .A2(n885), .ZN(n1004) );
  NAND2_X1 U930 ( .A1(n838), .A2(n1004), .ZN(n840) );
  NAND2_X1 U931 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U932 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U933 ( .A(n843), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U936 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G1), .A2(G3), .ZN(n847) );
  NAND2_X1 U938 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U939 ( .A(n848), .B(KEYINPUT114), .ZN(G188) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2072), .Z(n850) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2078), .ZN(n849) );
  XNOR2_X1 U942 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U943 ( .A(n851), .B(G2096), .Z(n853) );
  XNOR2_X1 U944 ( .A(G2084), .B(G2090), .ZN(n852) );
  XNOR2_X1 U945 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U946 ( .A(G2100), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U947 ( .A(KEYINPUT115), .B(G2678), .ZN(n854) );
  XNOR2_X1 U948 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U949 ( .A(n857), .B(n856), .Z(G227) );
  XOR2_X1 U950 ( .A(KEYINPUT117), .B(G1961), .Z(n859) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U952 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U953 ( .A(n860), .B(KEYINPUT41), .Z(n862) );
  XNOR2_X1 U954 ( .A(G1971), .B(G1976), .ZN(n861) );
  XNOR2_X1 U955 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U956 ( .A(G1981), .B(G1956), .Z(n864) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1966), .ZN(n863) );
  XNOR2_X1 U958 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U959 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U960 ( .A(KEYINPUT116), .B(G2474), .ZN(n867) );
  XNOR2_X1 U961 ( .A(n868), .B(n867), .ZN(G229) );
  NAND2_X1 U962 ( .A1(G124), .A2(n892), .ZN(n869) );
  XNOR2_X1 U963 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U964 ( .A1(G112), .A2(n525), .ZN(n870) );
  NAND2_X1 U965 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U966 ( .A1(n889), .A2(G100), .ZN(n873) );
  NAND2_X1 U967 ( .A1(G136), .A2(n534), .ZN(n872) );
  NAND2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U969 ( .A1(n875), .A2(n874), .ZN(G162) );
  NAND2_X1 U970 ( .A1(n892), .A2(G130), .ZN(n877) );
  NAND2_X1 U971 ( .A1(G118), .A2(n525), .ZN(n876) );
  NAND2_X1 U972 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U973 ( .A1(n889), .A2(G106), .ZN(n879) );
  NAND2_X1 U974 ( .A1(G142), .A2(n534), .ZN(n878) );
  NAND2_X1 U975 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U976 ( .A(n880), .B(KEYINPUT45), .Z(n881) );
  NOR2_X1 U977 ( .A1(n882), .A2(n881), .ZN(n884) );
  XOR2_X1 U978 ( .A(n884), .B(n883), .Z(n905) );
  XNOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n887) );
  XNOR2_X1 U980 ( .A(n885), .B(G162), .ZN(n886) );
  XNOR2_X1 U981 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U982 ( .A(G164), .B(n888), .ZN(n903) );
  NAND2_X1 U983 ( .A1(n889), .A2(G103), .ZN(n891) );
  NAND2_X1 U984 ( .A1(G139), .A2(n534), .ZN(n890) );
  NAND2_X1 U985 ( .A1(n891), .A2(n890), .ZN(n897) );
  NAND2_X1 U986 ( .A1(n892), .A2(G127), .ZN(n894) );
  NAND2_X1 U987 ( .A1(G115), .A2(n525), .ZN(n893) );
  NAND2_X1 U988 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n895), .Z(n896) );
  NOR2_X1 U990 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U991 ( .A(KEYINPUT118), .B(n898), .Z(n997) );
  XNOR2_X1 U992 ( .A(n997), .B(n986), .ZN(n901) );
  XOR2_X1 U993 ( .A(G160), .B(n899), .Z(n900) );
  XNOR2_X1 U994 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U995 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U996 ( .A(n905), .B(n904), .Z(n906) );
  NOR2_X1 U997 ( .A1(G37), .A2(n906), .ZN(G395) );
  XOR2_X1 U998 ( .A(n907), .B(G286), .Z(n909) );
  XOR2_X1 U999 ( .A(G301), .B(n940), .Z(n908) );
  XNOR2_X1 U1000 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1001 ( .A(n949), .B(n910), .ZN(n911) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n911), .ZN(n912) );
  XOR2_X1 U1003 ( .A(KEYINPUT119), .B(n912), .Z(G397) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(KEYINPUT120), .ZN(n914) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1006 ( .A(n914), .B(n913), .ZN(n925) );
  XOR2_X1 U1007 ( .A(G2451), .B(G2430), .Z(n916) );
  XNOR2_X1 U1008 ( .A(G2438), .B(G2443), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n916), .B(n915), .ZN(n922) );
  XOR2_X1 U1010 ( .A(G2435), .B(G2454), .Z(n918) );
  XNOR2_X1 U1011 ( .A(G1348), .B(G1341), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n920) );
  XOR2_X1 U1013 ( .A(G2446), .B(G2427), .Z(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1015 ( .A(n922), .B(n921), .Z(n923) );
  NAND2_X1 U1016 ( .A1(G14), .A2(n923), .ZN(n931) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n931), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(n927) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1020 ( .A1(n927), .A2(n926), .ZN(G225) );
  XNOR2_X1 U1021 ( .A(KEYINPUT121), .B(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(G96), .ZN(G221) );
  INV_X1 U1024 ( .A(n928), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(G325) );
  INV_X1 U1026 ( .A(G325), .ZN(G261) );
  INV_X1 U1027 ( .A(G69), .ZN(G235) );
  INV_X1 U1028 ( .A(n931), .ZN(G401) );
  INV_X1 U1029 ( .A(G16), .ZN(n979) );
  XOR2_X1 U1030 ( .A(n979), .B(KEYINPUT56), .Z(n955) );
  XNOR2_X1 U1031 ( .A(G1966), .B(G168), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(KEYINPUT57), .ZN(n953) );
  XOR2_X1 U1034 ( .A(G1971), .B(G303), .Z(n948) );
  XOR2_X1 U1035 ( .A(G299), .B(G1956), .Z(n936) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n946) );
  XOR2_X1 U1037 ( .A(G1961), .B(G171), .Z(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n944) );
  XOR2_X1 U1039 ( .A(n939), .B(KEYINPUT125), .Z(n942) );
  XOR2_X1 U1040 ( .A(G1348), .B(n940), .Z(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1045 ( .A(G1341), .B(n949), .Z(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n981) );
  XNOR2_X1 U1049 ( .A(G1341), .B(G19), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G1981), .B(G6), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT126), .B(n958), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(n959), .B(G20), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1055 ( .A(KEYINPUT59), .B(G1348), .Z(n962) );
  XNOR2_X1 U1056 ( .A(G4), .B(n962), .ZN(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT60), .B(n965), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G21), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G5), .B(G1961), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n976) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G22), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(G23), .B(G1976), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n973) );
  XOR2_X1 U1066 ( .A(G1986), .B(G24), .Z(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(KEYINPUT58), .B(n974), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(KEYINPUT61), .B(n977), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n982), .B(KEYINPUT127), .ZN(n1010) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1076 ( .A(KEYINPUT51), .B(n985), .Z(n993) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n991) );
  XOR2_X1 U1079 ( .A(G2084), .B(G160), .Z(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1083 ( .A(KEYINPUT122), .B(n996), .Z(n1002) );
  XOR2_X1 U1084 ( .A(G164), .B(G2078), .Z(n999) );
  XNOR2_X1 U1085 ( .A(G2072), .B(n997), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(KEYINPUT50), .B(n1000), .Z(n1001) );
  NOR2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(n1005), .B(KEYINPUT52), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(KEYINPUT123), .B(n1006), .ZN(n1007) );
  INV_X1 U1092 ( .A(KEYINPUT55), .ZN(n1027) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1027), .ZN(n1008) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(G29), .ZN(n1009) );
  NAND2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1034) );
  XNOR2_X1 U1096 ( .A(G1996), .B(G32), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G33), .B(G2072), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1020) );
  XOR2_X1 U1099 ( .A(G2067), .B(G26), .Z(n1013) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(G28), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(n1014), .B(G27), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(G1991), .B(G25), .Z(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1021), .B(KEYINPUT53), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(G2084), .B(G34), .Z(n1022) );
  XNOR2_X1 U1108 ( .A(KEYINPUT54), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(G35), .B(G2090), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(n1028), .B(n1027), .Z(n1030) );
  INV_X1 U1113 ( .A(G29), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1115 ( .A1(G11), .A2(n1031), .ZN(n1032) );
  XNOR2_X1 U1116 ( .A(KEYINPUT124), .B(n1032), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1035), .Z(G150) );
  INV_X1 U1119 ( .A(G150), .ZN(G311) );
endmodule

