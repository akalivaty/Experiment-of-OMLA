

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579;

  XOR2_X1 U323 ( .A(n418), .B(n417), .Z(n291) );
  XOR2_X1 U324 ( .A(n420), .B(G204GAT), .Z(n292) );
  XNOR2_X1 U325 ( .A(KEYINPUT26), .B(n446), .ZN(n527) );
  NOR2_X1 U326 ( .A1(n466), .A2(n465), .ZN(n478) );
  XOR2_X1 U327 ( .A(n426), .B(n425), .Z(n543) );
  INV_X1 U328 ( .A(G204GAT), .ZN(n451) );
  XNOR2_X1 U329 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n449) );
  XOR2_X1 U330 ( .A(KEYINPUT17), .B(G190GAT), .Z(n294) );
  XNOR2_X1 U331 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n293) );
  XNOR2_X1 U332 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U333 ( .A(KEYINPUT19), .B(n295), .Z(n440) );
  XOR2_X1 U334 ( .A(G169GAT), .B(G8GAT), .Z(n330) );
  XOR2_X1 U335 ( .A(n330), .B(KEYINPUT79), .Z(n297) );
  NAND2_X1 U336 ( .A1(G226GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U338 ( .A(G92GAT), .B(G64GAT), .Z(n299) );
  XNOR2_X1 U339 ( .A(G204GAT), .B(KEYINPUT73), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U341 ( .A(G176GAT), .B(n300), .Z(n320) );
  XOR2_X1 U342 ( .A(n301), .B(n320), .Z(n307) );
  XNOR2_X1 U343 ( .A(G211GAT), .B(KEYINPUT90), .ZN(n302) );
  XNOR2_X1 U344 ( .A(n302), .B(KEYINPUT21), .ZN(n303) );
  XOR2_X1 U345 ( .A(n303), .B(KEYINPUT91), .Z(n305) );
  XNOR2_X1 U346 ( .A(G197GAT), .B(G218GAT), .ZN(n304) );
  XNOR2_X1 U347 ( .A(n305), .B(n304), .ZN(n424) );
  XNOR2_X1 U348 ( .A(G36GAT), .B(n424), .ZN(n306) );
  XNOR2_X1 U349 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U350 ( .A(n440), .B(n308), .ZN(n509) );
  XNOR2_X1 U351 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n385) );
  XOR2_X1 U352 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n310) );
  XNOR2_X1 U353 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n309) );
  XNOR2_X1 U354 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U355 ( .A(G106GAT), .B(G78GAT), .Z(n418) );
  XOR2_X1 U356 ( .A(G99GAT), .B(G85GAT), .Z(n373) );
  XNOR2_X1 U357 ( .A(n418), .B(n373), .ZN(n312) );
  XOR2_X1 U358 ( .A(KEYINPUT72), .B(KEYINPUT74), .Z(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U360 ( .A(n314), .B(n313), .Z(n316) );
  NAND2_X1 U361 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n318) );
  XNOR2_X1 U363 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n317) );
  XNOR2_X1 U364 ( .A(n317), .B(KEYINPUT13), .ZN(n349) );
  XNOR2_X1 U365 ( .A(n318), .B(n349), .ZN(n322) );
  XNOR2_X1 U366 ( .A(G120GAT), .B(G148GAT), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n319), .B(G57GAT), .ZN(n400) );
  XNOR2_X1 U368 ( .A(n400), .B(n320), .ZN(n321) );
  XNOR2_X1 U369 ( .A(n322), .B(n321), .ZN(n454) );
  INV_X1 U370 ( .A(KEYINPUT41), .ZN(n323) );
  XNOR2_X1 U371 ( .A(n454), .B(n323), .ZN(n533) );
  XOR2_X1 U372 ( .A(KEYINPUT7), .B(KEYINPUT69), .Z(n325) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(G36GAT), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U375 ( .A(KEYINPUT8), .B(n326), .ZN(n381) );
  XOR2_X1 U376 ( .A(KEYINPUT66), .B(KEYINPUT68), .Z(n328) );
  XNOR2_X1 U377 ( .A(G197GAT), .B(G15GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U379 ( .A(n330), .B(n329), .Z(n332) );
  NAND2_X1 U380 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U382 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n334) );
  XNOR2_X1 U383 ( .A(KEYINPUT65), .B(KEYINPUT29), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U385 ( .A(n336), .B(n335), .Z(n340) );
  XNOR2_X1 U386 ( .A(G50GAT), .B(G22GAT), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n337), .B(G141GAT), .ZN(n421) );
  XNOR2_X1 U388 ( .A(G29GAT), .B(G113GAT), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n338), .B(G1GAT), .ZN(n411) );
  XNOR2_X1 U390 ( .A(n421), .B(n411), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n381), .B(n341), .ZN(n567) );
  NAND2_X1 U393 ( .A1(n533), .A2(n567), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n342), .B(KEYINPUT46), .ZN(n363) );
  XOR2_X1 U395 ( .A(G155GAT), .B(G127GAT), .Z(n344) );
  XNOR2_X1 U396 ( .A(G22GAT), .B(G183GAT), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U398 ( .A(KEYINPUT79), .B(G64GAT), .Z(n346) );
  XNOR2_X1 U399 ( .A(G8GAT), .B(G15GAT), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U401 ( .A(n348), .B(n347), .Z(n354) );
  XOR2_X1 U402 ( .A(G78GAT), .B(n349), .Z(n351) );
  NAND2_X1 U403 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U405 ( .A(G211GAT), .B(n352), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n362) );
  XOR2_X1 U407 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n356) );
  XNOR2_X1 U408 ( .A(G57GAT), .B(KEYINPUT15), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U410 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n358) );
  XNOR2_X1 U411 ( .A(G1GAT), .B(KEYINPUT82), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U413 ( .A(n360), .B(n359), .Z(n361) );
  XOR2_X1 U414 ( .A(n362), .B(n361), .Z(n572) );
  INV_X1 U415 ( .A(n572), .ZN(n557) );
  NAND2_X1 U416 ( .A1(n363), .A2(n557), .ZN(n364) );
  XNOR2_X1 U417 ( .A(n364), .B(KEYINPUT111), .ZN(n383) );
  XOR2_X1 U418 ( .A(G92GAT), .B(G162GAT), .Z(n366) );
  XNOR2_X1 U419 ( .A(G190GAT), .B(G134GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n380) );
  XOR2_X1 U421 ( .A(KEYINPUT78), .B(KEYINPUT76), .Z(n368) );
  XNOR2_X1 U422 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U424 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n370) );
  XNOR2_X1 U425 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U427 ( .A(n372), .B(n371), .Z(n378) );
  XOR2_X1 U428 ( .A(G29GAT), .B(n373), .Z(n375) );
  NAND2_X1 U429 ( .A1(G232GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U431 ( .A(G50GAT), .B(n376), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n382) );
  XNOR2_X1 U434 ( .A(n382), .B(n381), .ZN(n564) );
  NAND2_X1 U435 ( .A1(n383), .A2(n564), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n385), .B(n384), .ZN(n392) );
  XOR2_X1 U437 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n388) );
  XOR2_X1 U438 ( .A(KEYINPUT36), .B(KEYINPUT103), .Z(n386) );
  XOR2_X1 U439 ( .A(n564), .B(n386), .Z(n577) );
  NAND2_X1 U440 ( .A1(n572), .A2(n577), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U442 ( .A(KEYINPUT70), .B(n567), .Z(n549) );
  NAND2_X1 U443 ( .A1(n389), .A2(n549), .ZN(n390) );
  NOR2_X1 U444 ( .A1(n454), .A2(n390), .ZN(n391) );
  NOR2_X1 U445 ( .A1(n392), .A2(n391), .ZN(n393) );
  XNOR2_X1 U446 ( .A(KEYINPUT48), .B(n393), .ZN(n528) );
  NOR2_X1 U447 ( .A1(n509), .A2(n528), .ZN(n394) );
  XNOR2_X1 U448 ( .A(KEYINPUT54), .B(n394), .ZN(n414) );
  XOR2_X1 U449 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n396) );
  NAND2_X1 U450 ( .A1(G225GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U452 ( .A(n397), .B(KEYINPUT6), .Z(n402) );
  XOR2_X1 U453 ( .A(G127GAT), .B(KEYINPUT84), .Z(n399) );
  XNOR2_X1 U454 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n433) );
  XNOR2_X1 U456 ( .A(n433), .B(n400), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U458 ( .A(G85GAT), .B(KEYINPUT4), .Z(n404) );
  XNOR2_X1 U459 ( .A(G141GAT), .B(KEYINPUT94), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U461 ( .A(n406), .B(n405), .Z(n413) );
  XOR2_X1 U462 ( .A(KEYINPUT92), .B(G162GAT), .Z(n408) );
  XNOR2_X1 U463 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U465 ( .A(KEYINPUT2), .B(n409), .Z(n425) );
  INV_X1 U466 ( .A(n425), .ZN(n410) );
  XOR2_X1 U467 ( .A(n411), .B(n410), .Z(n412) );
  XOR2_X1 U468 ( .A(n413), .B(n412), .Z(n461) );
  XNOR2_X1 U469 ( .A(KEYINPUT95), .B(n461), .ZN(n505) );
  NAND2_X1 U470 ( .A1(n414), .A2(n505), .ZN(n544) );
  XOR2_X1 U471 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n416) );
  XNOR2_X1 U472 ( .A(KEYINPUT24), .B(G148GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n291), .B(n419), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(KEYINPUT93), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n292), .B(n422), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U479 ( .A(KEYINPUT89), .B(G120GAT), .Z(n428) );
  XNOR2_X1 U480 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U482 ( .A(KEYINPUT86), .B(G176GAT), .Z(n430) );
  XNOR2_X1 U483 ( .A(G113GAT), .B(G71GAT), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n444) );
  XOR2_X1 U486 ( .A(G99GAT), .B(n433), .Z(n435) );
  NAND2_X1 U487 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U489 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n437) );
  XNOR2_X1 U490 ( .A(G169GAT), .B(G15GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n439), .B(n438), .Z(n442) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X2 U495 ( .A(n444), .B(n443), .Z(n511) );
  NAND2_X1 U496 ( .A1(n543), .A2(n511), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n445), .B(KEYINPUT98), .ZN(n446) );
  NOR2_X1 U498 ( .A1(n544), .A2(n527), .ZN(n447) );
  XOR2_X1 U499 ( .A(n447), .B(KEYINPUT123), .Z(n576) );
  AND2_X1 U500 ( .A1(n576), .A2(n454), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(G1353GAT) );
  XOR2_X1 U503 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n453) );
  XNOR2_X1 U504 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(n471) );
  NOR2_X1 U506 ( .A1(n549), .A2(n454), .ZN(n482) );
  NOR2_X1 U507 ( .A1(n511), .A2(n509), .ZN(n455) );
  NOR2_X1 U508 ( .A1(n543), .A2(n455), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n456), .B(KEYINPUT99), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n457), .B(KEYINPUT25), .ZN(n460) );
  XNOR2_X1 U511 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n458), .B(n509), .ZN(n463) );
  NOR2_X1 U513 ( .A1(n463), .A2(n527), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n460), .A2(n459), .ZN(n462) );
  NOR2_X1 U515 ( .A1(n462), .A2(n461), .ZN(n466) );
  INV_X1 U516 ( .A(n511), .ZN(n548) );
  NOR2_X1 U517 ( .A1(n505), .A2(n463), .ZN(n464) );
  XOR2_X1 U518 ( .A(KEYINPUT97), .B(n464), .Z(n530) );
  XOR2_X1 U519 ( .A(KEYINPUT28), .B(n543), .Z(n514) );
  NAND2_X1 U520 ( .A1(n530), .A2(n514), .ZN(n517) );
  NOR2_X1 U521 ( .A1(n548), .A2(n517), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT83), .B(KEYINPUT16), .Z(n468) );
  NAND2_X1 U523 ( .A1(n572), .A2(n564), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n468), .B(n467), .ZN(n469) );
  NOR2_X1 U525 ( .A1(n478), .A2(n469), .ZN(n492) );
  NAND2_X1 U526 ( .A1(n482), .A2(n492), .ZN(n476) );
  NOR2_X1 U527 ( .A1(n505), .A2(n476), .ZN(n470) );
  XOR2_X1 U528 ( .A(n471), .B(n470), .Z(G1324GAT) );
  NOR2_X1 U529 ( .A1(n509), .A2(n476), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT102), .B(n472), .Z(n473) );
  XNOR2_X1 U531 ( .A(G8GAT), .B(n473), .ZN(G1325GAT) );
  NOR2_X1 U532 ( .A1(n511), .A2(n476), .ZN(n475) );
  XNOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  NOR2_X1 U535 ( .A1(n514), .A2(n476), .ZN(n477) );
  XOR2_X1 U536 ( .A(G22GAT), .B(n477), .Z(G1327GAT) );
  NOR2_X1 U537 ( .A1(n572), .A2(n478), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n577), .A2(n479), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(KEYINPUT37), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT104), .ZN(n503) );
  NAND2_X1 U541 ( .A1(n503), .A2(n482), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n483), .B(KEYINPUT38), .ZN(n490) );
  NOR2_X1 U543 ( .A1(n505), .A2(n490), .ZN(n486) );
  XOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT105), .Z(n484) );
  XNOR2_X1 U545 ( .A(KEYINPUT39), .B(n484), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  NOR2_X1 U547 ( .A1(n490), .A2(n509), .ZN(n487) );
  XOR2_X1 U548 ( .A(G36GAT), .B(n487), .Z(G1329GAT) );
  NOR2_X1 U549 ( .A1(n490), .A2(n511), .ZN(n488) );
  XOR2_X1 U550 ( .A(KEYINPUT40), .B(n488), .Z(n489) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(n489), .ZN(G1330GAT) );
  NOR2_X1 U552 ( .A1(n490), .A2(n514), .ZN(n491) );
  XOR2_X1 U553 ( .A(G50GAT), .B(n491), .Z(G1331GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT106), .B(n533), .Z(n551) );
  NOR2_X1 U555 ( .A1(n567), .A2(n551), .ZN(n502) );
  NAND2_X1 U556 ( .A1(n502), .A2(n492), .ZN(n499) );
  NOR2_X1 U557 ( .A1(n505), .A2(n499), .ZN(n494) );
  XNOR2_X1 U558 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U560 ( .A(G57GAT), .B(n495), .ZN(G1332GAT) );
  NOR2_X1 U561 ( .A1(n509), .A2(n499), .ZN(n496) );
  XOR2_X1 U562 ( .A(KEYINPUT108), .B(n496), .Z(n497) );
  XNOR2_X1 U563 ( .A(G64GAT), .B(n497), .ZN(G1333GAT) );
  NOR2_X1 U564 ( .A1(n511), .A2(n499), .ZN(n498) );
  XOR2_X1 U565 ( .A(G71GAT), .B(n498), .Z(G1334GAT) );
  NOR2_X1 U566 ( .A1(n514), .A2(n499), .ZN(n501) );
  XNOR2_X1 U567 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n501), .B(n500), .ZN(G1335GAT) );
  INV_X1 U569 ( .A(G85GAT), .ZN(n507) );
  NAND2_X1 U570 ( .A1(n503), .A2(n502), .ZN(n504) );
  XOR2_X1 U571 ( .A(KEYINPUT109), .B(n504), .Z(n513) );
  NOR2_X1 U572 ( .A1(n505), .A2(n513), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT110), .B(n508), .ZN(G1336GAT) );
  NOR2_X1 U575 ( .A1(n509), .A2(n513), .ZN(n510) );
  XOR2_X1 U576 ( .A(G92GAT), .B(n510), .Z(G1337GAT) );
  NOR2_X1 U577 ( .A1(n511), .A2(n513), .ZN(n512) );
  XOR2_X1 U578 ( .A(G99GAT), .B(n512), .Z(G1338GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n515) );
  XOR2_X1 U580 ( .A(KEYINPUT44), .B(n515), .Z(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G106GAT), .ZN(G1339GAT) );
  NOR2_X1 U582 ( .A1(n528), .A2(n517), .ZN(n518) );
  NAND2_X1 U583 ( .A1(n548), .A2(n518), .ZN(n524) );
  NOR2_X1 U584 ( .A1(n549), .A2(n524), .ZN(n519) );
  XOR2_X1 U585 ( .A(G113GAT), .B(n519), .Z(G1340GAT) );
  NOR2_X1 U586 ( .A1(n551), .A2(n524), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1341GAT) );
  NOR2_X1 U589 ( .A1(n557), .A2(n524), .ZN(n522) );
  XOR2_X1 U590 ( .A(KEYINPUT50), .B(n522), .Z(n523) );
  XNOR2_X1 U591 ( .A(G127GAT), .B(n523), .ZN(G1342GAT) );
  NOR2_X1 U592 ( .A1(n564), .A2(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(G1343GAT) );
  NOR2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(KEYINPUT113), .B(n531), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n567), .A2(n540), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G141GAT), .B(n532), .ZN(G1344GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n535) );
  NAND2_X1 U601 ( .A1(n540), .A2(n533), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G148GAT), .B(n536), .ZN(G1345GAT) );
  NAND2_X1 U604 ( .A1(n540), .A2(n572), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n537), .B(KEYINPUT114), .ZN(n538) );
  XNOR2_X1 U606 ( .A(G155GAT), .B(n538), .ZN(G1346GAT) );
  XOR2_X1 U607 ( .A(G162GAT), .B(KEYINPUT115), .Z(n542) );
  INV_X1 U608 ( .A(n564), .ZN(n539) );
  NAND2_X1 U609 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1347GAT) );
  NOR2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U612 ( .A(KEYINPUT55), .B(KEYINPUT116), .ZN(n545) );
  XOR2_X1 U613 ( .A(n546), .B(n545), .Z(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n563) );
  NOR2_X1 U615 ( .A1(n549), .A2(n563), .ZN(n550) );
  XOR2_X1 U616 ( .A(G169GAT), .B(n550), .Z(G1348GAT) );
  NOR2_X1 U617 ( .A1(n563), .A2(n551), .ZN(n556) );
  XOR2_X1 U618 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n553) );
  XNOR2_X1 U619 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(KEYINPUT56), .B(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n563), .ZN(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(n560), .ZN(G1350GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n562) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n566) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(n566), .B(n565), .Z(G1351GAT) );
  NAND2_X1 U632 ( .A1(n576), .A2(n567), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n574) );
  NAND2_X1 U638 ( .A1(n576), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

