

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, n1034, G284, G297, G282, G295, n516, n517, n518,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U551 ( .A(n625), .Z(n664) );
  NOR2_X1 U552 ( .A1(n714), .A2(n701), .ZN(n703) );
  AND2_X1 U553 ( .A1(n692), .A2(n691), .ZN(n693) );
  OR2_X1 U554 ( .A1(n690), .A2(n689), .ZN(n691) );
  INV_X1 U555 ( .A(n625), .ZN(n660) );
  NAND2_X1 U556 ( .A1(G8), .A2(n625), .ZN(n714) );
  NAND2_X1 U557 ( .A1(n609), .A2(n608), .ZN(n625) );
  BUF_X1 U558 ( .A(n533), .Z(n720) );
  INV_X1 U559 ( .A(G2104), .ZN(n526) );
  NAND2_X1 U560 ( .A1(n517), .A2(n518), .ZN(n516) );
  NAND2_X1 U561 ( .A1(n705), .A2(n704), .ZN(n517) );
  AND2_X1 U562 ( .A1(n521), .A2(n992), .ZN(n518) );
  NOR2_X1 U563 ( .A1(n542), .A2(n541), .ZN(G160) );
  NOR2_X1 U564 ( .A1(n542), .A2(n541), .ZN(n1034) );
  AND2_X1 U565 ( .A1(n716), .A2(n715), .ZN(n520) );
  OR2_X1 U566 ( .A1(n707), .A2(n714), .ZN(n521) );
  INV_X1 U567 ( .A(KEYINPUT92), .ZN(n636) );
  INV_X1 U568 ( .A(KEYINPUT28), .ZN(n653) );
  XNOR2_X1 U569 ( .A(n657), .B(KEYINPUT29), .ZN(n658) );
  XNOR2_X1 U570 ( .A(KEYINPUT32), .B(KEYINPUT96), .ZN(n695) );
  INV_X1 U571 ( .A(KEYINPUT64), .ZN(n702) );
  AND2_X2 U572 ( .A1(n526), .A2(G2105), .ZN(n876) );
  NOR2_X1 U573 ( .A1(n719), .A2(n718), .ZN(n744) );
  NOR2_X1 U574 ( .A1(G651), .A2(n581), .ZN(n791) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n875) );
  NAND2_X1 U576 ( .A1(G114), .A2(n875), .ZN(n523) );
  NAND2_X1 U577 ( .A1(G126), .A2(n876), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U579 ( .A(KEYINPUT80), .B(n524), .ZN(n530) );
  NOR2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XOR2_X1 U581 ( .A(KEYINPUT17), .B(n525), .Z(n538) );
  BUF_X1 U582 ( .A(n538), .Z(n879) );
  NAND2_X1 U583 ( .A1(G138), .A2(n879), .ZN(n528) );
  NOR2_X1 U584 ( .A1(G2105), .A2(n526), .ZN(n533) );
  NAND2_X1 U585 ( .A1(G102), .A2(n720), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U587 ( .A1(n530), .A2(n529), .ZN(G164) );
  INV_X1 U588 ( .A(KEYINPUT66), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n876), .A2(G125), .ZN(n531) );
  XNOR2_X1 U590 ( .A(n532), .B(n531), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n533), .A2(G101), .ZN(n534) );
  XNOR2_X1 U592 ( .A(KEYINPUT23), .B(n534), .ZN(n535) );
  NOR2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U594 ( .A(n537), .B(KEYINPUT67), .ZN(n542) );
  NAND2_X1 U595 ( .A1(G113), .A2(n875), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G137), .A2(n538), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U598 ( .A(G543), .B(KEYINPUT0), .Z(n581) );
  NAND2_X1 U599 ( .A1(G53), .A2(n791), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT70), .B(n543), .Z(n550) );
  NOR2_X1 U601 ( .A1(G543), .A2(G651), .ZN(n544) );
  XOR2_X2 U602 ( .A(KEYINPUT65), .B(n544), .Z(n797) );
  NAND2_X1 U603 ( .A1(G91), .A2(n797), .ZN(n547) );
  INV_X1 U604 ( .A(G651), .ZN(n551) );
  OR2_X1 U605 ( .A1(n551), .A2(n581), .ZN(n545) );
  XOR2_X2 U606 ( .A(KEYINPUT68), .B(n545), .Z(n794) );
  NAND2_X1 U607 ( .A1(G78), .A2(n794), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U609 ( .A(KEYINPUT69), .B(n548), .Z(n549) );
  NOR2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n554) );
  NOR2_X1 U611 ( .A1(G543), .A2(n551), .ZN(n552) );
  XOR2_X2 U612 ( .A(KEYINPUT1), .B(n552), .Z(n793) );
  NAND2_X1 U613 ( .A1(n793), .A2(G65), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(G299) );
  NAND2_X1 U615 ( .A1(G52), .A2(n791), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G64), .A2(n793), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G90), .A2(n797), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G77), .A2(n794), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n559), .Z(n560) );
  NOR2_X1 U622 ( .A1(n561), .A2(n560), .ZN(G171) );
  INV_X1 U623 ( .A(G171), .ZN(G301) );
  NAND2_X1 U624 ( .A1(n797), .A2(G89), .ZN(n562) );
  XNOR2_X1 U625 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G76), .A2(n794), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U629 ( .A1(G51), .A2(n791), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G63), .A2(n793), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U634 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U635 ( .A1(G88), .A2(n797), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G75), .A2(n794), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G50), .A2(n791), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G62), .A2(n793), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(G166) );
  XNOR2_X1 U642 ( .A(KEYINPUT81), .B(G166), .ZN(G303) );
  XOR2_X1 U643 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U644 ( .A1(G49), .A2(n791), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G74), .A2(G651), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U647 ( .A1(n793), .A2(n580), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n581), .A2(G87), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(G288) );
  NAND2_X1 U650 ( .A1(G86), .A2(n797), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G48), .A2(n791), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n794), .A2(G73), .ZN(n586) );
  XOR2_X1 U654 ( .A(KEYINPUT2), .B(n586), .Z(n587) );
  NOR2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n793), .A2(G61), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(G305) );
  AND2_X1 U658 ( .A1(G72), .A2(n794), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G85), .A2(n797), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G47), .A2(n791), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n793), .A2(G60), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n596), .A2(n595), .ZN(G290) );
  NOR2_X1 U665 ( .A1(G164), .A2(G1384), .ZN(n608) );
  NAND2_X1 U666 ( .A1(n1034), .A2(G40), .ZN(n607) );
  NOR2_X1 U667 ( .A1(n608), .A2(n607), .ZN(n757) );
  XNOR2_X1 U668 ( .A(KEYINPUT82), .B(KEYINPUT34), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G140), .A2(n879), .ZN(n598) );
  NAND2_X1 U670 ( .A1(G104), .A2(n720), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n600), .B(n599), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G116), .A2(n875), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G128), .A2(n876), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U676 ( .A(KEYINPUT35), .B(n603), .Z(n604) );
  NOR2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U678 ( .A(KEYINPUT36), .B(n606), .Z(n895) );
  XOR2_X1 U679 ( .A(G2067), .B(KEYINPUT37), .Z(n753) );
  AND2_X1 U680 ( .A1(n895), .A2(n753), .ZN(n954) );
  NAND2_X1 U681 ( .A1(n757), .A2(n954), .ZN(n751) );
  INV_X1 U682 ( .A(n751), .ZN(n719) );
  XNOR2_X1 U683 ( .A(KEYINPUT89), .B(n607), .ZN(n609) );
  NOR2_X1 U684 ( .A1(G1966), .A2(n714), .ZN(n673) );
  NAND2_X1 U685 ( .A1(G1996), .A2(n660), .ZN(n610) );
  XNOR2_X1 U686 ( .A(n610), .B(KEYINPUT26), .ZN(n628) );
  NAND2_X1 U687 ( .A1(n793), .A2(G56), .ZN(n611) );
  XOR2_X1 U688 ( .A(KEYINPUT14), .B(n611), .Z(n613) );
  AND2_X1 U689 ( .A1(G43), .A2(n791), .ZN(n612) );
  NOR2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n623) );
  NAND2_X1 U691 ( .A1(n797), .A2(G81), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT12), .ZN(n616) );
  NAND2_X1 U693 ( .A1(G68), .A2(n794), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n617), .A2(KEYINPUT13), .ZN(n621) );
  INV_X1 U696 ( .A(n617), .ZN(n619) );
  INV_X1 U697 ( .A(KEYINPUT13), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n622) );
  AND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U701 ( .A(KEYINPUT73), .B(n624), .Z(n766) );
  NAND2_X1 U702 ( .A1(G1341), .A2(n664), .ZN(n626) );
  AND2_X1 U703 ( .A1(n766), .A2(n626), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n642) );
  NAND2_X1 U705 ( .A1(G54), .A2(n791), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G66), .A2(n793), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U708 ( .A1(G92), .A2(n797), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G79), .A2(n794), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U712 ( .A(n635), .B(KEYINPUT15), .Z(n983) );
  INV_X1 U713 ( .A(n983), .ZN(n773) );
  NOR2_X1 U714 ( .A1(n642), .A2(n773), .ZN(n637) );
  XNOR2_X1 U715 ( .A(n637), .B(n636), .ZN(n641) );
  NOR2_X1 U716 ( .A1(n660), .A2(G1348), .ZN(n639) );
  NOR2_X1 U717 ( .A1(G2067), .A2(n664), .ZN(n638) );
  NOR2_X1 U718 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n642), .A2(n773), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n651) );
  INV_X1 U722 ( .A(G299), .ZN(n808) );
  XOR2_X1 U723 ( .A(KEYINPUT90), .B(KEYINPUT27), .Z(n646) );
  NAND2_X1 U724 ( .A1(n660), .A2(G2072), .ZN(n645) );
  XOR2_X1 U725 ( .A(n646), .B(n645), .Z(n649) );
  NAND2_X1 U726 ( .A1(G1956), .A2(n664), .ZN(n647) );
  XNOR2_X1 U727 ( .A(n647), .B(KEYINPUT91), .ZN(n648) );
  NOR2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n808), .A2(n652), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n656) );
  NOR2_X1 U731 ( .A1(n808), .A2(n652), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n659) );
  XOR2_X1 U734 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n657) );
  XNOR2_X1 U735 ( .A(n659), .B(n658), .ZN(n688) );
  XOR2_X1 U736 ( .A(KEYINPUT25), .B(G2078), .Z(n927) );
  NOR2_X1 U737 ( .A1(n927), .A2(n664), .ZN(n662) );
  NOR2_X1 U738 ( .A1(n660), .A2(G1961), .ZN(n661) );
  NOR2_X1 U739 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U740 ( .A1(G301), .A2(n663), .ZN(n686) );
  NOR2_X1 U741 ( .A1(n688), .A2(n686), .ZN(n671) );
  AND2_X1 U742 ( .A1(G301), .A2(n663), .ZN(n669) );
  NOR2_X1 U743 ( .A1(G2084), .A2(n664), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n673), .A2(n676), .ZN(n665) );
  NAND2_X1 U745 ( .A1(G8), .A2(n665), .ZN(n666) );
  XNOR2_X1 U746 ( .A(KEYINPUT30), .B(n666), .ZN(n667) );
  NOR2_X1 U747 ( .A1(G168), .A2(n667), .ZN(n668) );
  NOR2_X1 U748 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U749 ( .A(n670), .B(KEYINPUT31), .ZN(n690) );
  NOR2_X1 U750 ( .A1(n671), .A2(n690), .ZN(n672) );
  NOR2_X1 U751 ( .A1(n673), .A2(n672), .ZN(n675) );
  INV_X1 U752 ( .A(KEYINPUT95), .ZN(n674) );
  XNOR2_X1 U753 ( .A(n675), .B(n674), .ZN(n678) );
  NAND2_X1 U754 ( .A1(n676), .A2(G8), .ZN(n677) );
  NAND2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n698) );
  INV_X1 U756 ( .A(G8), .ZN(n683) );
  NOR2_X1 U757 ( .A1(G1971), .A2(n714), .ZN(n680) );
  NOR2_X1 U758 ( .A1(G2090), .A2(n664), .ZN(n679) );
  NOR2_X1 U759 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U760 ( .A1(n681), .A2(G303), .ZN(n682) );
  NOR2_X1 U761 ( .A1(n683), .A2(n682), .ZN(n689) );
  AND2_X1 U762 ( .A1(G286), .A2(G8), .ZN(n684) );
  OR2_X1 U763 ( .A1(n689), .A2(n684), .ZN(n692) );
  INV_X1 U764 ( .A(n692), .ZN(n685) );
  OR2_X1 U765 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U766 ( .A1(n688), .A2(n687), .ZN(n694) );
  NOR2_X1 U767 ( .A1(n694), .A2(n693), .ZN(n696) );
  XNOR2_X1 U768 ( .A(n696), .B(n695), .ZN(n697) );
  NAND2_X1 U769 ( .A1(n698), .A2(n697), .ZN(n708) );
  NOR2_X1 U770 ( .A1(G1976), .A2(G288), .ZN(n706) );
  NOR2_X1 U771 ( .A1(G1971), .A2(G303), .ZN(n699) );
  NOR2_X1 U772 ( .A1(n706), .A2(n699), .ZN(n981) );
  NAND2_X1 U773 ( .A1(n708), .A2(n981), .ZN(n700) );
  NAND2_X1 U774 ( .A1(G1976), .A2(G288), .ZN(n977) );
  NAND2_X1 U775 ( .A1(n700), .A2(n977), .ZN(n701) );
  XNOR2_X1 U776 ( .A(n703), .B(n702), .ZN(n705) );
  INV_X1 U777 ( .A(KEYINPUT33), .ZN(n704) );
  NAND2_X1 U778 ( .A1(n706), .A2(KEYINPUT33), .ZN(n707) );
  XOR2_X1 U779 ( .A(G1981), .B(G305), .Z(n992) );
  NOR2_X1 U780 ( .A1(G2090), .A2(G303), .ZN(n709) );
  NAND2_X1 U781 ( .A1(G8), .A2(n709), .ZN(n710) );
  NAND2_X1 U782 ( .A1(n708), .A2(n710), .ZN(n711) );
  NAND2_X1 U783 ( .A1(n711), .A2(n714), .ZN(n716) );
  NOR2_X1 U784 ( .A1(G1981), .A2(G305), .ZN(n712) );
  XOR2_X1 U785 ( .A(n712), .B(KEYINPUT24), .Z(n713) );
  OR2_X1 U786 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U787 ( .A1(n516), .A2(n520), .ZN(n717) );
  XNOR2_X1 U788 ( .A(n717), .B(KEYINPUT97), .ZN(n718) );
  NAND2_X1 U789 ( .A1(G105), .A2(n720), .ZN(n721) );
  XNOR2_X1 U790 ( .A(n721), .B(KEYINPUT38), .ZN(n722) );
  XNOR2_X1 U791 ( .A(n722), .B(KEYINPUT86), .ZN(n724) );
  NAND2_X1 U792 ( .A1(G129), .A2(n876), .ZN(n723) );
  NAND2_X1 U793 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U794 ( .A1(G141), .A2(n879), .ZN(n725) );
  XNOR2_X1 U795 ( .A(KEYINPUT87), .B(n725), .ZN(n726) );
  NOR2_X1 U796 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U797 ( .A1(G117), .A2(n875), .ZN(n728) );
  XOR2_X1 U798 ( .A(KEYINPUT85), .B(n728), .Z(n729) );
  NAND2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n891) );
  NAND2_X1 U800 ( .A1(G1996), .A2(n891), .ZN(n731) );
  XOR2_X1 U801 ( .A(KEYINPUT88), .B(n731), .Z(n741) );
  INV_X1 U802 ( .A(G1991), .ZN(n838) );
  NAND2_X1 U803 ( .A1(G119), .A2(n876), .ZN(n733) );
  NAND2_X1 U804 ( .A1(G95), .A2(n720), .ZN(n732) );
  NAND2_X1 U805 ( .A1(n733), .A2(n732), .ZN(n739) );
  NAND2_X1 U806 ( .A1(G131), .A2(n879), .ZN(n734) );
  XNOR2_X1 U807 ( .A(n734), .B(KEYINPUT84), .ZN(n737) );
  NAND2_X1 U808 ( .A1(G107), .A2(n875), .ZN(n735) );
  XOR2_X1 U809 ( .A(KEYINPUT83), .B(n735), .Z(n736) );
  NAND2_X1 U810 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U811 ( .A1(n739), .A2(n738), .ZN(n887) );
  NOR2_X1 U812 ( .A1(n838), .A2(n887), .ZN(n740) );
  NOR2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n745) );
  XOR2_X1 U814 ( .A(G1986), .B(G290), .Z(n978) );
  NAND2_X1 U815 ( .A1(n745), .A2(n978), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n742), .A2(n757), .ZN(n743) );
  NAND2_X1 U817 ( .A1(n744), .A2(n743), .ZN(n760) );
  NOR2_X1 U818 ( .A1(G1996), .A2(n891), .ZN(n949) );
  INV_X1 U819 ( .A(n745), .ZN(n961) );
  AND2_X1 U820 ( .A1(n887), .A2(n838), .ZN(n746) );
  XNOR2_X1 U821 ( .A(n746), .B(KEYINPUT98), .ZN(n945) );
  NOR2_X1 U822 ( .A1(G1986), .A2(G290), .ZN(n747) );
  NOR2_X1 U823 ( .A1(n945), .A2(n747), .ZN(n748) );
  NOR2_X1 U824 ( .A1(n961), .A2(n748), .ZN(n749) );
  NOR2_X1 U825 ( .A1(n949), .A2(n749), .ZN(n750) );
  XNOR2_X1 U826 ( .A(n750), .B(KEYINPUT39), .ZN(n752) );
  NAND2_X1 U827 ( .A1(n752), .A2(n751), .ZN(n755) );
  NOR2_X1 U828 ( .A1(n753), .A2(n895), .ZN(n754) );
  XNOR2_X1 U829 ( .A(n754), .B(KEYINPUT99), .ZN(n966) );
  NAND2_X1 U830 ( .A1(n755), .A2(n966), .ZN(n756) );
  XNOR2_X1 U831 ( .A(KEYINPUT100), .B(n756), .ZN(n758) );
  NAND2_X1 U832 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U833 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U834 ( .A(n761), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U835 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U836 ( .A(G132), .ZN(G219) );
  INV_X1 U837 ( .A(G82), .ZN(G220) );
  INV_X1 U838 ( .A(G57), .ZN(G237) );
  INV_X1 U839 ( .A(G108), .ZN(G238) );
  INV_X1 U840 ( .A(G69), .ZN(G235) );
  XOR2_X1 U841 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n765) );
  XOR2_X1 U842 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n763) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n762) );
  XOR2_X1 U844 ( .A(n763), .B(n762), .Z(n921) );
  NAND2_X1 U845 ( .A1(G567), .A2(n921), .ZN(n764) );
  XNOR2_X1 U846 ( .A(n765), .B(n764), .ZN(G234) );
  BUF_X1 U847 ( .A(n766), .Z(n989) );
  NAND2_X1 U848 ( .A1(n989), .A2(G860), .ZN(G153) );
  NAND2_X1 U849 ( .A1(G868), .A2(G301), .ZN(n768) );
  INV_X1 U850 ( .A(G868), .ZN(n814) );
  NAND2_X1 U851 ( .A1(n773), .A2(n814), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n768), .A2(n767), .ZN(G284) );
  NOR2_X1 U853 ( .A1(G868), .A2(G299), .ZN(n770) );
  NOR2_X1 U854 ( .A1(G286), .A2(n814), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U856 ( .A(KEYINPUT74), .B(n771), .ZN(G297) );
  INV_X1 U857 ( .A(G559), .ZN(n775) );
  NOR2_X1 U858 ( .A1(G860), .A2(n775), .ZN(n772) );
  NOR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U860 ( .A(KEYINPUT16), .B(n774), .Z(G148) );
  NAND2_X1 U861 ( .A1(n775), .A2(n983), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n776), .A2(G868), .ZN(n779) );
  INV_X1 U863 ( .A(n989), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n777), .A2(n814), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(G282) );
  NAND2_X1 U866 ( .A1(G123), .A2(n876), .ZN(n780) );
  XOR2_X1 U867 ( .A(KEYINPUT75), .B(n780), .Z(n781) );
  XNOR2_X1 U868 ( .A(n781), .B(KEYINPUT18), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G111), .A2(n875), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G135), .A2(n879), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G99), .A2(n720), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n946) );
  XNOR2_X1 U875 ( .A(n946), .B(G2096), .ZN(n788) );
  INV_X1 U876 ( .A(G2100), .ZN(n855) );
  NAND2_X1 U877 ( .A1(n788), .A2(n855), .ZN(G156) );
  NAND2_X1 U878 ( .A1(G559), .A2(n983), .ZN(n789) );
  XOR2_X1 U879 ( .A(KEYINPUT76), .B(n789), .Z(n811) );
  XNOR2_X1 U880 ( .A(n811), .B(n989), .ZN(n790) );
  NOR2_X1 U881 ( .A1(G860), .A2(n790), .ZN(n803) );
  NAND2_X1 U882 ( .A1(G55), .A2(n791), .ZN(n792) );
  XNOR2_X1 U883 ( .A(n792), .B(KEYINPUT78), .ZN(n802) );
  NAND2_X1 U884 ( .A1(n793), .A2(G67), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G80), .A2(n794), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G93), .A2(n797), .ZN(n798) );
  XNOR2_X1 U888 ( .A(KEYINPUT77), .B(n798), .ZN(n799) );
  NOR2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n813) );
  XOR2_X1 U891 ( .A(n803), .B(n813), .Z(G145) );
  XNOR2_X1 U892 ( .A(KEYINPUT19), .B(G288), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n804), .B(n813), .ZN(n807) );
  XNOR2_X1 U894 ( .A(G166), .B(G290), .ZN(n805) );
  XNOR2_X1 U895 ( .A(n805), .B(G305), .ZN(n806) );
  XNOR2_X1 U896 ( .A(n807), .B(n806), .ZN(n810) );
  XOR2_X1 U897 ( .A(n989), .B(n808), .Z(n809) );
  XNOR2_X1 U898 ( .A(n810), .B(n809), .ZN(n899) );
  XNOR2_X1 U899 ( .A(n811), .B(n899), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n812), .A2(G868), .ZN(n816) );
  NAND2_X1 U901 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U902 ( .A1(n816), .A2(n815), .ZN(G295) );
  NAND2_X1 U903 ( .A1(G2078), .A2(G2084), .ZN(n817) );
  XOR2_X1 U904 ( .A(KEYINPUT20), .B(n817), .Z(n818) );
  NAND2_X1 U905 ( .A1(G2090), .A2(n818), .ZN(n819) );
  XNOR2_X1 U906 ( .A(KEYINPUT21), .B(n819), .ZN(n820) );
  NAND2_X1 U907 ( .A1(n820), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U908 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U909 ( .A1(G235), .A2(G238), .ZN(n821) );
  NAND2_X1 U910 ( .A1(G120), .A2(n821), .ZN(n822) );
  NOR2_X1 U911 ( .A1(n822), .A2(G237), .ZN(n823) );
  XNOR2_X1 U912 ( .A(n823), .B(KEYINPUT79), .ZN(n835) );
  NAND2_X1 U913 ( .A1(n835), .A2(G567), .ZN(n828) );
  NOR2_X1 U914 ( .A1(G220), .A2(G219), .ZN(n824) );
  XOR2_X1 U915 ( .A(KEYINPUT22), .B(n824), .Z(n825) );
  NOR2_X1 U916 ( .A1(G218), .A2(n825), .ZN(n826) );
  NAND2_X1 U917 ( .A1(G96), .A2(n826), .ZN(n834) );
  NAND2_X1 U918 ( .A1(n834), .A2(G2106), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(n837) );
  NAND2_X1 U920 ( .A1(G661), .A2(G483), .ZN(n829) );
  NOR2_X1 U921 ( .A1(n837), .A2(n829), .ZN(n833) );
  NAND2_X1 U922 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(n921), .A2(G2106), .ZN(n830) );
  XOR2_X1 U924 ( .A(KEYINPUT103), .B(n830), .Z(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U926 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  XOR2_X1 U929 ( .A(G120), .B(KEYINPUT104), .Z(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U933 ( .A(n836), .B(KEYINPUT105), .Z(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n837), .ZN(G319) );
  XNOR2_X1 U936 ( .A(G1996), .B(G2474), .ZN(n848) );
  XOR2_X1 U937 ( .A(G1976), .B(G1956), .Z(n840) );
  XOR2_X1 U938 ( .A(n838), .B(G1971), .Z(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U940 ( .A(G1981), .B(G1966), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1961), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U944 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(G229) );
  XOR2_X1 U947 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n850) );
  XNOR2_X1 U948 ( .A(G2678), .B(KEYINPUT43), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U950 ( .A(KEYINPUT42), .B(G2072), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U953 ( .A(n854), .B(n853), .Z(n857) );
  XOR2_X1 U954 ( .A(G2096), .B(n855), .Z(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n859) );
  XOR2_X1 U956 ( .A(G2078), .B(G2084), .Z(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(G227) );
  NAND2_X1 U958 ( .A1(G124), .A2(n876), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U960 ( .A1(n875), .A2(G112), .ZN(n861) );
  NAND2_X1 U961 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U962 ( .A1(G136), .A2(n879), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G100), .A2(n720), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U965 ( .A1(n866), .A2(n865), .ZN(G162) );
  NAND2_X1 U966 ( .A1(G139), .A2(n879), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G103), .A2(n720), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U969 ( .A1(G115), .A2(n875), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G127), .A2(n876), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U972 ( .A(KEYINPUT47), .B(n871), .ZN(n872) );
  XNOR2_X1 U973 ( .A(KEYINPUT109), .B(n872), .ZN(n873) );
  NOR2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n955) );
  XNOR2_X1 U975 ( .A(n955), .B(G162), .ZN(n886) );
  NAND2_X1 U976 ( .A1(G118), .A2(n875), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G130), .A2(n876), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G142), .A2(n879), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G106), .A2(n720), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n882), .Z(n883) );
  NOR2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n888) );
  XOR2_X1 U985 ( .A(n888), .B(n887), .Z(n890) );
  XNOR2_X1 U986 ( .A(G164), .B(G160), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n897) );
  XNOR2_X1 U988 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n891), .B(n946), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U991 ( .A(n895), .B(n894), .Z(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U993 ( .A1(G37), .A2(n898), .ZN(G395) );
  XOR2_X1 U994 ( .A(KEYINPUT110), .B(n899), .Z(n901) );
  XOR2_X1 U995 ( .A(G301), .B(n983), .Z(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U997 ( .A(G286), .B(n902), .Z(n903) );
  NOR2_X1 U998 ( .A1(G37), .A2(n903), .ZN(G397) );
  XNOR2_X1 U999 ( .A(G2451), .B(G2427), .ZN(n913) );
  XOR2_X1 U1000 ( .A(KEYINPUT101), .B(G2443), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G2435), .B(G2438), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1003 ( .A(G2454), .B(G2430), .Z(n907) );
  XNOR2_X1 U1004 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1006 ( .A(n909), .B(n908), .Z(n911) );
  XNOR2_X1 U1007 ( .A(G2446), .B(KEYINPUT102), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n914), .A2(G14), .ZN(n920) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n920), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(n920), .ZN(G401) );
  INV_X1 U1019 ( .A(n921), .ZN(G223) );
  XOR2_X1 U1020 ( .A(KEYINPUT55), .B(KEYINPUT115), .Z(n941) );
  XNOR2_X1 U1021 ( .A(G2090), .B(G35), .ZN(n936) );
  XOR2_X1 U1022 ( .A(G25), .B(G1991), .Z(n922) );
  NAND2_X1 U1023 ( .A1(n922), .A2(G28), .ZN(n933) );
  XOR2_X1 U1024 ( .A(G2067), .B(G26), .Z(n923) );
  XNOR2_X1 U1025 ( .A(KEYINPUT113), .B(n923), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(G33), .B(G2072), .ZN(n924) );
  NOR2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(KEYINPUT114), .B(n926), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G1996), .B(G32), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n927), .B(G27), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(KEYINPUT53), .B(n934), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1036 ( .A(G2084), .B(G34), .Z(n937) );
  XNOR2_X1 U1037 ( .A(KEYINPUT54), .B(n937), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(n941), .B(n940), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(G29), .A2(n942), .ZN(n943) );
  XOR2_X1 U1041 ( .A(KEYINPUT116), .B(n943), .Z(n944) );
  NAND2_X1 U1042 ( .A1(G11), .A2(n944), .ZN(n973) );
  INV_X1 U1043 ( .A(G29), .ZN(n971) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G2090), .B(G162), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(n947), .B(KEYINPUT111), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1048 ( .A(KEYINPUT51), .B(n950), .Z(n951) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n965) );
  XOR2_X1 U1050 ( .A(G160), .B(G2084), .Z(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n963) );
  XOR2_X1 U1052 ( .A(G164), .B(G2078), .Z(n958) );
  XOR2_X1 U1053 ( .A(n955), .B(KEYINPUT112), .Z(n956) );
  XNOR2_X1 U1054 ( .A(G2072), .B(n956), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1056 ( .A(KEYINPUT50), .B(n959), .Z(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT52), .B(n968), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(KEYINPUT55), .A2(n969), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n1000) );
  XNOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .ZN(n998) );
  XOR2_X1 U1066 ( .A(G301), .B(G1961), .Z(n974) );
  XNOR2_X1 U1067 ( .A(n974), .B(KEYINPUT118), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(G1971), .A2(G303), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n988) );
  XOR2_X1 U1072 ( .A(G299), .B(G1956), .Z(n982) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G1348), .B(n983), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT117), .B(n984), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1078 ( .A(G1341), .B(n989), .Z(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n996) );
  XNOR2_X1 U1080 ( .A(G168), .B(G1966), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(n994), .B(KEYINPUT57), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1032) );
  XOR2_X1 U1086 ( .A(G16), .B(KEYINPUT119), .Z(n1029) );
  XOR2_X1 U1087 ( .A(G1986), .B(G24), .Z(n1004) );
  XNOR2_X1 U1088 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G23), .B(G1976), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(KEYINPUT58), .B(n1005), .ZN(n1025) );
  XNOR2_X1 U1093 ( .A(KEYINPUT121), .B(G1341), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(n1006), .B(G19), .ZN(n1013) );
  XOR2_X1 U1095 ( .A(KEYINPUT123), .B(G4), .Z(n1008) );
  XNOR2_X1 U1096 ( .A(G1348), .B(KEYINPUT59), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1008), .B(n1007), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(KEYINPUT122), .B(n1009), .Z(n1011) );
  XNOR2_X1 U1099 ( .A(G1981), .B(G6), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT120), .B(G1956), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(G20), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT124), .B(n1017), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(n1018), .B(KEYINPUT60), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(G1961), .B(G5), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(G21), .B(G1966), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1111 ( .A(n1023), .B(KEYINPUT125), .Z(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1113 ( .A(KEYINPUT126), .B(n1026), .Z(n1027) );
  XNOR2_X1 U1114 ( .A(n1027), .B(KEYINPUT61), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1116 ( .A(KEYINPUT127), .B(n1030), .Z(n1031) );
  NOR2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1033), .Z(G150) );
  INV_X1 U1119 ( .A(G150), .ZN(G311) );
endmodule

