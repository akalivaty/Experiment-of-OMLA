

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n601), .A2(n571), .ZN(n816) );
  AND2_X1 U556 ( .A1(n551), .A2(G2104), .ZN(n1028) );
  NOR2_X1 U557 ( .A1(G651), .A2(n601), .ZN(n820) );
  NAND2_X2 U558 ( .A1(n629), .A2(G8), .ZN(n743) );
  OR2_X1 U559 ( .A1(n665), .A2(n986), .ZN(n666) );
  OR2_X1 U560 ( .A1(n663), .A2(n662), .ZN(n667) );
  NOR2_X2 U561 ( .A1(n551), .A2(G2104), .ZN(n1023) );
  NOR2_X2 U562 ( .A1(G651), .A2(G543), .ZN(n815) );
  NOR2_X2 U563 ( .A1(G2105), .A2(G2104), .ZN(n554) );
  NOR2_X1 U564 ( .A1(n743), .A2(G1966), .ZN(n689) );
  XNOR2_X1 U565 ( .A(n539), .B(KEYINPUT32), .ZN(n694) );
  NAND2_X1 U566 ( .A1(n535), .A2(n532), .ZN(n539) );
  NAND2_X1 U567 ( .A1(n534), .A2(n533), .ZN(n532) );
  AND2_X1 U568 ( .A1(n537), .A2(n522), .ZN(n535) );
  INV_X1 U569 ( .A(KEYINPUT33), .ZN(n544) );
  XNOR2_X1 U570 ( .A(n676), .B(n527), .ZN(n526) );
  INV_X1 U571 ( .A(KEYINPUT28), .ZN(n527) );
  OR2_X1 U572 ( .A1(n685), .A2(KEYINPUT94), .ZN(n536) );
  INV_X1 U573 ( .A(KEYINPUT94), .ZN(n533) );
  INV_X1 U574 ( .A(KEYINPUT64), .ZN(n529) );
  INV_X1 U575 ( .A(KEYINPUT95), .ZN(n695) );
  NAND2_X1 U576 ( .A1(n543), .A2(n523), .ZN(n753) );
  NAND2_X1 U577 ( .A1(n545), .A2(n544), .ZN(n543) );
  XNOR2_X1 U578 ( .A(n542), .B(n541), .ZN(n540) );
  INV_X1 U579 ( .A(KEYINPUT65), .ZN(n541) );
  XNOR2_X1 U580 ( .A(n560), .B(n559), .ZN(n561) );
  INV_X1 U581 ( .A(KEYINPUT23), .ZN(n559) );
  INV_X1 U582 ( .A(n629), .ZN(n669) );
  AND2_X1 U583 ( .A1(n536), .A2(G8), .ZN(n522) );
  NOR2_X1 U584 ( .A1(n737), .A2(n738), .ZN(n523) );
  NAND2_X1 U585 ( .A1(n524), .A2(n679), .ZN(n680) );
  XNOR2_X1 U586 ( .A(n525), .B(n677), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n528), .A2(n526), .ZN(n525) );
  NAND2_X1 U588 ( .A1(n673), .A2(n672), .ZN(n528) );
  XNOR2_X2 U589 ( .A(n530), .B(n529), .ZN(n629) );
  NOR2_X2 U590 ( .A1(n722), .A2(n531), .ZN(n530) );
  INV_X1 U591 ( .A(n723), .ZN(n531) );
  NAND2_X1 U592 ( .A1(G160), .A2(G40), .ZN(n722) );
  INV_X1 U593 ( .A(n686), .ZN(n534) );
  NAND2_X1 U594 ( .A1(n686), .A2(n538), .ZN(n537) );
  AND2_X1 U595 ( .A1(n685), .A2(KEYINPUT94), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n561), .A2(n540), .ZN(n565) );
  NAND2_X1 U597 ( .A1(n1027), .A2(G137), .ZN(n542) );
  XNOR2_X2 U598 ( .A(n554), .B(n553), .ZN(n1027) );
  NAND2_X1 U599 ( .A1(n702), .A2(n701), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n669), .A2(n782), .ZN(n659) );
  OR2_X1 U601 ( .A1(n990), .A2(n919), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n752), .A2(n751), .ZN(n547) );
  AND2_X1 U603 ( .A1(G8), .A2(n624), .ZN(n548) );
  INV_X1 U604 ( .A(KEYINPUT90), .ZN(n658) );
  INV_X1 U605 ( .A(KEYINPUT29), .ZN(n677) );
  INV_X1 U606 ( .A(n929), .ZN(n700) );
  NOR2_X1 U607 ( .A1(n700), .A2(n743), .ZN(n701) );
  INV_X1 U608 ( .A(KEYINPUT13), .ZN(n644) );
  INV_X1 U609 ( .A(KEYINPUT97), .ZN(n754) );
  XNOR2_X1 U610 ( .A(n645), .B(n644), .ZN(n646) );
  INV_X1 U611 ( .A(KEYINPUT17), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n650), .A2(n649), .ZN(n990) );
  INV_X1 U613 ( .A(G2105), .ZN(n551) );
  NAND2_X1 U614 ( .A1(G102), .A2(n1028), .ZN(n550) );
  AND2_X1 U615 ( .A1(G2105), .A2(G2104), .ZN(n1024) );
  NAND2_X1 U616 ( .A1(G114), .A2(n1024), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n1023), .A2(G126), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(KEYINPUT84), .ZN(n556) );
  NAND2_X1 U620 ( .A1(G138), .A2(n1027), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X2 U622 ( .A1(n558), .A2(n557), .ZN(G164) );
  NAND2_X1 U623 ( .A1(G101), .A2(n1028), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G125), .A2(n1023), .ZN(n563) );
  NAND2_X1 U625 ( .A1(G113), .A2(n1024), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X2 U627 ( .A1(n565), .A2(n564), .ZN(G160) );
  INV_X1 U628 ( .A(G651), .ZN(n571) );
  NOR2_X1 U629 ( .A1(G543), .A2(n571), .ZN(n566) );
  XOR2_X2 U630 ( .A(KEYINPUT1), .B(n566), .Z(n819) );
  NAND2_X1 U631 ( .A1(G63), .A2(n819), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT0), .B(G543), .Z(n601) );
  NAND2_X1 U633 ( .A1(G51), .A2(n820), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT6), .B(n569), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n815), .A2(G89), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G76), .A2(n816), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT5), .B(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT71), .B(n575), .ZN(n576) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT7), .B(n578), .Z(G168) );
  XOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U645 ( .A1(n815), .A2(G90), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT67), .B(n579), .Z(n581) );
  NAND2_X1 U647 ( .A1(n816), .A2(G77), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U649 ( .A(KEYINPUT9), .B(n582), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G64), .A2(n819), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G52), .A2(n820), .ZN(n583) );
  AND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(G301) );
  INV_X1 U654 ( .A(G301), .ZN(G171) );
  NAND2_X1 U655 ( .A1(G91), .A2(n815), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G65), .A2(n819), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U658 ( .A1(n816), .A2(G78), .ZN(n589) );
  XOR2_X1 U659 ( .A(KEYINPUT68), .B(n589), .Z(n590) );
  NOR2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U661 ( .A1(n820), .A2(G53), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n593), .A2(n592), .ZN(G299) );
  NAND2_X1 U663 ( .A1(n816), .A2(G75), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G88), .A2(n815), .ZN(n594) );
  XOR2_X1 U665 ( .A(KEYINPUT79), .B(n594), .Z(n595) );
  NAND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G62), .A2(n819), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G50), .A2(n820), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U670 ( .A1(n600), .A2(n599), .ZN(G166) );
  INV_X1 U671 ( .A(G166), .ZN(G303) );
  NAND2_X1 U672 ( .A1(n601), .A2(G87), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G49), .A2(n820), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G74), .A2(G651), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U676 ( .A1(n819), .A2(n604), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U678 ( .A(KEYINPUT77), .B(n607), .Z(G288) );
  NAND2_X1 U679 ( .A1(G61), .A2(n819), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(KEYINPUT78), .ZN(n615) );
  NAND2_X1 U681 ( .A1(G86), .A2(n815), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G48), .A2(n820), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n816), .A2(G73), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT2), .B(n611), .Z(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(G305) );
  NAND2_X1 U688 ( .A1(G85), .A2(n815), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G72), .A2(n816), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G60), .A2(n819), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G47), .A2(n820), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U695 ( .A(KEYINPUT66), .B(n622), .Z(G290) );
  NOR2_X1 U696 ( .A1(G164), .A2(G1384), .ZN(n723) );
  NOR2_X1 U697 ( .A1(n629), .A2(G2084), .ZN(n690) );
  INV_X1 U698 ( .A(n690), .ZN(n624) );
  INV_X1 U699 ( .A(n689), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n548), .A2(n625), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(KEYINPUT30), .ZN(n627) );
  NOR2_X1 U702 ( .A1(G168), .A2(n627), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT91), .ZN(n633) );
  XNOR2_X1 U704 ( .A(G2078), .B(KEYINPUT25), .ZN(n896) );
  NAND2_X1 U705 ( .A1(n669), .A2(n896), .ZN(n631) );
  XNOR2_X1 U706 ( .A(G1961), .B(KEYINPUT89), .ZN(n966) );
  NAND2_X1 U707 ( .A1(n629), .A2(n966), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n678) );
  OR2_X1 U709 ( .A1(n678), .A2(G171), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n635) );
  XNOR2_X1 U711 ( .A(KEYINPUT31), .B(KEYINPUT92), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n635), .B(n634), .ZN(n681) );
  NAND2_X1 U713 ( .A1(n669), .A2(G1996), .ZN(n636) );
  XNOR2_X1 U714 ( .A(n636), .B(KEYINPUT26), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n629), .A2(G1341), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n664) );
  NAND2_X1 U717 ( .A1(n819), .A2(G56), .ZN(n639) );
  XOR2_X1 U718 ( .A(KEYINPUT14), .B(n639), .Z(n647) );
  NAND2_X1 U719 ( .A1(G81), .A2(n815), .ZN(n640) );
  XOR2_X1 U720 ( .A(KEYINPUT12), .B(n640), .Z(n641) );
  XNOR2_X1 U721 ( .A(n641), .B(KEYINPUT69), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G68), .A2(n816), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n645) );
  NOR2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U725 ( .A(n648), .B(KEYINPUT70), .ZN(n650) );
  NAND2_X1 U726 ( .A1(G43), .A2(n820), .ZN(n649) );
  NAND2_X1 U727 ( .A1(G92), .A2(n815), .ZN(n652) );
  NAND2_X1 U728 ( .A1(G79), .A2(n816), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U730 ( .A1(G66), .A2(n819), .ZN(n654) );
  NAND2_X1 U731 ( .A1(G54), .A2(n820), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U734 ( .A(KEYINPUT15), .B(n657), .Z(n986) );
  INV_X1 U735 ( .A(n986), .ZN(n919) );
  NOR2_X1 U736 ( .A1(n664), .A2(n546), .ZN(n663) );
  INV_X1 U737 ( .A(G1348), .ZN(n782) );
  XNOR2_X1 U738 ( .A(n659), .B(n658), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n669), .A2(G2067), .ZN(n660) );
  AND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U741 ( .A1(n990), .A2(n664), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n667), .A2(n666), .ZN(n673) );
  INV_X1 U743 ( .A(G299), .ZN(n674) );
  NAND2_X1 U744 ( .A1(G2072), .A2(n669), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n668), .B(KEYINPUT27), .ZN(n671) );
  INV_X1 U746 ( .A(G1956), .ZN(n945) );
  NOR2_X1 U747 ( .A1(n669), .A2(n945), .ZN(n670) );
  NOR2_X1 U748 ( .A1(n671), .A2(n670), .ZN(n675) );
  NAND2_X1 U749 ( .A1(n674), .A2(n675), .ZN(n672) );
  NOR2_X1 U750 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n678), .A2(G171), .ZN(n679) );
  NAND2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n687) );
  NAND2_X1 U753 ( .A1(n687), .A2(G286), .ZN(n686) );
  NOR2_X1 U754 ( .A1(G2090), .A2(n629), .ZN(n747) );
  NOR2_X1 U755 ( .A1(G1971), .A2(n743), .ZN(n682) );
  XOR2_X1 U756 ( .A(KEYINPUT93), .B(n682), .Z(n683) );
  NOR2_X1 U757 ( .A1(n747), .A2(n683), .ZN(n684) );
  NAND2_X1 U758 ( .A1(n684), .A2(G303), .ZN(n685) );
  INV_X1 U759 ( .A(n687), .ZN(n688) );
  NOR2_X1 U760 ( .A1(n689), .A2(n688), .ZN(n692) );
  NAND2_X1 U761 ( .A1(G8), .A2(n690), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n696) );
  XNOR2_X1 U764 ( .A(n696), .B(n695), .ZN(n742) );
  NOR2_X1 U765 ( .A1(G1976), .A2(G288), .ZN(n927) );
  NOR2_X1 U766 ( .A1(G1971), .A2(G303), .ZN(n697) );
  NOR2_X1 U767 ( .A1(n927), .A2(n697), .ZN(n698) );
  NAND2_X1 U768 ( .A1(n742), .A2(n698), .ZN(n699) );
  XNOR2_X1 U769 ( .A(n699), .B(KEYINPUT96), .ZN(n702) );
  NAND2_X1 U770 ( .A1(G1976), .A2(G288), .ZN(n929) );
  XOR2_X1 U771 ( .A(G1981), .B(G305), .Z(n924) );
  INV_X1 U772 ( .A(n924), .ZN(n705) );
  NAND2_X1 U773 ( .A1(n927), .A2(KEYINPUT33), .ZN(n703) );
  NOR2_X1 U774 ( .A1(n743), .A2(n703), .ZN(n704) );
  OR2_X1 U775 ( .A1(n705), .A2(n704), .ZN(n737) );
  NAND2_X1 U776 ( .A1(G131), .A2(n1027), .ZN(n707) );
  NAND2_X1 U777 ( .A1(G95), .A2(n1028), .ZN(n706) );
  NAND2_X1 U778 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U779 ( .A1(G119), .A2(n1023), .ZN(n709) );
  NAND2_X1 U780 ( .A1(G107), .A2(n1024), .ZN(n708) );
  NAND2_X1 U781 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U782 ( .A1(n711), .A2(n710), .ZN(n1014) );
  INV_X1 U783 ( .A(G1991), .ZN(n894) );
  NOR2_X1 U784 ( .A1(n1014), .A2(n894), .ZN(n721) );
  XOR2_X1 U785 ( .A(KEYINPUT38), .B(KEYINPUT86), .Z(n713) );
  NAND2_X1 U786 ( .A1(G105), .A2(n1028), .ZN(n712) );
  XNOR2_X1 U787 ( .A(n713), .B(n712), .ZN(n717) );
  NAND2_X1 U788 ( .A1(G141), .A2(n1027), .ZN(n715) );
  NAND2_X1 U789 ( .A1(G117), .A2(n1024), .ZN(n714) );
  NAND2_X1 U790 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U791 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U792 ( .A1(n1023), .A2(G129), .ZN(n718) );
  NAND2_X1 U793 ( .A1(n719), .A2(n718), .ZN(n1016) );
  AND2_X1 U794 ( .A1(n1016), .A2(G1996), .ZN(n720) );
  NOR2_X1 U795 ( .A1(n721), .A2(n720), .ZN(n881) );
  NOR2_X1 U796 ( .A1(n723), .A2(n722), .ZN(n769) );
  XNOR2_X1 U797 ( .A(KEYINPUT87), .B(n769), .ZN(n724) );
  NOR2_X1 U798 ( .A1(n881), .A2(n724), .ZN(n762) );
  INV_X1 U799 ( .A(n762), .ZN(n736) );
  NAND2_X1 U800 ( .A1(G140), .A2(n1027), .ZN(n726) );
  NAND2_X1 U801 ( .A1(G104), .A2(n1028), .ZN(n725) );
  NAND2_X1 U802 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U803 ( .A(KEYINPUT34), .B(n727), .ZN(n732) );
  NAND2_X1 U804 ( .A1(G128), .A2(n1023), .ZN(n729) );
  NAND2_X1 U805 ( .A1(G116), .A2(n1024), .ZN(n728) );
  NAND2_X1 U806 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U807 ( .A(n730), .B(KEYINPUT35), .Z(n731) );
  NOR2_X1 U808 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U809 ( .A(KEYINPUT36), .B(n733), .Z(n734) );
  XNOR2_X1 U810 ( .A(KEYINPUT85), .B(n734), .ZN(n1037) );
  XNOR2_X1 U811 ( .A(G2067), .B(KEYINPUT37), .ZN(n767) );
  NOR2_X1 U812 ( .A1(n1037), .A2(n767), .ZN(n885) );
  NAND2_X1 U813 ( .A1(n769), .A2(n885), .ZN(n735) );
  NAND2_X1 U814 ( .A1(n736), .A2(n735), .ZN(n738) );
  INV_X1 U815 ( .A(n738), .ZN(n752) );
  NOR2_X1 U816 ( .A1(G1981), .A2(G305), .ZN(n739) );
  XOR2_X1 U817 ( .A(n739), .B(KEYINPUT24), .Z(n740) );
  NOR2_X1 U818 ( .A1(n743), .A2(n740), .ZN(n741) );
  XNOR2_X1 U819 ( .A(n741), .B(KEYINPUT88), .ZN(n746) );
  INV_X1 U820 ( .A(n743), .ZN(n744) );
  NOR2_X1 U821 ( .A1(n742), .A2(n744), .ZN(n745) );
  NOR2_X1 U822 ( .A1(n746), .A2(n745), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n747), .A2(G8), .ZN(n748) );
  OR2_X1 U824 ( .A1(G303), .A2(n748), .ZN(n749) );
  NAND2_X1 U825 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U826 ( .A1(n753), .A2(n547), .ZN(n755) );
  XNOR2_X1 U827 ( .A(n755), .B(n754), .ZN(n757) );
  XNOR2_X1 U828 ( .A(G1986), .B(G290), .ZN(n932) );
  NAND2_X1 U829 ( .A1(n932), .A2(n769), .ZN(n756) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n772) );
  NOR2_X1 U831 ( .A1(n1016), .A2(G1996), .ZN(n758) );
  XNOR2_X1 U832 ( .A(n758), .B(KEYINPUT98), .ZN(n876) );
  NOR2_X1 U833 ( .A1(G1986), .A2(G290), .ZN(n760) );
  NAND2_X1 U834 ( .A1(n894), .A2(n1014), .ZN(n880) );
  INV_X1 U835 ( .A(n880), .ZN(n759) );
  NOR2_X1 U836 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U837 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U838 ( .A1(n876), .A2(n763), .ZN(n764) );
  XOR2_X1 U839 ( .A(KEYINPUT39), .B(n764), .Z(n765) );
  NOR2_X1 U840 ( .A1(n885), .A2(n765), .ZN(n766) );
  XNOR2_X1 U841 ( .A(n766), .B(KEYINPUT99), .ZN(n768) );
  NAND2_X1 U842 ( .A1(n1037), .A2(n767), .ZN(n873) );
  NAND2_X1 U843 ( .A1(n768), .A2(n873), .ZN(n770) );
  NAND2_X1 U844 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U846 ( .A(n773), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U847 ( .A(G2435), .B(KEYINPUT102), .Z(n775) );
  XNOR2_X1 U848 ( .A(KEYINPUT101), .B(G2438), .ZN(n774) );
  XNOR2_X1 U849 ( .A(n775), .B(n774), .ZN(n779) );
  XOR2_X1 U850 ( .A(G2451), .B(G2443), .Z(n777) );
  XNOR2_X1 U851 ( .A(G1341), .B(KEYINPUT100), .ZN(n776) );
  XNOR2_X1 U852 ( .A(n777), .B(n776), .ZN(n778) );
  XOR2_X1 U853 ( .A(n779), .B(n778), .Z(n781) );
  XNOR2_X1 U854 ( .A(G2427), .B(G2446), .ZN(n780) );
  XNOR2_X1 U855 ( .A(n781), .B(n780), .ZN(n785) );
  XNOR2_X1 U856 ( .A(G2430), .B(G2454), .ZN(n783) );
  XNOR2_X1 U857 ( .A(n783), .B(n782), .ZN(n784) );
  XOR2_X1 U858 ( .A(n785), .B(n784), .Z(n786) );
  AND2_X1 U859 ( .A1(G14), .A2(n786), .ZN(G401) );
  AND2_X1 U860 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U861 ( .A(G132), .ZN(G219) );
  INV_X1 U862 ( .A(G82), .ZN(G220) );
  INV_X1 U863 ( .A(G57), .ZN(G237) );
  NAND2_X1 U864 ( .A1(G7), .A2(G661), .ZN(n787) );
  XNOR2_X1 U865 ( .A(n787), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U866 ( .A(G223), .ZN(n847) );
  NAND2_X1 U867 ( .A1(n847), .A2(G567), .ZN(n788) );
  XOR2_X1 U868 ( .A(KEYINPUT11), .B(n788), .Z(G234) );
  INV_X1 U869 ( .A(G860), .ZN(n980) );
  OR2_X1 U870 ( .A1(n990), .A2(n980), .ZN(G153) );
  NAND2_X1 U871 ( .A1(G868), .A2(G301), .ZN(n790) );
  INV_X1 U872 ( .A(G868), .ZN(n830) );
  NAND2_X1 U873 ( .A1(n919), .A2(n830), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(G284) );
  NOR2_X1 U875 ( .A1(G286), .A2(n830), .ZN(n792) );
  NOR2_X1 U876 ( .A1(G868), .A2(G299), .ZN(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(G297) );
  NAND2_X1 U878 ( .A1(n980), .A2(G559), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n793), .A2(n986), .ZN(n794) );
  XNOR2_X1 U880 ( .A(n794), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U881 ( .A1(G868), .A2(n990), .ZN(n797) );
  NAND2_X1 U882 ( .A1(G868), .A2(n986), .ZN(n795) );
  NOR2_X1 U883 ( .A1(G559), .A2(n795), .ZN(n796) );
  NOR2_X1 U884 ( .A1(n797), .A2(n796), .ZN(G282) );
  NAND2_X1 U885 ( .A1(n1023), .A2(G123), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n798), .B(KEYINPUT18), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G135), .A2(n1027), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U889 ( .A(KEYINPUT72), .B(n801), .ZN(n804) );
  NAND2_X1 U890 ( .A1(G99), .A2(n1028), .ZN(n802) );
  XNOR2_X1 U891 ( .A(KEYINPUT73), .B(n802), .ZN(n803) );
  NOR2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n1024), .A2(G111), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n1034) );
  XOR2_X1 U895 ( .A(G2096), .B(KEYINPUT74), .Z(n807) );
  XNOR2_X1 U896 ( .A(n1034), .B(n807), .ZN(n809) );
  INV_X1 U897 ( .A(G2100), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(G156) );
  XOR2_X1 U899 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n811) );
  XNOR2_X1 U900 ( .A(G166), .B(KEYINPUT19), .ZN(n810) );
  XNOR2_X1 U901 ( .A(n811), .B(n810), .ZN(n814) );
  XNOR2_X1 U902 ( .A(G290), .B(G305), .ZN(n812) );
  XNOR2_X1 U903 ( .A(n812), .B(G299), .ZN(n813) );
  XNOR2_X1 U904 ( .A(n814), .B(n813), .ZN(n827) );
  NAND2_X1 U905 ( .A1(G93), .A2(n815), .ZN(n818) );
  NAND2_X1 U906 ( .A1(G80), .A2(n816), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n818), .A2(n817), .ZN(n824) );
  NAND2_X1 U908 ( .A1(G67), .A2(n819), .ZN(n822) );
  NAND2_X1 U909 ( .A1(G55), .A2(n820), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U911 ( .A1(n824), .A2(n823), .ZN(n825) );
  XOR2_X1 U912 ( .A(KEYINPUT76), .B(n825), .Z(n979) );
  XNOR2_X1 U913 ( .A(G288), .B(n979), .ZN(n826) );
  XNOR2_X1 U914 ( .A(n827), .B(n826), .ZN(n989) );
  NAND2_X1 U915 ( .A1(G559), .A2(n986), .ZN(n828) );
  XOR2_X1 U916 ( .A(n990), .B(n828), .Z(n981) );
  XOR2_X1 U917 ( .A(n989), .B(n981), .Z(n829) );
  NOR2_X1 U918 ( .A1(n830), .A2(n829), .ZN(n832) );
  NOR2_X1 U919 ( .A1(n979), .A2(G868), .ZN(n831) );
  NOR2_X1 U920 ( .A1(n832), .A2(n831), .ZN(G295) );
  NAND2_X1 U921 ( .A1(G2078), .A2(G2084), .ZN(n833) );
  XOR2_X1 U922 ( .A(KEYINPUT20), .B(n833), .Z(n834) );
  NAND2_X1 U923 ( .A1(G2090), .A2(n834), .ZN(n835) );
  XNOR2_X1 U924 ( .A(KEYINPUT21), .B(n835), .ZN(n836) );
  NAND2_X1 U925 ( .A1(n836), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U926 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U927 ( .A1(G120), .A2(G69), .ZN(n837) );
  NOR2_X1 U928 ( .A1(G237), .A2(n837), .ZN(n838) );
  NAND2_X1 U929 ( .A1(G108), .A2(n838), .ZN(n984) );
  NAND2_X1 U930 ( .A1(n984), .A2(G567), .ZN(n844) );
  NOR2_X1 U931 ( .A1(G220), .A2(G219), .ZN(n839) );
  XNOR2_X1 U932 ( .A(KEYINPUT22), .B(n839), .ZN(n840) );
  NAND2_X1 U933 ( .A1(n840), .A2(G96), .ZN(n841) );
  NOR2_X1 U934 ( .A1(G218), .A2(n841), .ZN(n842) );
  XOR2_X1 U935 ( .A(KEYINPUT82), .B(n842), .Z(n985) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n985), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n844), .A2(n843), .ZN(n1049) );
  NAND2_X1 U938 ( .A1(G661), .A2(G483), .ZN(n845) );
  XOR2_X1 U939 ( .A(KEYINPUT83), .B(n845), .Z(n846) );
  NOR2_X1 U940 ( .A1(n1049), .A2(n846), .ZN(n849) );
  NAND2_X1 U941 ( .A1(n849), .A2(G36), .ZN(G176) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n847), .ZN(G217) );
  AND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n848) );
  NAND2_X1 U944 ( .A1(G661), .A2(n848), .ZN(G259) );
  NAND2_X1 U945 ( .A1(G3), .A2(G1), .ZN(n850) );
  NAND2_X1 U946 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT103), .B(n851), .Z(G188) );
  XOR2_X1 U948 ( .A(G69), .B(KEYINPUT104), .Z(G235) );
  NAND2_X1 U950 ( .A1(G100), .A2(n1028), .ZN(n853) );
  NAND2_X1 U951 ( .A1(G112), .A2(n1024), .ZN(n852) );
  NAND2_X1 U952 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U953 ( .A(KEYINPUT106), .B(n854), .ZN(n859) );
  NAND2_X1 U954 ( .A1(n1023), .A2(G124), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G136), .A2(n1027), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U958 ( .A1(n859), .A2(n858), .ZN(G162) );
  INV_X1 U959 ( .A(KEYINPUT55), .ZN(n915) );
  XOR2_X1 U960 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n872) );
  NAND2_X1 U961 ( .A1(G139), .A2(n1027), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G103), .A2(n1028), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n867) );
  NAND2_X1 U964 ( .A1(n1024), .A2(G115), .ZN(n862) );
  XOR2_X1 U965 ( .A(KEYINPUT107), .B(n862), .Z(n864) );
  NAND2_X1 U966 ( .A1(n1023), .A2(G127), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U968 ( .A(KEYINPUT47), .B(n865), .Z(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n1019) );
  XOR2_X1 U970 ( .A(G2072), .B(n1019), .Z(n869) );
  XOR2_X1 U971 ( .A(G164), .B(G2078), .Z(n868) );
  NOR2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n870), .B(KEYINPUT114), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n879) );
  XOR2_X1 U976 ( .A(G2090), .B(G162), .Z(n875) );
  NOR2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n877), .B(KEYINPUT51), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n888) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n883) );
  XOR2_X1 U981 ( .A(G160), .B(G2084), .Z(n882) );
  NOR2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n884), .A2(n1034), .ZN(n886) );
  NOR2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n887) );
  NAND2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U986 ( .A(KEYINPUT116), .B(n889), .ZN(n890) );
  XOR2_X1 U987 ( .A(KEYINPUT52), .B(n890), .Z(n891) );
  NAND2_X1 U988 ( .A1(n915), .A2(n891), .ZN(n892) );
  NAND2_X1 U989 ( .A1(n892), .A2(G29), .ZN(n977) );
  XOR2_X1 U990 ( .A(G2090), .B(G35), .Z(n893) );
  XNOR2_X1 U991 ( .A(KEYINPUT117), .B(n893), .ZN(n909) );
  XOR2_X1 U992 ( .A(G32), .B(G1996), .Z(n901) );
  XNOR2_X1 U993 ( .A(G25), .B(n894), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n895), .A2(G28), .ZN(n899) );
  XNOR2_X1 U995 ( .A(G27), .B(n896), .ZN(n897) );
  XNOR2_X1 U996 ( .A(KEYINPUT119), .B(n897), .ZN(n898) );
  NOR2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n900) );
  NAND2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n906) );
  XNOR2_X1 U999 ( .A(G2067), .B(G26), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(G2072), .B(G33), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1002 ( .A(KEYINPUT118), .B(n904), .Z(n905) );
  NOR2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n907), .B(KEYINPUT53), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n910), .B(KEYINPUT120), .ZN(n913) );
  XOR2_X1 U1007 ( .A(G2084), .B(G34), .Z(n911) );
  XNOR2_X1 U1008 ( .A(KEYINPUT54), .B(n911), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n917) );
  INV_X1 U1011 ( .A(G29), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1013 ( .A1(G11), .A2(n918), .ZN(n975) );
  XNOR2_X1 U1014 ( .A(G16), .B(KEYINPUT56), .ZN(n944) );
  XNOR2_X1 U1015 ( .A(G301), .B(G1961), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(n919), .B(G1348), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT122), .B(n922), .ZN(n942) );
  XOR2_X1 U1019 ( .A(G1966), .B(G168), .Z(n923) );
  XNOR2_X1 U1020 ( .A(KEYINPUT121), .B(n923), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(n926), .B(KEYINPUT57), .ZN(n938) );
  XNOR2_X1 U1023 ( .A(G166), .B(G1971), .ZN(n934) );
  INV_X1 U1024 ( .A(n927), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1026 ( .A(KEYINPUT123), .B(n930), .Z(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(G1956), .B(G299), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n940) );
  XNOR2_X1 U1032 ( .A(G1341), .B(n990), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n973) );
  INV_X1 U1036 ( .A(G16), .ZN(n971) );
  XNOR2_X1 U1037 ( .A(G20), .B(n945), .ZN(n949) );
  XNOR2_X1 U1038 ( .A(G1981), .B(G6), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(G1341), .B(G19), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n952) );
  XOR2_X1 U1042 ( .A(KEYINPUT59), .B(G1348), .Z(n950) );
  XNOR2_X1 U1043 ( .A(G4), .B(n950), .ZN(n951) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(n953), .B(KEYINPUT60), .ZN(n956) );
  XOR2_X1 U1046 ( .A(G1966), .B(G21), .Z(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT124), .B(n954), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(n957), .B(KEYINPUT125), .ZN(n965) );
  XOR2_X1 U1050 ( .A(G1976), .B(KEYINPUT126), .Z(n958) );
  XNOR2_X1 U1051 ( .A(G23), .B(n958), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G1986), .B(G24), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1056 ( .A(KEYINPUT58), .B(n963), .Z(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n968) );
  XOR2_X1 U1058 ( .A(G5), .B(n966), .Z(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(KEYINPUT61), .B(n969), .ZN(n970) );
  NAND2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1062 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1063 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1064 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1065 ( .A(KEYINPUT62), .B(n978), .Z(G311) );
  XNOR2_X1 U1066 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  XOR2_X1 U1067 ( .A(n979), .B(KEYINPUT75), .Z(n983) );
  NAND2_X1 U1068 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1069 ( .A(n983), .B(n982), .ZN(G145) );
  INV_X1 U1070 ( .A(G120), .ZN(G236) );
  INV_X1 U1071 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(G325) );
  INV_X1 U1073 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1074 ( .A(KEYINPUT111), .B(G286), .Z(n988) );
  XNOR2_X1 U1075 ( .A(G171), .B(n986), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(n988), .B(n987), .ZN(n992) );
  XOR2_X1 U1077 ( .A(n990), .B(n989), .Z(n991) );
  XNOR2_X1 U1078 ( .A(n992), .B(n991), .ZN(n993) );
  NOR2_X1 U1079 ( .A1(G37), .A2(n993), .ZN(G397) );
  XOR2_X1 U1080 ( .A(KEYINPUT43), .B(G2100), .Z(n995) );
  XNOR2_X1 U1081 ( .A(G2067), .B(G2084), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(n995), .B(n994), .ZN(n996) );
  XOR2_X1 U1083 ( .A(n996), .B(KEYINPUT42), .Z(n998) );
  XNOR2_X1 U1084 ( .A(G2090), .B(KEYINPUT105), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(n998), .B(n997), .ZN(n1002) );
  XOR2_X1 U1086 ( .A(G2096), .B(G2678), .Z(n1000) );
  XNOR2_X1 U1087 ( .A(G2078), .B(G2072), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(n1000), .B(n999), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(n1002), .B(n1001), .Z(G227) );
  XOR2_X1 U1090 ( .A(G1976), .B(G1971), .Z(n1004) );
  XNOR2_X1 U1091 ( .A(G1996), .B(G1981), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1004), .B(n1003), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(n1005), .B(G2474), .Z(n1007) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G1956), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1007), .B(n1006), .ZN(n1011) );
  XOR2_X1 U1096 ( .A(KEYINPUT41), .B(G1961), .Z(n1009) );
  XNOR2_X1 U1097 ( .A(G1991), .B(G1986), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(n1009), .B(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(n1011), .B(n1010), .ZN(G229) );
  XOR2_X1 U1100 ( .A(KEYINPUT46), .B(KEYINPUT108), .Z(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT109), .B(KEYINPUT48), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(n1013), .B(n1012), .ZN(n1015) );
  XOR2_X1 U1103 ( .A(n1015), .B(n1014), .Z(n1018) );
  XOR2_X1 U1104 ( .A(G164), .B(n1016), .Z(n1017) );
  XNOR2_X1 U1105 ( .A(n1018), .B(n1017), .ZN(n1020) );
  XOR2_X1 U1106 ( .A(n1020), .B(n1019), .Z(n1022) );
  XNOR2_X1 U1107 ( .A(G160), .B(G162), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1022), .B(n1021), .ZN(n1039) );
  NAND2_X1 U1109 ( .A1(G130), .A2(n1023), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(G118), .A2(n1024), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1033) );
  NAND2_X1 U1112 ( .A1(G142), .A2(n1027), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(G106), .A2(n1028), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(n1031), .B(KEYINPUT45), .Z(n1032) );
  NOR2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1035) );
  XNOR2_X1 U1117 ( .A(n1035), .B(n1034), .ZN(n1036) );
  XOR2_X1 U1118 ( .A(n1037), .B(n1036), .Z(n1038) );
  XNOR2_X1 U1119 ( .A(n1039), .B(n1038), .ZN(n1040) );
  NOR2_X1 U1120 ( .A1(G37), .A2(n1040), .ZN(n1041) );
  XNOR2_X1 U1121 ( .A(KEYINPUT110), .B(n1041), .ZN(G395) );
  NOR2_X1 U1122 ( .A1(G401), .A2(n1049), .ZN(n1046) );
  NOR2_X1 U1123 ( .A1(G227), .A2(G229), .ZN(n1043) );
  XNOR2_X1 U1124 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n1042) );
  XNOR2_X1 U1125 ( .A(n1043), .B(n1042), .ZN(n1044) );
  NOR2_X1 U1126 ( .A1(G397), .A2(n1044), .ZN(n1045) );
  NAND2_X1 U1127 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NOR2_X1 U1128 ( .A1(n1047), .A2(G395), .ZN(n1048) );
  XNOR2_X1 U1129 ( .A(n1048), .B(KEYINPUT113), .ZN(G225) );
  INV_X1 U1130 ( .A(G225), .ZN(G308) );
  INV_X1 U1131 ( .A(n1049), .ZN(G319) );
  INV_X1 U1132 ( .A(G108), .ZN(G238) );
endmodule

