//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G77), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n219), .A2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G58), .A2(G232), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n202), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n239), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  OAI211_X1 g0048(.A(G1), .B(G13), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G222), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT66), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  AND3_X1   g0057(.A1(new_n255), .A2(new_n257), .A3(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n257), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n258), .A2(G223), .B1(new_n219), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n249), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n248), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT65), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT65), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G41), .A2(G45), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n249), .A2(G274), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n263), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G226), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n261), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n215), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n206), .A2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n281), .A2(G50), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n207), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G150), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n207), .A2(new_n247), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n288), .A2(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G58), .A2(G68), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n207), .B1(new_n293), .B2(new_n240), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n279), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n261), .A2(new_n274), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n277), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(KEYINPUT67), .A2(KEYINPUT9), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT67), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n296), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n287), .A2(new_n303), .A3(new_n304), .A4(new_n295), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n275), .A2(G200), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  NOR4_X1   g0109(.A1(new_n261), .A2(KEYINPUT68), .A3(new_n309), .A4(new_n274), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT68), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n297), .B2(G190), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT10), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n308), .B(new_n315), .C1(new_n310), .C2(new_n312), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n301), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n272), .A2(G244), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n258), .A2(G238), .B1(G107), .B2(new_n259), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n270), .B(new_n318), .C1(new_n321), .C2(new_n249), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G200), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n283), .A2(G77), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n282), .A2(new_n324), .B1(new_n219), .B2(new_n281), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT15), .B(G87), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n289), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(G20), .B2(new_n219), .ZN(new_n328));
  INV_X1    g0128(.A(new_n288), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G20), .A2(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n325), .B1(new_n332), .B2(new_n279), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n323), .B(new_n333), .C1(new_n309), .C2(new_n322), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n322), .A2(G179), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n333), .B1(new_n322), .B2(new_n276), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n317), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT7), .B1(new_n259), .B2(new_n207), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT7), .ZN(new_n340));
  AOI211_X1 g0140(.A(new_n340), .B(G20), .C1(new_n255), .C2(new_n257), .ZN(new_n341));
  OAI21_X1  g0141(.A(G68), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G58), .A2(G68), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G20), .B1(new_n344), .B2(new_n293), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n330), .A2(G159), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n280), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n340), .B1(new_n250), .B2(G20), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n207), .B1(new_n203), .B2(new_n343), .ZN(new_n354));
  INV_X1    g0154(.A(G159), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n291), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT73), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT73), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n345), .A2(new_n358), .A3(new_n346), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n353), .A2(G68), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n350), .B1(new_n360), .B2(KEYINPUT16), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n359), .ZN(new_n362));
  AND4_X1   g0162(.A1(new_n350), .A2(new_n342), .A3(KEYINPUT16), .A4(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n349), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n255), .A2(new_n257), .A3(G226), .A4(G1698), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT75), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n250), .A2(KEYINPUT75), .A3(G226), .A4(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n255), .A2(new_n257), .A3(G223), .A4(new_n251), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n249), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n272), .A2(G232), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n270), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(G200), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n268), .A2(new_n269), .B1(new_n272), .B2(G232), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n372), .B1(new_n367), .B2(new_n368), .ZN(new_n379));
  OAI211_X1 g0179(.A(G190), .B(new_n378), .C1(new_n379), .C2(new_n249), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n329), .A2(new_n283), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n382), .A2(new_n282), .B1(new_n281), .B2(new_n329), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n364), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT77), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n342), .A2(new_n362), .A3(KEYINPUT16), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT74), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n360), .A2(new_n350), .A3(KEYINPUT16), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n383), .B1(new_n392), .B2(new_n349), .ZN(new_n393));
  NAND2_X1  g0193(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n386), .A2(new_n387), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n381), .A4(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(G169), .B1(new_n374), .B2(new_n376), .ZN(new_n398));
  OAI211_X1 g0198(.A(G179), .B(new_n378), .C1(new_n379), .C2(new_n249), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT18), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT76), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n202), .B1(new_n351), .B2(new_n352), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n345), .A2(new_n346), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n348), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n279), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n391), .B2(new_n390), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n404), .B(new_n400), .C1(new_n409), .C2(new_n383), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n402), .A2(new_n403), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n403), .B1(new_n402), .B2(new_n410), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n397), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n330), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n415));
  INV_X1    g0215(.A(G77), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(new_n289), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT11), .B1(new_n417), .B2(new_n279), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n280), .A2(G68), .A3(new_n281), .A4(new_n283), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT12), .ZN(new_n421));
  INV_X1    g0221(.A(new_n281), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(new_n202), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n281), .A2(KEYINPUT12), .A3(G68), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n420), .B(KEYINPUT71), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n417), .A2(KEYINPUT11), .A3(new_n279), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n419), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT71), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n414), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n426), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n418), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n429), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n433), .A2(KEYINPUT72), .A3(new_n434), .A4(new_n425), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n250), .A2(G232), .A3(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G97), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n255), .A2(new_n257), .A3(G226), .A4(new_n251), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n271), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n268), .A2(new_n269), .B1(new_n272), .B2(G238), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(KEYINPUT70), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT70), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n443), .A2(new_n449), .A3(new_n445), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(G169), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n451), .A2(KEYINPUT14), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT14), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n448), .A2(new_n453), .A3(G169), .A4(new_n450), .ZN(new_n454));
  INV_X1    g0254(.A(new_n447), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT13), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n441), .B2(new_n442), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G179), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n436), .B1(new_n452), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n458), .A2(G190), .B1(new_n431), .B2(new_n435), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n448), .A2(G200), .A3(new_n450), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n338), .A2(new_n413), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G107), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n351), .B2(new_n352), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n469), .A2(KEYINPUT78), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n353), .A2(KEYINPUT78), .A3(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(KEYINPUT6), .A3(G97), .ZN(new_n472));
  INV_X1    g0272(.A(G97), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n472), .B1(new_n476), .B2(KEYINPUT6), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n477), .A2(G20), .B1(G77), .B2(new_n330), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n470), .A2(new_n471), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n206), .A2(G33), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n280), .A2(new_n281), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G97), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(G97), .B2(new_n422), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n482), .B(KEYINPUT79), .C1(G97), .C2(new_n422), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n479), .A2(new_n279), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT82), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(KEYINPUT5), .B2(new_n248), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT5), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n492), .A2(KEYINPUT80), .A3(G41), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT80), .B1(new_n492), .B2(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n490), .A2(new_n248), .A3(KEYINPUT5), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT81), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n262), .A2(G1), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n492), .A2(G41), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n249), .A2(G274), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n488), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n501), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(KEYINPUT82), .A3(new_n494), .A4(new_n497), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n255), .A2(new_n257), .A3(G244), .A4(new_n251), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n250), .A2(G250), .A3(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n508), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n495), .A2(new_n496), .A3(new_n499), .A4(new_n500), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n513), .A2(new_n249), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n512), .A2(new_n271), .B1(new_n514), .B2(G257), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n505), .A2(new_n515), .A3(KEYINPUT83), .A4(G190), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT83), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n505), .A2(new_n515), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(G200), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n309), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n487), .B(new_n516), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n471), .A2(new_n478), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n469), .A2(KEYINPUT78), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n279), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n485), .A2(new_n486), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n505), .A2(new_n515), .A3(new_n298), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n518), .A2(new_n276), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n249), .A2(G274), .A3(new_n499), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n206), .A2(G45), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n247), .A2(new_n248), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(G250), .C1(new_n532), .C2(new_n215), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT84), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n255), .A2(new_n257), .A3(G244), .A4(G1698), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n255), .A2(new_n257), .A3(G238), .A4(new_n251), .ZN(new_n537));
  INV_X1    g0337(.A(G116), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n247), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n271), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT84), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n530), .A2(new_n533), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n535), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G169), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n298), .B2(new_n545), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n207), .B1(new_n438), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G87), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n475), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n255), .A2(new_n257), .A3(new_n207), .A4(G68), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n548), .B1(new_n289), .B2(new_n473), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n279), .B1(new_n422), .B2(new_n326), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n481), .B2(new_n326), .ZN(new_n557));
  INV_X1    g0357(.A(new_n481), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G87), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n545), .B2(G200), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n530), .A2(new_n533), .A3(new_n543), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n543), .B1(new_n530), .B2(new_n533), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(G190), .A3(new_n542), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n547), .A2(new_n557), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n521), .A2(new_n529), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT87), .ZN(new_n568));
  XNOR2_X1  g0368(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n250), .A2(new_n569), .A3(new_n207), .A4(G87), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n255), .A2(new_n257), .A3(new_n207), .A4(G87), .ZN(new_n571));
  XOR2_X1   g0371(.A(KEYINPUT86), .B(KEYINPUT22), .Z(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT23), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n207), .B2(G107), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n468), .A2(KEYINPUT23), .A3(G20), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n539), .A2(new_n207), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n568), .B1(new_n574), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n580), .B1(new_n570), .B2(new_n573), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n568), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT24), .B1(new_n585), .B2(new_n568), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n584), .B(new_n279), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n422), .A2(new_n468), .ZN(new_n590));
  NOR2_X1   g0390(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n590), .B2(new_n591), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n592), .A2(new_n594), .B1(new_n558), .B2(G107), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n258), .A2(G257), .B1(G33), .B2(G294), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n255), .A2(new_n257), .A3(G250), .A4(new_n251), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT89), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n271), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n514), .A2(G264), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n505), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n298), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n502), .A2(new_n504), .B1(G264), .B2(new_n514), .ZN(new_n607));
  AOI21_X1  g0407(.A(G169), .B1(new_n607), .B2(new_n603), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n596), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n595), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n574), .A2(new_n581), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT87), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(KEYINPUT24), .A3(new_n586), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n280), .B1(new_n582), .B2(new_n583), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n505), .A2(new_n603), .A3(new_n604), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(G190), .ZN(new_n618));
  AOI21_X1  g0418(.A(G200), .B1(new_n607), .B2(new_n603), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n510), .B(new_n207), .C1(G33), .C2(new_n473), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n622), .B(new_n279), .C1(new_n207), .C2(G116), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT20), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n281), .A2(G116), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n558), .B2(G116), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n255), .A2(new_n257), .A3(G257), .A4(new_n251), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n250), .A2(KEYINPUT85), .A3(G257), .A4(new_n251), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n258), .A2(G264), .B1(G303), .B2(new_n259), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n271), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n514), .A2(G270), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n505), .A2(new_n637), .A3(G190), .A4(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n505), .A2(new_n637), .A3(new_n638), .ZN(new_n640));
  INV_X1    g0440(.A(G200), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n629), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(G179), .A3(new_n628), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT21), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n505), .A2(new_n637), .A3(new_n638), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n276), .B1(new_n625), .B2(new_n627), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n645), .A2(new_n644), .A3(new_n646), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n642), .B(new_n643), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n567), .A2(new_n621), .A3(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n467), .A2(new_n650), .ZN(G372));
  NAND2_X1  g0451(.A1(new_n364), .A2(new_n384), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n404), .B1(new_n652), .B2(new_n400), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n393), .A2(KEYINPUT18), .A3(new_n401), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n337), .B1(new_n463), .B2(new_n462), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n451), .A2(KEYINPUT14), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n459), .A3(new_n454), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n436), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n388), .A2(new_n396), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n661), .A2(new_n662), .B1(new_n314), .B2(new_n316), .ZN(new_n663));
  OAI211_X1 g0463(.A(KEYINPUT90), .B(new_n655), .C1(new_n659), .C2(new_n660), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n301), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n276), .B1(new_n564), .B2(new_n542), .ZN(new_n667));
  AND4_X1   g0467(.A1(G179), .A2(new_n535), .A3(new_n542), .A4(new_n544), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n557), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n560), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n535), .A2(new_n542), .A3(new_n544), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n565), .B(new_n670), .C1(new_n641), .C2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n666), .B1(new_n529), .B2(new_n673), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n524), .A2(new_n525), .B1(new_n518), .B2(new_n276), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n566), .A2(KEYINPUT26), .A3(new_n675), .A4(new_n527), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n643), .B1(new_n648), .B2(new_n647), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n298), .A2(new_n505), .A3(new_n603), .A4(new_n604), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n616), .A2(new_n679), .A3(new_n608), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n620), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n677), .B(new_n669), .C1(new_n681), .C2(new_n567), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n467), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n665), .A2(new_n683), .ZN(G369));
  INV_X1    g0484(.A(new_n649), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n688), .A3(G213), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n628), .A2(new_n691), .ZN(new_n692));
  MUX2_X1   g0492(.A(new_n678), .B(new_n685), .S(new_n692), .Z(new_n693));
  XNOR2_X1  g0493(.A(KEYINPUT91), .B(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n610), .A2(new_n620), .ZN(new_n697));
  INV_X1    g0497(.A(new_n691), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT92), .B1(new_n616), .B2(new_n698), .ZN(new_n699));
  OR3_X1    g0499(.A1(new_n616), .A2(KEYINPUT92), .A3(new_n698), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n610), .B2(new_n698), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT93), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n678), .A2(new_n698), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n701), .A2(new_n705), .B1(new_n610), .B2(new_n691), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n704), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n210), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n551), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n213), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n671), .A2(G179), .A3(new_n515), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n605), .A3(new_n640), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n716), .A2(new_n605), .A3(new_n640), .A4(KEYINPUT30), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n671), .A2(G179), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n617), .A3(new_n645), .A4(new_n518), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n691), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n650), .A2(new_n698), .B1(new_n715), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n698), .A2(new_n715), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n719), .A2(new_n722), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT94), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n720), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n727), .A2(KEYINPUT94), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n694), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n682), .A2(new_n698), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT29), .B1(new_n733), .B2(KEYINPUT95), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT95), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n735), .B(new_n736), .C1(new_n682), .C2(new_n698), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n732), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT96), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n714), .B1(new_n739), .B2(G1), .ZN(G364));
  AND2_X1   g0540(.A1(new_n207), .A2(G13), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n206), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n709), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n693), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n215), .B1(G20), .B2(new_n276), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT97), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT98), .Z(new_n755));
  NOR2_X1   g0555(.A1(new_n708), .A2(new_n250), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n214), .A2(new_n262), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n756), .B(new_n757), .C1(new_n262), .C2(new_n245), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n708), .A2(new_n259), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n759), .A2(G355), .B1(new_n538), .B2(new_n708), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n755), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(G20), .A2(G179), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT99), .Z(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n309), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n641), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(G200), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G68), .A2(new_n765), .B1(new_n766), .B2(new_n219), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n763), .A2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n767), .B1(new_n201), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G179), .A2(G200), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(G20), .A3(new_n309), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G159), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT32), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(G190), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n207), .A2(new_n309), .A3(new_n641), .A4(G179), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n250), .B1(new_n779), .B2(new_n473), .C1(new_n781), .C2(new_n550), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n768), .A2(new_n641), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR4_X1   g0584(.A1(new_n207), .A2(new_n641), .A3(G179), .A4(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n784), .A2(new_n240), .B1(new_n789), .B2(new_n468), .ZN(new_n790));
  NOR4_X1   g0590(.A1(new_n771), .A2(new_n776), .A3(new_n782), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT101), .ZN(new_n793));
  INV_X1    g0593(.A(new_n789), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G283), .B1(G326), .B2(new_n783), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n250), .B1(new_n774), .B2(G329), .ZN(new_n796));
  INV_X1    g0596(.A(G294), .ZN(new_n797));
  INV_X1    g0597(.A(G303), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(new_n779), .B2(new_n797), .C1(new_n798), .C2(new_n781), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT33), .B(G317), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(new_n765), .B2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G311), .A2(new_n766), .B1(new_n769), .B2(G322), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n795), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n792), .A2(KEYINPUT101), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n793), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n761), .B1(new_n805), .B2(new_n751), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n745), .B1(new_n750), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n696), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n693), .A2(new_n695), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n807), .B1(new_n745), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT102), .ZN(G396));
  OAI21_X1  g0612(.A(new_n334), .B1(new_n333), .B2(new_n698), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n337), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n337), .A2(new_n691), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n733), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n725), .A2(new_n731), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n695), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n819), .A2(new_n821), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n822), .A2(new_n745), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT104), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n818), .A2(new_n747), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT103), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n250), .B1(new_n780), .B2(G107), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n765), .A2(G283), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G311), .A2(new_n774), .B1(new_n778), .B2(G97), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n829), .B(new_n830), .C1(new_n798), .C2(new_n784), .ZN(new_n831));
  INV_X1    g0631(.A(new_n766), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n832), .A2(new_n538), .B1(new_n827), .B2(new_n828), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n789), .A2(new_n550), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n770), .A2(new_n797), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n831), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G143), .A2(new_n769), .B1(new_n766), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  INV_X1    g0638(.A(new_n765), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n838), .B2(new_n784), .C1(new_n290), .C2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT34), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n250), .B1(new_n842), .B2(new_n773), .C1(new_n781), .C2(new_n240), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n789), .A2(new_n202), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n843), .B(new_n844), .C1(G58), .C2(new_n778), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n836), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n752), .A2(new_n747), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n846), .A2(new_n752), .B1(G77), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n744), .B1(new_n826), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n824), .A2(new_n825), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n825), .B1(new_n824), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(G384));
  OR2_X1    g0652(.A1(new_n477), .A2(KEYINPUT35), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n477), .A2(KEYINPUT35), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n853), .A2(G116), .A3(new_n216), .A4(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT36), .Z(new_n856));
  NAND3_X1  g0656(.A1(new_n214), .A2(new_n219), .A3(new_n343), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n206), .B(G13), .C1(new_n857), .C2(new_n241), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n279), .B1(new_n360), .B2(KEYINPUT16), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n391), .B2(new_n390), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n400), .B1(new_n861), .B2(new_n383), .ZN(new_n862));
  INV_X1    g0662(.A(new_n689), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n861), .B2(new_n383), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n864), .A3(new_n385), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n400), .B1(new_n409), .B2(new_n383), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT37), .B1(new_n867), .B2(KEYINPUT105), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT105), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n870), .B(new_n400), .C1(new_n409), .C2(new_n383), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n689), .B(KEYINPUT106), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n409), .B2(new_n383), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n385), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n866), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT76), .B1(new_n653), .B2(new_n654), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n402), .A2(new_n403), .A3(new_n410), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n660), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n875), .B1(new_n878), .B2(new_n864), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT38), .B(new_n875), .C1(new_n878), .C2(new_n864), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n867), .A2(new_n873), .A3(new_n385), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n869), .B2(new_n874), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n388), .A2(new_n396), .A3(new_n402), .A4(new_n410), .ZN(new_n887));
  INV_X1    g0687(.A(new_n873), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n880), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n882), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n461), .A2(new_n691), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n883), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n655), .A2(new_n872), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n881), .A2(new_n882), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n436), .A2(new_n691), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n461), .A2(new_n465), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n436), .B(new_n691), .C1(new_n658), .C2(new_n464), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n682), .A2(new_n818), .A3(new_n698), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n904), .B2(new_n816), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n897), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n896), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n467), .B1(new_n734), .B2(new_n737), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n665), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n907), .B(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n817), .B1(new_n900), .B2(new_n901), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n521), .A2(new_n529), .A3(new_n566), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n912), .A2(new_n685), .A3(new_n697), .A4(new_n698), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n724), .A2(new_n715), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n723), .A2(new_n726), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT40), .B1(new_n881), .B2(new_n882), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n892), .A2(new_n917), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n917), .A2(new_n918), .B1(new_n919), .B2(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n467), .A2(new_n916), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n920), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n910), .B1(new_n922), .B2(new_n694), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n206), .B2(new_n741), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n910), .A2(new_n922), .A3(new_n694), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n859), .B1(new_n924), .B2(new_n925), .ZN(G367));
  NOR2_X1   g0726(.A1(new_n670), .A2(new_n698), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n547), .A2(new_n557), .A3(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n928), .B(KEYINPUT107), .C1(new_n673), .C2(new_n927), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(KEYINPUT107), .B2(new_n928), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n748), .ZN(new_n931));
  INV_X1    g0731(.A(new_n326), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n754), .B1(new_n708), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n756), .A2(new_n235), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n745), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI22_X1  g0735(.A1(G50), .A2(new_n766), .B1(new_n783), .B2(G143), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n355), .B2(new_n839), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n770), .A2(new_n290), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n250), .B1(new_n838), .B2(new_n773), .C1(new_n781), .C2(new_n201), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n202), .A2(new_n779), .B1(new_n786), .B2(new_n218), .ZN(new_n940));
  NOR4_X1   g0740(.A1(new_n937), .A2(new_n938), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT111), .Z(new_n942));
  NAND2_X1  g0742(.A1(new_n780), .A2(G116), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT46), .Z(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(G303), .B2(new_n769), .ZN(new_n945));
  INV_X1    g0745(.A(G317), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n259), .B1(new_n946), .B2(new_n773), .C1(new_n786), .C2(new_n473), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT110), .Z(new_n948));
  AOI22_X1  g0748(.A1(G283), .A2(new_n766), .B1(new_n783), .B2(G311), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n765), .A2(G294), .B1(G107), .B2(new_n778), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n945), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n942), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT112), .Z(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT47), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n931), .B(new_n935), .C1(new_n954), .C2(new_n752), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n521), .B(new_n529), .C1(new_n487), .C2(new_n698), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n675), .A2(new_n527), .A3(new_n691), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n706), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT45), .Z(new_n961));
  NOR2_X1   g0761(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n962));
  INV_X1    g0762(.A(new_n706), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n962), .B1(new_n963), .B2(new_n958), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n706), .B(new_n959), .C1(KEYINPUT108), .C2(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g0765(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n704), .A2(new_n961), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n704), .B1(new_n961), .B2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n701), .A2(new_n705), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT109), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n702), .B1(new_n678), .B2(new_n698), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(KEYINPUT109), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n808), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n739), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n739), .B1(new_n971), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n709), .B(KEYINPUT41), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n743), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT43), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n930), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n972), .A2(new_n959), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n529), .B1(new_n956), .B2(new_n610), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n985), .A2(KEYINPUT42), .B1(new_n698), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n984), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n930), .A2(new_n983), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n704), .A2(new_n958), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n955), .B1(new_n982), .B2(new_n995), .ZN(G387));
  OR2_X1    g0796(.A1(new_n702), .A2(new_n749), .ZN(new_n997));
  INV_X1    g0797(.A(new_n711), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n759), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(G107), .B2(new_n210), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n232), .A2(new_n262), .ZN(new_n1001));
  AOI211_X1 g0801(.A(G45), .B(new_n998), .C1(G68), .C2(G77), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n288), .A2(G50), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n708), .B(new_n250), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1000), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n744), .B1(new_n1006), .B2(new_n755), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n259), .B1(new_n774), .B2(G150), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n218), .B2(new_n781), .C1(new_n789), .C2(new_n473), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT113), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G68), .A2(new_n766), .B1(new_n765), .B2(new_n329), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT114), .Z(new_n1012));
  NOR2_X1   g0812(.A1(new_n779), .A2(new_n326), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n770), .B2(new_n240), .C1(new_n355), .C2(new_n784), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n1010), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n250), .B1(new_n774), .B2(G326), .ZN(new_n1017));
  INV_X1    g0817(.A(G283), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n781), .A2(new_n797), .B1(new_n779), .B2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G311), .A2(new_n765), .B1(new_n783), .B2(G322), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n798), .B2(new_n832), .C1(new_n946), .C2(new_n770), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT48), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n1022), .B2(new_n1021), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT49), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1017), .B1(new_n538), .B2(new_n786), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1016), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT115), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n752), .B1(new_n1028), .B2(KEYINPUT115), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1007), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n977), .A2(new_n743), .B1(new_n997), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n978), .A2(new_n709), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n739), .A2(new_n977), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(G393));
  AOI21_X1  g0835(.A(new_n754), .B1(G97), .B2(new_n708), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n756), .A2(new_n239), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n745), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n250), .B1(new_n774), .B2(G322), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n779), .B2(new_n538), .C1(new_n1018), .C2(new_n781), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n797), .A2(new_n832), .B1(new_n839), .B2(new_n798), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G107), .C2(new_n794), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G311), .A2(new_n769), .B1(new_n783), .B2(G317), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  AOI22_X1  g0844(.A1(G150), .A2(new_n783), .B1(new_n769), .B2(G159), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT51), .Z(new_n1046));
  NOR2_X1   g0846(.A1(new_n779), .A2(new_n416), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n259), .B(new_n1047), .C1(G143), .C2(new_n774), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n202), .B2(new_n781), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n240), .A2(new_n839), .B1(new_n832), .B2(new_n288), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1049), .A2(new_n834), .A3(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1042), .A2(new_n1044), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1038), .B1(new_n752), .B2(new_n1052), .C1(new_n958), .C2(new_n749), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n971), .A2(new_n978), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n709), .B1(new_n971), .B2(new_n978), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1053), .B1(new_n742), .B2(new_n971), .C1(new_n1054), .C2(new_n1055), .ZN(G390));
  NAND2_X1  g0856(.A1(new_n904), .A2(new_n816), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n895), .B1(new_n1057), .B2(new_n902), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n892), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n732), .A2(new_n818), .A3(new_n902), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n883), .A2(new_n894), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1059), .B(new_n1060), .C1(new_n1061), .C2(new_n1058), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n916), .A2(G330), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n1063), .A2(new_n817), .A3(new_n903), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1058), .B1(new_n883), .B2(new_n894), .ZN(new_n1065));
  AOI21_X1  g0865(.A(KEYINPUT38), .B1(new_n886), .B2(new_n889), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n871), .A2(new_n385), .A3(new_n873), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1067), .A2(new_n868), .B1(new_n865), .B2(KEYINPUT37), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n864), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n413), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1066), .B1(new_n1070), .B2(KEYINPUT38), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n905), .A2(new_n1071), .A3(new_n895), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1064), .B1(new_n1065), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1062), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n742), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1061), .A2(new_n747), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n744), .B1(new_n329), .B2(new_n847), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n259), .B1(new_n774), .B2(G125), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n779), .B2(new_n355), .C1(new_n240), .C2(new_n786), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G132), .A2(new_n769), .B1(new_n765), .B2(G137), .ZN(new_n1080));
  INV_X1    g0880(.A(G128), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT54), .B(G143), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n784), .C1(new_n832), .C2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT53), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n781), .B2(new_n290), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n780), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1079), .B(new_n1083), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT116), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G107), .A2(new_n765), .B1(new_n769), .B2(G116), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n473), .B2(new_n832), .C1(new_n1018), .C2(new_n784), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n259), .B1(new_n797), .B2(new_n773), .C1(new_n781), .C2(new_n550), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n1090), .A2(new_n844), .A3(new_n1047), .A4(new_n1091), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT117), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n752), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1077), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1075), .B1(new_n1076), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n902), .B1(new_n732), .B2(new_n818), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1057), .B1(new_n1099), .B2(new_n1064), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1057), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n903), .B1(new_n1063), .B2(new_n817), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1060), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1063), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n467), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n908), .A2(new_n665), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1074), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1062), .A2(new_n1111), .A3(new_n1073), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n709), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1098), .A2(new_n1113), .ZN(G378));
  XOR2_X1   g0914(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n296), .A2(new_n863), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT55), .Z(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n317), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n317), .A2(new_n1119), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1116), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1122), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1124), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT40), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n882), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n413), .A2(new_n1069), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT38), .B1(new_n1130), .B2(new_n875), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1128), .B(new_n917), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n911), .A2(new_n916), .ZN(new_n1133));
  OAI21_X1  g0933(.A(KEYINPUT40), .B1(new_n1071), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1127), .B1(new_n1135), .B2(G330), .ZN(new_n1136));
  INV_X1    g0936(.A(G330), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1137), .B(new_n1126), .C1(new_n1132), .C2(new_n1134), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n907), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1126), .B1(new_n920), .B2(new_n1137), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n907), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1135), .A2(new_n1127), .A3(G330), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT120), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1139), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n1112), .B2(new_n1108), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1140), .A2(KEYINPUT120), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1139), .A2(new_n1143), .B1(new_n1112), .B2(new_n1108), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n709), .C1(KEYINPUT57), .C2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1136), .A2(new_n1138), .A3(new_n907), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1141), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n743), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1126), .A2(new_n746), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n744), .B1(G50), .B2(new_n847), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n781), .A2(new_n1082), .B1(new_n779), .B2(new_n290), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G125), .A2(new_n783), .B1(new_n769), .B2(G128), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n838), .B2(new_n832), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(G132), .C2(new_n765), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT59), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n785), .A2(G159), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n774), .C2(G124), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n786), .A2(new_n201), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n250), .A2(G41), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n1018), .B2(new_n773), .C1(new_n779), .C2(new_n202), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(new_n219), .C2(new_n780), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n326), .B2(new_n832), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G107), .A2(new_n769), .B1(new_n783), .B2(G116), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n473), .B2(new_n839), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT58), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1175), .A2(KEYINPUT58), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1169), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n240), .C1(G33), .C2(G41), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1167), .A2(new_n1176), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1157), .B1(new_n1180), .B2(new_n751), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1156), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1154), .A2(new_n1155), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n742), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1182), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT119), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1151), .A2(new_n1187), .ZN(G375));
  NAND2_X1  g0988(.A1(new_n903), .A2(new_n746), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n744), .B1(G68), .B2(new_n847), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n769), .A2(G137), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n839), .B2(new_n1082), .C1(new_n842), .C2(new_n784), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT123), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n250), .B1(new_n773), .B2(new_n1081), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1194), .B(new_n1168), .C1(G159), .C2(new_n780), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n766), .A2(G150), .B1(G50), .B2(new_n778), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT124), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1192), .B2(KEYINPUT123), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n781), .A2(new_n473), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1014), .B(new_n259), .C1(new_n798), .C2(new_n773), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G294), .C2(new_n783), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n468), .A2(new_n832), .B1(new_n839), .B2(new_n538), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT122), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n794), .A2(G77), .B1(G283), .B2(new_n769), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1202), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1196), .A2(new_n1199), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1190), .B1(new_n1209), .B2(new_n751), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1104), .A2(new_n743), .B1(new_n1189), .B2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n980), .B(KEYINPUT121), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1109), .A2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1211), .B1(new_n1213), .B2(new_n1214), .ZN(G381));
  NOR2_X1   g1015(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1053), .B1(new_n971), .B2(new_n742), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(G384), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(G393), .A2(G396), .A3(G381), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  OR4_X1    g1021(.A1(G387), .A2(new_n1221), .A3(G375), .A4(G378), .ZN(G407));
  INV_X1    g1022(.A(G378), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n690), .A2(G213), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT125), .Z(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(G407), .B(G213), .C1(G375), .C2(new_n1226), .ZN(G409));
  NAND2_X1  g1027(.A1(new_n1225), .A2(G2897), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1100), .A2(new_n1107), .A3(KEYINPUT60), .A4(new_n1103), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1109), .A2(new_n709), .A3(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT60), .B1(new_n1231), .B2(new_n1107), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1211), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1219), .ZN(new_n1234));
  OAI211_X1 g1034(.A(G384), .B(new_n1211), .C1(new_n1232), .C2(new_n1230), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT126), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1228), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1228), .ZN(new_n1239));
  AOI211_X1 g1039(.A(KEYINPUT126), .B(new_n1239), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1238), .A2(new_n1240), .B1(new_n1237), .B2(new_n1236), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1151), .A2(new_n1187), .A3(G378), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1150), .A2(new_n1212), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1145), .A2(new_n743), .A3(new_n1148), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n1182), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1223), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1225), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT61), .B1(new_n1242), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1250), .B2(new_n1236), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G390), .B(new_n955), .C1(new_n982), .C2(new_n995), .ZN(new_n1254));
  XOR2_X1   g1054(.A(G393), .B(G396), .Z(new_n1255));
  NAND2_X1  g1055(.A1(G387), .A2(new_n1218), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1225), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1236), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1251), .A2(new_n1253), .A3(new_n1259), .A4(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1260), .A2(new_n1264), .A3(new_n1261), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT61), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1260), .B2(new_n1241), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1264), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1265), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1263), .B1(new_n1269), .B2(new_n1259), .ZN(G405));
  INV_X1    g1070(.A(new_n1243), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G378), .B1(new_n1151), .B2(new_n1187), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1261), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1261), .A2(new_n1274), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1236), .A2(KEYINPUT127), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1276), .B(new_n1277), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1275), .A2(new_n1259), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1259), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(G402));
endmodule


