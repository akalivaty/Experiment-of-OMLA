//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(KEYINPUT64), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n466), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n463), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  AND3_X1   g051(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(KEYINPUT3), .B1(new_n470), .B2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(new_n463), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n481), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n469), .B2(new_n471), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT4), .B1(new_n490), .B2(new_n468), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n469), .B2(new_n471), .ZN(new_n494));
  NAND2_X1  g069(.A1(G102), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n463), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT4), .B1(new_n461), .B2(G138), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n492), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT5), .B1(new_n502), .B2(KEYINPUT65), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(G543), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n507), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n513), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(new_n512), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT66), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT66), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n519), .B(new_n524), .C1(new_n520), .C2(new_n512), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n507), .A2(new_n508), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n525), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n523), .A2(new_n530), .ZN(G168));
  XNOR2_X1  g106(.A(KEYINPUT67), .B(G90), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n503), .A2(new_n506), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n508), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G52), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n533), .A2(new_n538), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n509), .A2(new_n543), .B1(new_n544), .B2(new_n512), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n507), .A2(G56), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n514), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT68), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT69), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT71), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n503), .A2(new_n506), .A3(G65), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n557), .B1(new_n560), .B2(G651), .ZN(new_n561));
  AOI211_X1 g136(.A(KEYINPUT71), .B(new_n514), .C1(new_n558), .C2(new_n559), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT6), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n564), .A2(new_n566), .A3(G53), .A4(G543), .ZN(new_n567));
  AND2_X1   g142(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n568));
  NOR2_X1   g143(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n508), .A2(G53), .A3(G543), .A4(new_n568), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n508), .A2(G91), .A3(new_n503), .A4(new_n506), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n563), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n539), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(G87), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n509), .ZN(G288));
  AOI22_X1  g156(.A1(new_n528), .A2(G86), .B1(G48), .B2(new_n539), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n503), .A2(new_n506), .A3(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n514), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT72), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n582), .A2(new_n587), .A3(new_n588), .ZN(G305));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n509), .A2(new_n590), .B1(new_n591), .B2(new_n512), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n507), .A2(G60), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n514), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n507), .A2(G92), .A3(new_n508), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  XOR2_X1   g177(.A(KEYINPUT73), .B(G66), .Z(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n535), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(G54), .B2(new_n539), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G299), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G168), .B2(new_n610), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(G168), .B2(new_n610), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  INV_X1    g190(.A(new_n549), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n610), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n606), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n480), .A2(G135), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n482), .A2(G123), .ZN(new_n622));
  NOR2_X1   g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND3_X1  g201(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT74), .B(G2100), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT75), .Z(G156));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XOR2_X1   g210(.A(G1341), .B(G1348), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT76), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n639), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT77), .B(KEYINPUT18), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  MUX2_X1   g234(.A(new_n656), .B(new_n651), .S(new_n659), .Z(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n664), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(G1986), .Z(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  INV_X1    g252(.A(G1981), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G24), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n596), .B2(new_n681), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1986), .ZN(new_n684));
  INV_X1    g259(.A(G29), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G25), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n480), .A2(G131), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n482), .A2(G119), .ZN(new_n688));
  OR2_X1    g263(.A1(G95), .A2(G2105), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n689), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n686), .B1(new_n692), .B2(new_n685), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT35), .B(G1991), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT78), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n693), .B(new_n695), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n681), .A2(G6), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n507), .A2(G86), .A3(new_n508), .ZN(new_n698));
  INV_X1    g273(.A(G48), .ZN(new_n699));
  OAI221_X1 g274(.A(new_n698), .B1(new_n699), .B2(new_n512), .C1(new_n585), .C2(new_n586), .ZN(new_n700));
  INV_X1    g275(.A(new_n588), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n697), .B1(new_n702), .B2(new_n681), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT80), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  MUX2_X1   g283(.A(G23), .B(G288), .S(G16), .Z(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT81), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n709), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n681), .A2(G22), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G166), .B2(new_n681), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(G1971), .Z(new_n715));
  NAND4_X1  g290(.A1(new_n707), .A2(new_n708), .A3(new_n712), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT79), .B(KEYINPUT34), .Z(new_n717));
  AOI211_X1 g292(.A(new_n684), .B(new_n696), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT36), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n718), .A2(new_n722), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n685), .A2(G32), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n480), .A2(G141), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n482), .A2(G129), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT87), .B(KEYINPUT26), .Z(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n726), .A2(new_n727), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n725), .B1(new_n733), .B2(new_n685), .ZN(new_n734));
  INV_X1    g309(.A(G1996), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT88), .B(KEYINPUT27), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT31), .B(G11), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT89), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G28), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n685), .B1(new_n741), .B2(G28), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n740), .B1(new_n742), .B2(new_n743), .C1(new_n625), .C2(new_n685), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT90), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n681), .A2(G21), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G168), .B2(new_n681), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(G1966), .ZN(new_n748));
  NAND2_X1  g323(.A1(G164), .A2(G29), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G27), .B2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G2078), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n745), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n681), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n549), .B2(new_n681), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT83), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1341), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n681), .A2(G20), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT23), .ZN(new_n759));
  INV_X1    g334(.A(G299), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n681), .ZN(new_n761));
  INV_X1    g336(.A(G1956), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n738), .A2(new_n753), .A3(new_n757), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n681), .A2(G4), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n607), .B2(new_n681), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT82), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1348), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n685), .A2(G35), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G162), .B2(new_n685), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT29), .B(G2090), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n681), .A2(G5), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G171), .B2(new_n681), .ZN(new_n774));
  INV_X1    g349(.A(G1961), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n750), .A2(new_n751), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n747), .A2(G1966), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n772), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n685), .A2(G26), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT86), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT28), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n480), .A2(G140), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT84), .ZN(new_n784));
  OR2_X1    g359(.A1(G104), .A2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n785), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT85), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G128), .B2(new_n482), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n782), .B1(new_n789), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT24), .ZN(new_n792));
  INV_X1    g367(.A(G34), .ZN(new_n793));
  AOI21_X1  g368(.A(G29), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G160), .B2(new_n685), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G2084), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n685), .A2(G33), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n480), .A2(G139), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT25), .Z(new_n802));
  AOI22_X1  g377(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n800), .B(new_n802), .C1(new_n463), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n799), .B1(new_n804), .B2(G29), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n797), .A2(new_n798), .B1(new_n806), .B2(G2072), .ZN(new_n807));
  INV_X1    g382(.A(G2072), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n796), .A2(G2084), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n791), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n764), .A2(new_n768), .A3(new_n779), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n724), .A2(new_n811), .ZN(G150));
  INV_X1    g387(.A(G150), .ZN(G311));
  AOI22_X1  g388(.A1(new_n528), .A2(G93), .B1(G55), .B2(new_n539), .ZN(new_n814));
  NAND2_X1  g389(.A1(G80), .A2(G543), .ZN(new_n815));
  INV_X1    g390(.A(G67), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n535), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G651), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT92), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n819), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NOR2_X1   g401(.A1(new_n606), .A2(new_n614), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n616), .B1(new_n821), .B2(new_n822), .ZN(new_n830));
  INV_X1    g405(.A(new_n822), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n831), .A2(new_n549), .A3(new_n820), .A4(new_n814), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n829), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT93), .Z(new_n836));
  AOI21_X1  g411(.A(G860), .B1(new_n834), .B2(KEYINPUT39), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n836), .A2(KEYINPUT94), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(KEYINPUT94), .B1(new_n836), .B2(new_n837), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n826), .B1(new_n838), .B2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(new_n500), .B(KEYINPUT95), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n804), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n480), .A2(G142), .ZN(new_n843));
  NOR2_X1   g418(.A1(G106), .A2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n482), .A2(KEYINPUT96), .A3(G130), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT96), .B1(new_n482), .B2(G130), .ZN(new_n847));
  OAI221_X1 g422(.A(new_n843), .B1(new_n844), .B2(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n628), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n842), .B(new_n849), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n789), .B(new_n732), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n692), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n851), .B(new_n691), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n842), .B(new_n849), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(G160), .B(new_n625), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G162), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n858), .B1(new_n853), .B2(new_n856), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT97), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n864), .A2(new_n865), .A3(new_n860), .A4(new_n859), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT40), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(new_n866), .A3(KEYINPUT40), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(G395));
  XNOR2_X1  g446(.A(G166), .B(KEYINPUT101), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n702), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n596), .B(G288), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n873), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT42), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n830), .A2(new_n879), .A3(new_n832), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n879), .B1(new_n830), .B2(new_n832), .ZN(new_n882));
  OAI22_X1  g457(.A1(new_n881), .A2(new_n882), .B1(G559), .B2(new_n606), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n618), .A3(new_n880), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n760), .A2(new_n606), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n607), .A2(G299), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(KEYINPUT99), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT41), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n886), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n883), .A2(new_n885), .A3(new_n889), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n886), .A2(KEYINPUT100), .A3(new_n891), .A4(new_n895), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT102), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n898), .A2(new_n899), .A3(new_n903), .A4(new_n900), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n878), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n877), .B1(KEYINPUT102), .B2(new_n901), .ZN(new_n906));
  OAI21_X1  g481(.A(G868), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n824), .A2(new_n610), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(G295));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n908), .ZN(G331));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n911));
  INV_X1    g486(.A(new_n530), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(new_n522), .A3(G301), .ZN(new_n913));
  OAI21_X1  g488(.A(G171), .B1(new_n523), .B2(new_n530), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n915), .A2(new_n833), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n833), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n889), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n892), .A2(new_n894), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n920), .B2(new_n918), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n876), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n873), .B(new_n874), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n895), .A2(new_n891), .A3(new_n916), .A4(new_n917), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n919), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n922), .A2(new_n925), .A3(new_n926), .A4(new_n860), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(new_n860), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(new_n919), .B2(new_n924), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n927), .A2(new_n928), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n911), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n922), .A2(new_n925), .A3(new_n860), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(new_n926), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT44), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n939), .ZN(G397));
  INV_X1    g515(.A(G2067), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n789), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n735), .B2(new_n733), .ZN(new_n943));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT45), .B1(new_n500), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n474), .A2(G40), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(new_n464), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT104), .Z(new_n949));
  NAND2_X1  g524(.A1(new_n943), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n948), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n735), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n732), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n691), .B(new_n695), .Z(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(new_n949), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n596), .B(G1986), .Z(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n951), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n500), .A2(new_n944), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT50), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n500), .A2(new_n961), .A3(new_n944), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n960), .A2(new_n798), .A3(new_n947), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  INV_X1    g541(.A(new_n493), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n477), .B2(new_n478), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n495), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n498), .B1(new_n969), .B2(new_n463), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n970), .B2(new_n492), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n966), .B(new_n947), .C1(new_n971), .C2(KEYINPUT45), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n474), .A2(G40), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n465), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT110), .B1(new_n945), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n965), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(G168), .B(new_n963), .C1(new_n976), .C2(G1966), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(KEYINPUT120), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n979), .A2(KEYINPUT120), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n977), .A2(new_n980), .A3(new_n982), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n963), .B1(new_n976), .B2(G1966), .ZN(new_n986));
  NOR2_X1   g561(.A1(G168), .A2(new_n978), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n965), .A2(new_n945), .A3(new_n974), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n960), .A2(new_n947), .A3(new_n962), .ZN(new_n990));
  OAI22_X1  g565(.A1(new_n989), .A2(G1971), .B1(new_n990), .B2(G2090), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT55), .B(G8), .C1(new_n513), .C2(new_n517), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n992), .A2(KEYINPUT105), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G166), .B2(new_n978), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(KEYINPUT105), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(G8), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT106), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n991), .A2(new_n1000), .A3(new_n997), .A4(G8), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n947), .A2(new_n944), .A3(new_n500), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT107), .B(G1976), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(G288), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n528), .A2(G87), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1006), .A2(G1976), .A3(new_n579), .A4(new_n578), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1003), .A2(new_n1005), .A3(G8), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT108), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n978), .B1(new_n971), .B2(new_n947), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n1007), .A4(new_n1005), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1007), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT52), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n582), .A2(new_n587), .A3(new_n678), .A4(new_n588), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n698), .B1(new_n699), .B2(new_n512), .ZN(new_n1017));
  OAI21_X1  g592(.A(G1981), .B1(new_n1017), .B2(new_n585), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1016), .A2(KEYINPUT49), .A3(new_n1018), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1010), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1013), .A2(new_n1015), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n997), .B1(new_n991), .B2(G8), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n959), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1029), .A2(new_n751), .A3(new_n964), .A4(new_n947), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1027), .A2(new_n1030), .B1(new_n990), .B2(new_n775), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n972), .A2(new_n975), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n964), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n751), .A2(KEYINPUT53), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(G301), .B(KEYINPUT54), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G113), .A2(G2104), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT3), .B(G2104), .Z(new_n1038));
  INV_X1    g613(.A(G125), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n463), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n462), .A2(KEYINPUT121), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n973), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT122), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(KEYINPUT122), .A3(new_n973), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT123), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT53), .B1(new_n1049), .B2(new_n751), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n1049), .B2(new_n751), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1047), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n965), .A2(new_n945), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1036), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1035), .A2(new_n1036), .B1(new_n1031), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1002), .A2(new_n1026), .A3(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n988), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(KEYINPUT57), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n574), .B(new_n1060), .C1(new_n561), .C2(new_n562), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(KEYINPUT57), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n962), .A2(new_n947), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n961), .B1(new_n500), .B2(new_n944), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n762), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT56), .B(G2072), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1029), .A2(new_n964), .A3(new_n947), .A4(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1066), .A2(new_n1069), .A3(KEYINPUT113), .A4(new_n1071), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1066), .A2(KEYINPUT115), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1069), .A2(KEYINPUT114), .A3(new_n1071), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT114), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1348), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n990), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n971), .A2(new_n941), .A3(new_n947), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n606), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1076), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1072), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1066), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(KEYINPUT61), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1089), .A2(KEYINPUT61), .B1(new_n1076), .B2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1029), .A2(new_n735), .A3(new_n964), .A4(new_n947), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(G1341), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1003), .A2(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1093), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1094), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n549), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT119), .B1(new_n1101), .B2(KEYINPUT59), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1085), .A2(new_n606), .A3(new_n1086), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT60), .B1(new_n1104), .B2(new_n1087), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1085), .A2(new_n1086), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1102), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n549), .B(new_n1108), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1088), .B1(new_n1092), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1057), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1025), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n978), .A2(KEYINPUT63), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1113), .A2(G168), .A3(new_n986), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1024), .B1(new_n1115), .B2(new_n1002), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n991), .A2(G8), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT111), .ZN(new_n1119));
  INV_X1    g694(.A(new_n997), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT111), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n991), .A2(new_n1121), .A3(G8), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n986), .A2(G168), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1013), .A2(G8), .A3(new_n1015), .A4(new_n1023), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1117), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G288), .A2(G1976), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1023), .A2(new_n1128), .B1(new_n678), .B2(new_n702), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1010), .B1(new_n1129), .B2(KEYINPUT109), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(KEYINPUT109), .B2(new_n1129), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1116), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1002), .A2(G171), .A3(new_n1026), .A4(new_n1035), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n986), .A2(new_n987), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n977), .A2(new_n980), .A3(new_n982), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n982), .B1(new_n977), .B2(new_n980), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT62), .B(new_n1134), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1133), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1112), .B(new_n1132), .C1(new_n1141), .C2(KEYINPUT124), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1143), .B(new_n1133), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n958), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n948), .A2(G1986), .A3(G290), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT48), .Z(new_n1147));
  NAND2_X1  g722(.A1(new_n955), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n942), .A2(new_n733), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n949), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT126), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT47), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n952), .B(KEYINPUT46), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1152), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1148), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n692), .A2(new_n695), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n953), .A2(new_n1157), .B1(G2067), .B2(new_n789), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1156), .B1(new_n949), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1145), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g737(.A1(new_n864), .A2(new_n860), .A3(new_n859), .ZN(new_n1164));
  NOR3_X1   g738(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1165));
  XOR2_X1   g739(.A(new_n1165), .B(KEYINPUT127), .Z(new_n1166));
  NOR2_X1   g740(.A1(new_n1166), .A2(G229), .ZN(new_n1167));
  OAI211_X1 g741(.A(new_n1164), .B(new_n1167), .C1(new_n933), .C2(new_n934), .ZN(G225));
  INV_X1    g742(.A(G225), .ZN(G308));
endmodule


