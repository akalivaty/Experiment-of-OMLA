//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1199, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G97), .C2(G257), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G1), .B2(G20), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT1), .Z(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NOR3_X1   g0025(.A1(new_n217), .A2(new_n221), .A3(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n228), .B(new_n229), .Z(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n230), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G68), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  XOR2_X1   g0044(.A(KEYINPUT8), .B(G58), .Z(new_n245));
  NAND2_X1  g0045(.A1(new_n219), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n245), .A2(new_n247), .B1(G20), .B2(new_n203), .ZN(new_n248));
  INV_X1    g0048(.A(G150), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n248), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(KEYINPUT69), .B1(new_n222), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT69), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n255), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n220), .A3(new_n256), .ZN(new_n257));
  AND3_X1   g0057(.A1(new_n254), .A2(new_n220), .A3(new_n256), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT68), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT68), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n252), .A2(new_n257), .B1(G50), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(G50), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(G222), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G223), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(new_n277), .B2(new_n275), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n253), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n278), .B(new_n279), .C1(G77), .C2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n287), .A2(new_n259), .A3(G274), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n263), .A2(new_n287), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT67), .B1(new_n253), .B2(new_n285), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT67), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G33), .A3(G41), .ZN(new_n292));
  INV_X1    g0092(.A(new_n220), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n288), .B1(new_n295), .B2(G226), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n284), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G200), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n269), .A2(new_n270), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n284), .A2(G190), .A3(new_n296), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n271), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n284), .A2(new_n305), .A3(new_n296), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n269), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT70), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n283), .A2(G232), .A3(new_n275), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n274), .A2(new_n213), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(G1698), .ZN(new_n312));
  INV_X1    g0112(.A(G107), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n312), .B1(new_n309), .B2(new_n310), .C1(new_n313), .C2(new_n283), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n279), .ZN(new_n315));
  INV_X1    g0115(.A(new_n288), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n295), .A2(G244), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n303), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  XOR2_X1   g0120(.A(KEYINPUT15), .B(G87), .Z(new_n321));
  AOI22_X1  g0121(.A1(new_n250), .A2(new_n245), .B1(new_n321), .B2(new_n247), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n219), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n257), .ZN(new_n325));
  INV_X1    g0125(.A(new_n268), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n323), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n266), .A2(G77), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n318), .B2(G179), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n320), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n318), .A2(G200), .ZN(new_n333));
  INV_X1    g0133(.A(new_n329), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(new_n318), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n308), .B1(KEYINPUT71), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(G226), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n283), .A2(KEYINPUT72), .A3(G226), .A4(new_n275), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n283), .A2(G232), .A3(G1698), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n279), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n295), .A2(G238), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n316), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n345), .A2(new_n279), .B1(G238), .B2(new_n295), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT13), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(new_n316), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n349), .A2(KEYINPUT74), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n349), .B1(KEYINPUT74), .B2(new_n352), .ZN(new_n354));
  OAI21_X1  g0154(.A(G190), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n247), .A2(G77), .B1(new_n250), .B2(G50), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n219), .B2(G68), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n357), .A2(new_n257), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(KEYINPUT11), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(KEYINPUT11), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n212), .C2(new_n265), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n268), .A2(G68), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT12), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n349), .A2(KEYINPUT73), .A3(new_n352), .ZN(new_n365));
  OR3_X1    g0165(.A1(new_n348), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(G200), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n355), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n364), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(new_n366), .A3(G169), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n372));
  OAI21_X1  g0172(.A(G179), .B1(new_n353), .B2(new_n354), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n365), .A2(new_n366), .A3(new_n374), .A4(G169), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n369), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT7), .B1(new_n274), .B2(new_n219), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n219), .A4(new_n282), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G58), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(new_n212), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n383), .B2(new_n201), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n250), .A2(G159), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n283), .B2(G20), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT75), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n379), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n274), .A2(KEYINPUT75), .A3(KEYINPUT7), .A4(new_n219), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n386), .B1(new_n394), .B2(G68), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n257), .B(new_n388), .C1(new_n395), .C2(KEYINPUT16), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n289), .A2(new_n294), .A3(G232), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT76), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n277), .A2(new_n275), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n211), .A2(G1698), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n272), .C2(new_n273), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n288), .B1(new_n404), .B2(new_n279), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n289), .A2(new_n294), .A3(KEYINPUT76), .A4(G232), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n399), .A2(new_n405), .A3(G190), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n265), .A2(new_n245), .ZN(new_n408));
  INV_X1    g0208(.A(new_n245), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n268), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n399), .A2(new_n405), .A3(new_n406), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G200), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n396), .A2(new_n407), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n414), .B(KEYINPUT17), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n303), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n399), .A2(new_n405), .A3(new_n305), .A4(new_n406), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT77), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n396), .A2(new_n411), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT77), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n420), .A2(KEYINPUT18), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT78), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(new_n425), .A3(new_n428), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n416), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n337), .A2(KEYINPUT71), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n338), .A2(new_n377), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n283), .A2(G238), .A3(new_n275), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n283), .A2(G244), .A3(G1698), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n436), .B(new_n437), .C1(new_n253), .C2(new_n207), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n279), .ZN(new_n439));
  INV_X1    g0239(.A(G250), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n263), .B2(G45), .ZN(new_n441));
  INV_X1    g0241(.A(G274), .ZN(new_n442));
  AOI211_X1 g0242(.A(new_n286), .B(new_n442), .C1(new_n260), .C2(new_n262), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n294), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n263), .A2(G33), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n258), .A2(new_n268), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n321), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n268), .A2(new_n321), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT19), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n219), .B1(new_n343), .B2(new_n451), .ZN(new_n452));
  NOR4_X1   g0252(.A1(KEYINPUT80), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT80), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G87), .A2(G97), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(new_n313), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n452), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n283), .A2(new_n219), .A3(G68), .ZN(new_n458));
  INV_X1    g0258(.A(G97), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n451), .B1(new_n246), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT81), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT81), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n451), .C1(new_n246), .C2(new_n459), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n457), .A2(new_n458), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n450), .B1(new_n464), .B2(new_n257), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n445), .A2(new_n305), .B1(new_n449), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(G169), .B2(new_n445), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n445), .A2(G190), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n258), .A2(G87), .A3(new_n268), .A4(new_n446), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G200), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n468), .B(new_n470), .C1(new_n471), .C2(new_n445), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n251), .A2(new_n323), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n394), .B2(G107), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT6), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n459), .A2(new_n313), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n313), .A2(KEYINPUT6), .A3(G97), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n219), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n258), .B1(new_n476), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n268), .A2(G97), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n459), .B2(new_n447), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n474), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n487), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n475), .B(new_n482), .C1(new_n394), .C2(G107), .ZN(new_n490));
  OAI211_X1 g0290(.A(KEYINPUT79), .B(new_n489), .C1(new_n490), .C2(new_n258), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n283), .A2(G250), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n275), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(G1698), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(G244), .C1(new_n273), .C2(new_n272), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  INV_X1    g0297(.A(G244), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n281), .B2(new_n282), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n496), .B(new_n497), .C1(new_n499), .C2(KEYINPUT4), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n279), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g0301(.A(KEYINPUT5), .B(G41), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n263), .A2(new_n502), .A3(G45), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n503), .A2(new_n294), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G257), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n443), .A2(new_n294), .A3(new_n502), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n507), .A2(G190), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n471), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n488), .A2(new_n491), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(G169), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n501), .A2(new_n505), .A3(G179), .A4(new_n506), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n394), .A2(G107), .ZN(new_n513));
  INV_X1    g0313(.A(new_n475), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n483), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n257), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n511), .A2(new_n512), .B1(new_n516), .B2(new_n489), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n473), .A2(new_n510), .A3(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G257), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n519));
  OAI211_X1 g0319(.A(G250), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G294), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n279), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n503), .A2(G264), .A3(new_n294), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n506), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(G190), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n524), .B(KEYINPUT85), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n523), .A2(new_n506), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n526), .B1(new_n529), .B2(new_n471), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n219), .B(G87), .C1(new_n272), .C2(new_n273), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT22), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT22), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n283), .A2(new_n534), .A3(new_n219), .A4(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n247), .A2(G116), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT23), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n538), .A2(new_n219), .A3(G107), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT23), .B1(new_n313), .B2(G20), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AND4_X1   g0342(.A1(new_n531), .A2(new_n536), .A3(new_n537), .A4(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n541), .B1(new_n533), .B2(new_n535), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n531), .B1(new_n544), .B2(new_n537), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n257), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n448), .A2(G107), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n326), .B(new_n313), .C1(KEYINPUT83), .C2(KEYINPUT25), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n326), .A2(KEYINPUT83), .A3(KEYINPUT25), .A4(new_n313), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n530), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n525), .A2(G169), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT84), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT85), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n524), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n504), .A2(KEYINPUT85), .A3(G264), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n528), .A2(G179), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT84), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n525), .A2(new_n561), .A3(G169), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n556), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT86), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT86), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n553), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n554), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n326), .A2(new_n207), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n258), .A2(G116), .A3(new_n268), .A4(new_n446), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n207), .A2(G20), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n497), .B(new_n219), .C1(G33), .C2(new_n459), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n257), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT20), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n569), .B(new_n570), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G264), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT82), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT82), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n283), .A2(new_n580), .A3(G264), .A4(G1698), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n283), .A2(G257), .A3(new_n275), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n274), .A2(G303), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n579), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n279), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n504), .A2(G270), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n506), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n577), .A2(new_n587), .A3(G169), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n587), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(G179), .A3(new_n577), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n577), .A2(new_n587), .A3(KEYINPUT21), .A4(G169), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n587), .A2(G200), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n335), .B2(new_n587), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n596), .A2(new_n577), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n435), .A2(new_n518), .A3(new_n568), .A4(new_n598), .ZN(G372));
  INV_X1    g0399(.A(KEYINPUT92), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n376), .A2(new_n370), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n368), .A2(new_n331), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n603), .A2(KEYINPUT91), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(KEYINPUT91), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n415), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n429), .A2(new_n424), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n302), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n600), .B(new_n307), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n606), .B2(new_n607), .ZN(new_n611));
  INV_X1    g0411(.A(new_n307), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT92), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n517), .ZN(new_n615));
  XNOR2_X1  g0415(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n473), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n444), .A2(KEYINPUT87), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT87), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n619), .B(new_n294), .C1(new_n441), .C2(new_n443), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n439), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G200), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n464), .A2(new_n257), .ZN(new_n623));
  INV_X1    g0423(.A(new_n450), .ZN(new_n624));
  AND4_X1   g0424(.A1(KEYINPUT88), .A2(new_n623), .A3(new_n624), .A4(new_n469), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT88), .B1(new_n465), .B2(new_n469), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT89), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT89), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n629), .B(new_n622), .C1(new_n625), .C2(new_n626), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n468), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n621), .A2(new_n303), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n466), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n511), .A2(new_n512), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n488), .A2(new_n634), .A3(new_n491), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n631), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n617), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n564), .A2(new_n592), .A3(new_n590), .A4(new_n593), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n488), .A2(new_n491), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n508), .A2(new_n509), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n517), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n554), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n631), .A2(new_n639), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n633), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n435), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n614), .A2(new_n647), .ZN(G369));
  INV_X1    g0448(.A(new_n553), .ZN(new_n649));
  INV_X1    g0449(.A(new_n263), .ZN(new_n650));
  INV_X1    g0450(.A(G13), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(G20), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OR3_X1    g0453(.A1(new_n650), .A2(KEYINPUT27), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT27), .B1(new_n650), .B2(new_n653), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n568), .B1(new_n649), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n553), .A2(new_n563), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT94), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT94), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n660), .A2(new_n664), .A3(new_n661), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n594), .A2(new_n658), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n553), .A2(new_n563), .A3(new_n659), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n666), .ZN(new_n671));
  INV_X1    g0471(.A(new_n594), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n577), .A2(new_n658), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n673), .B(KEYINPUT93), .Z(new_n674));
  MUX2_X1   g0474(.A(new_n598), .B(new_n672), .S(new_n674), .Z(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT95), .Z(G399));
  NOR2_X1   g0479(.A1(new_n453), .A2(new_n456), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n207), .ZN(new_n681));
  INV_X1    g0481(.A(new_n223), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n681), .A2(new_n259), .A3(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT96), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT96), .ZN(new_n686));
  INV_X1    g0486(.A(new_n683), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n685), .B(new_n686), .C1(new_n218), .C2(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n518), .A2(new_n598), .A3(new_n568), .A4(new_n659), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT98), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND4_X1   g0493(.A1(new_n445), .A2(new_n523), .A3(new_n527), .A4(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n512), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(new_n591), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n691), .B2(new_n692), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n691), .A2(new_n692), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n694), .A2(new_n695), .A3(new_n591), .A4(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n621), .A2(new_n305), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n529), .A2(KEYINPUT97), .A3(new_n507), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT97), .B1(new_n529), .B2(new_n507), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n587), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n697), .B(new_n699), .C1(new_n700), .C2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n658), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n690), .A2(new_n705), .A3(KEYINPUT31), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n707), .A3(new_n658), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  INV_X1    g0510(.A(new_n633), .ZN(new_n711));
  AND4_X1   g0511(.A1(KEYINPUT26), .A2(new_n488), .A3(new_n634), .A4(new_n491), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n631), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n616), .B1(new_n473), .B2(new_n615), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n553), .A2(new_n563), .A3(new_n566), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n566), .B1(new_n553), .B2(new_n563), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n594), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n642), .A3(new_n643), .A4(new_n631), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n658), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n646), .A2(new_n659), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(KEYINPUT29), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n710), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n689), .B1(new_n725), .B2(G1), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT99), .ZN(G364));
  AOI21_X1  g0527(.A(new_n259), .B1(new_n652), .B2(G45), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n683), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n676), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n675), .A2(G330), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n293), .B1(new_n219), .B2(G169), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT100), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n219), .A2(G190), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G159), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT32), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n274), .B1(new_n742), .B2(KEYINPUT32), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n305), .A2(new_n471), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n738), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G68), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n219), .B1(new_n739), .B2(G190), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G97), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n743), .A2(new_n744), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n219), .A2(new_n335), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(new_n305), .A3(G200), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n745), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n755), .A2(G87), .B1(new_n757), .B2(G50), .ZN(new_n758));
  NOR4_X1   g0558(.A1(new_n219), .A2(new_n471), .A3(G179), .A4(G190), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT102), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(KEYINPUT102), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n305), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n753), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT101), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n764), .A2(new_n765), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n758), .B1(new_n762), .B2(new_n313), .C1(new_n382), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n763), .A2(new_n738), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n752), .B(new_n770), .C1(G77), .C2(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G311), .A2(new_n772), .B1(new_n741), .B2(G329), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n757), .A2(G326), .ZN(new_n775));
  INV_X1    g0575(.A(G317), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(KEYINPUT33), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n776), .A2(KEYINPUT33), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n747), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n283), .B1(new_n750), .B2(G294), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n774), .A2(new_n775), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n769), .B1(new_n762), .B2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n781), .B(new_n784), .C1(G303), .C2(new_n755), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n737), .B1(new_n773), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n682), .A2(new_n283), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n218), .A2(G45), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(new_n240), .C2(new_n286), .ZN(new_n789));
  INV_X1    g0589(.A(G355), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n283), .A2(new_n223), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(G116), .B2(new_n223), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n737), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n795), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n786), .B(new_n797), .C1(new_n675), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n730), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n734), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT103), .Z(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NOR3_X1   g0603(.A1(new_n320), .A2(new_n330), .A3(new_n658), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n329), .A2(new_n658), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n336), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n804), .B1(new_n332), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n723), .B(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(new_n710), .Z(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n731), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G150), .A2(new_n747), .B1(new_n772), .B2(G159), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  INV_X1    g0612(.A(G143), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(new_n812), .B2(new_n756), .C1(new_n769), .C2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT34), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n283), .B1(new_n749), .B2(new_n382), .C1(new_n816), .C2(new_n740), .ZN(new_n817));
  INV_X1    g0617(.A(new_n762), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(G68), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n815), .B(new_n819), .C1(new_n202), .C2(new_n754), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n757), .A2(G303), .B1(new_n741), .B2(G311), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n821), .B1(new_n207), .B2(new_n771), .C1(new_n783), .C2(new_n746), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G97), .B2(new_n750), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n818), .A2(G87), .ZN(new_n824));
  INV_X1    g0624(.A(new_n769), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G294), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n283), .B1(new_n755), .B2(G107), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n823), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n736), .B1(new_n820), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n737), .A2(new_n793), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(new_n323), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n831), .B(new_n730), .C1(new_n807), .C2(new_n794), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n810), .A2(new_n832), .ZN(G384));
  INV_X1    g0633(.A(KEYINPUT40), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT16), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n212), .B1(new_n390), .B2(new_n379), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n386), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(new_n257), .A3(new_n388), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n411), .ZN(new_n840));
  INV_X1    g0640(.A(new_n656), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n430), .A2(new_n431), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n415), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n422), .B1(new_n417), .B2(new_n418), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n408), .A2(new_n410), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n390), .A2(new_n379), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n386), .B1(new_n847), .B2(G68), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n258), .B1(new_n848), .B2(KEYINPUT16), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n846), .B1(new_n849), .B2(new_n838), .ZN(new_n850));
  INV_X1    g0650(.A(new_n423), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n845), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n842), .A2(new_n414), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT37), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT105), .ZN(new_n855));
  XNOR2_X1  g0655(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n421), .A2(new_n841), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n427), .A2(new_n414), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT105), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n860), .B(KEYINPUT37), .C1(new_n852), .C2(new_n853), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n855), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n835), .B1(new_n844), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n855), .A2(new_n859), .A3(new_n861), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n864), .B(KEYINPUT38), .C1(new_n432), .C2(new_n842), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n601), .B(new_n368), .C1(new_n364), .C2(new_n659), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n370), .B(new_n658), .C1(new_n369), .C2(new_n376), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n870), .A2(new_n708), .A3(new_n706), .A4(new_n807), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n834), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n427), .A2(new_n858), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n856), .B1(new_n873), .B2(KEYINPUT108), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n427), .A2(new_n414), .A3(new_n858), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n873), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n877), .A2(KEYINPUT108), .A3(new_n414), .A4(new_n856), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n858), .B1(new_n607), .B2(new_n415), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n835), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n834), .B1(new_n881), .B2(new_n865), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n882), .A2(new_n709), .A3(new_n807), .A4(new_n870), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n872), .A2(G330), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n435), .A2(new_n710), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT110), .Z(new_n887));
  NAND4_X1  g0687(.A1(new_n872), .A2(new_n435), .A3(new_n709), .A4(new_n883), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT109), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n435), .A2(new_n724), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n614), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n890), .B(new_n892), .Z(new_n893));
  OAI211_X1 g0693(.A(new_n659), .B(new_n807), .C1(new_n638), .C2(new_n645), .ZN(new_n894));
  INV_X1    g0694(.A(new_n804), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n870), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT104), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n894), .A2(new_n895), .B1(new_n868), .B2(new_n869), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT104), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n898), .A2(new_n866), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n429), .A2(new_n424), .A3(new_n656), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT39), .B1(new_n881), .B2(new_n865), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n376), .A2(new_n370), .A3(new_n659), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT107), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n376), .A2(KEYINPUT107), .A3(new_n370), .A4(new_n659), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n905), .B(new_n910), .C1(new_n866), .C2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n902), .A2(new_n903), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n893), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n263), .B2(new_n652), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n480), .A2(new_n481), .ZN(new_n916));
  OAI211_X1 g0716(.A(G20), .B(new_n293), .C1(new_n916), .C2(KEYINPUT35), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n207), .B(new_n917), .C1(KEYINPUT35), .C2(new_n916), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT36), .Z(new_n919));
  OAI21_X1  g0719(.A(G77), .B1(new_n382), .B2(new_n212), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n920), .A2(new_n218), .B1(G50), .B2(new_n212), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n651), .A3(new_n650), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n915), .A2(new_n919), .A3(new_n922), .ZN(G367));
  OAI21_X1  g0723(.A(new_n642), .B1(new_n640), .B2(new_n659), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n635), .A2(new_n658), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n677), .A2(new_n927), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n668), .A2(KEYINPUT42), .A3(new_n926), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n565), .A2(new_n567), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n615), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(KEYINPUT111), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(KEYINPUT111), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n659), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT42), .B1(new_n668), .B2(new_n926), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n929), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n625), .A2(new_n626), .A3(new_n659), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n631), .A2(new_n633), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n633), .B2(new_n937), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n928), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n936), .A2(new_n928), .A3(new_n940), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n943), .B1(new_n942), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n683), .B(KEYINPUT41), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n670), .A2(new_n926), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT44), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT44), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n670), .A2(new_n952), .A3(new_n926), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n668), .A2(new_n669), .A3(new_n927), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT45), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n677), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n955), .B(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n677), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n959), .A2(new_n960), .A3(new_n951), .A4(new_n953), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n676), .B(KEYINPUT112), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n676), .A2(KEYINPUT112), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n666), .A2(new_n667), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n668), .ZN(new_n965));
  MUX2_X1   g0765(.A(new_n962), .B(new_n963), .S(new_n965), .Z(new_n966));
  NAND4_X1  g0766(.A1(new_n957), .A2(new_n961), .A3(new_n725), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n949), .B1(new_n967), .B2(new_n725), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n728), .B(KEYINPUT113), .Z(new_n969));
  OAI21_X1  g0769(.A(new_n947), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n818), .A2(G77), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n212), .B2(new_n749), .C1(new_n249), .C2(new_n769), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n771), .A2(new_n202), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n755), .A2(G58), .B1(new_n741), .B2(G137), .ZN(new_n974));
  INV_X1    g0774(.A(G159), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n974), .B1(new_n813), .B2(new_n756), .C1(new_n975), .C2(new_n746), .ZN(new_n976));
  NOR4_X1   g0776(.A1(new_n972), .A2(new_n274), .A3(new_n973), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n741), .A2(G317), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n755), .A2(G116), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT46), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n283), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n980), .B2(new_n979), .C1(new_n313), .C2(new_n749), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G311), .A2(new_n757), .B1(new_n772), .B2(G283), .ZN(new_n983));
  INV_X1    g0783(.A(G303), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(new_n762), .B2(new_n459), .C1(new_n984), .C2(new_n769), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n982), .B(new_n985), .C1(G294), .C2(new_n747), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n977), .B1(new_n978), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT47), .Z(new_n988));
  AOI21_X1  g0788(.A(new_n731), .B1(new_n988), .B2(new_n737), .ZN(new_n989));
  INV_X1    g0789(.A(new_n321), .ZN(new_n990));
  INV_X1    g0790(.A(new_n787), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n796), .B1(new_n223), .B2(new_n990), .C1(new_n235), .C2(new_n991), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n989), .B(new_n992), .C1(new_n798), .C2(new_n939), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n970), .A2(KEYINPUT114), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT114), .B1(new_n970), .B2(new_n993), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(G387));
  OR2_X1    g0797(.A1(new_n966), .A2(new_n725), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n966), .A2(new_n725), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(new_n683), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(G311), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n756), .A2(new_n782), .B1(new_n746), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT117), .Z(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n984), .B2(new_n771), .C1(new_n776), .C2(new_n769), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT48), .ZN(new_n1005));
  INV_X1    g0805(.A(G294), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1005), .B1(new_n783), .B2(new_n749), .C1(new_n1006), .C2(new_n754), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT49), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n741), .A2(G326), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n283), .B1(new_n818), .B2(G116), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G68), .A2(new_n772), .B1(new_n741), .B2(G150), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n323), .B2(new_n754), .C1(new_n975), .C2(new_n756), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n274), .B(new_n1015), .C1(new_n245), .C2(new_n747), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G50), .A2(new_n825), .B1(new_n818), .B2(G97), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n990), .C2(new_n749), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n736), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n666), .A2(new_n798), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n681), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1021), .A2(new_n791), .B1(G107), .B2(new_n223), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT115), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n409), .A2(G50), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(G45), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(G68), .A2(G77), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1021), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n991), .B1(new_n230), .B2(G45), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1023), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1031), .A2(new_n737), .A3(new_n795), .ZN(new_n1032));
  NOR4_X1   g0832(.A1(new_n1019), .A2(new_n1020), .A3(new_n731), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n966), .B2(new_n969), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1000), .A2(new_n1034), .ZN(G393));
  NAND2_X1  g0835(.A1(new_n957), .A2(new_n961), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n687), .B1(new_n1036), .B2(new_n999), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1037), .A2(new_n967), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n796), .B1(new_n459), .B2(new_n223), .C1(new_n243), .C2(new_n991), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n769), .A2(new_n975), .B1(new_n249), .B2(new_n756), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT51), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n749), .A2(new_n323), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n747), .A2(G50), .B1(new_n741), .B2(G143), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n212), .B2(new_n754), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(new_n245), .C2(new_n772), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n283), .A3(new_n1045), .A4(new_n824), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n769), .A2(new_n1001), .B1(new_n776), .B2(new_n756), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT52), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n746), .A2(new_n984), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n274), .B1(new_n749), .B2(new_n207), .C1(new_n1006), .C2(new_n771), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n818), .C2(G107), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n754), .A2(new_n783), .B1(new_n740), .B2(new_n782), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT118), .Z(new_n1053));
  NAND3_X1  g0853(.A1(new_n1048), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1046), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n731), .B1(new_n1055), .B2(new_n737), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1039), .B(new_n1056), .C1(new_n927), .C2(new_n798), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n969), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1057), .B1(new_n1036), .B2(new_n1058), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1038), .A2(new_n1059), .ZN(G390));
  AND3_X1   g0860(.A1(new_n863), .A2(KEYINPUT39), .A3(new_n865), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1061), .A2(new_n904), .B1(new_n899), .B2(new_n910), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n334), .B1(new_n1063), .B2(new_n305), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n336), .A2(new_n805), .B1(new_n319), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n658), .B(new_n1065), .C1(new_n715), .C2(new_n719), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n870), .B1(new_n1066), .B2(new_n804), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT119), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n910), .B1(new_n881), .B2(new_n865), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1068), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1062), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT120), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n706), .A2(G330), .A3(new_n708), .A4(new_n807), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n868), .A2(new_n869), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1062), .B(KEYINPUT120), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1074), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1072), .A2(new_n1073), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n896), .B1(new_n1083), .B2(new_n1077), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1066), .A2(new_n804), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1080), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n614), .A2(new_n891), .A3(new_n885), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1082), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1079), .A2(new_n1089), .A3(new_n1081), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n683), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1082), .A2(new_n969), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n793), .B1(new_n1061), .B2(new_n904), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n731), .B1(new_n830), .B2(new_n409), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT121), .Z(new_n1097));
  AOI22_X1  g0897(.A1(new_n757), .A2(G283), .B1(new_n741), .B2(G294), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n459), .B2(new_n771), .C1(new_n313), .C2(new_n746), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G87), .B2(new_n755), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G116), .A2(new_n825), .B1(new_n818), .B2(G68), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1042), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n274), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n755), .A2(G150), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT53), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G159), .B2(new_n750), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n274), .B1(new_n757), .B2(G128), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n740), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n818), .B2(G50), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n747), .A2(G137), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT122), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n825), .A2(G132), .B1(new_n772), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1106), .A2(new_n1110), .A3(new_n1111), .A4(new_n1114), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1103), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1095), .B(new_n1097), .C1(new_n736), .C2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1093), .A2(new_n1094), .A3(new_n1117), .ZN(G378));
  INV_X1    g0918(.A(KEYINPUT57), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n614), .A2(new_n891), .A3(new_n885), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n872), .A2(G330), .A3(new_n883), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n913), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n308), .B(KEYINPUT55), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n269), .A2(new_n841), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT56), .Z(new_n1126));
  XNOR2_X1  g0926(.A(new_n1124), .B(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n884), .A2(new_n903), .A3(new_n912), .A4(new_n902), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1123), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1127), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1119), .B1(new_n1121), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1127), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1123), .A2(new_n1128), .A3(new_n1127), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1089), .B1(new_n1081), .B2(new_n1079), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1137), .B(KEYINPUT57), .C1(new_n1120), .C2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1132), .A2(new_n1139), .A3(new_n683), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n969), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n830), .A2(new_n202), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n285), .B(new_n274), .C1(new_n754), .C2(new_n323), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n747), .A2(G97), .B1(new_n772), .B2(new_n321), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n207), .B2(new_n756), .C1(new_n783), .C2(new_n740), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(G68), .C2(new_n750), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n382), .B2(new_n762), .C1(new_n313), .C2(new_n769), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT58), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n202), .B1(new_n272), .B2(G41), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n825), .A2(G128), .B1(new_n755), .B2(new_n1113), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n756), .A2(new_n1108), .B1(new_n771), .B2(new_n812), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G150), .B2(new_n750), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(new_n816), .C2(new_n746), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT59), .Z(new_n1154));
  AOI21_X1  g0954(.A(G41), .B1(new_n818), .B2(G159), .ZN(new_n1155));
  AOI21_X1  g0955(.A(G33), .B1(new_n741), .B2(G124), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1148), .A2(new_n1149), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n731), .B1(new_n1158), .B2(new_n737), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1142), .B(new_n1159), .C1(new_n1134), .C2(new_n794), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1141), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1140), .A2(new_n1162), .ZN(G375));
  INV_X1    g0963(.A(KEYINPUT123), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n1058), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n283), .B1(new_n749), .B2(new_n202), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n755), .A2(G159), .B1(new_n772), .B2(G150), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n816), .B2(new_n756), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(G128), .C2(new_n741), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1113), .A2(new_n747), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G137), .A2(new_n825), .B1(new_n818), .B2(G58), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n769), .A2(new_n783), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n755), .A2(G97), .B1(new_n741), .B2(G303), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n207), .B2(new_n746), .C1(new_n1006), .C2(new_n756), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n321), .B2(new_n750), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n283), .B1(new_n772), .B2(G107), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n971), .A3(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1173), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1180), .A2(new_n737), .B1(new_n212), .B2(new_n830), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n730), .B(new_n1181), .C1(new_n870), .C2(new_n794), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1088), .A2(KEYINPUT123), .A3(new_n969), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1166), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT124), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1120), .A2(new_n1165), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n948), .A3(new_n1089), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT125), .Z(G381));
  XNOR2_X1  g0989(.A(G375), .B(KEYINPUT127), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT126), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(G378), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1093), .A2(KEYINPUT126), .A3(new_n1094), .A4(new_n1117), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1190), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n994), .A2(new_n995), .A3(G390), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OR4_X1    g0996(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1196), .A2(new_n1197), .ZN(G407));
  NAND2_X1  g0998(.A1(new_n1194), .A2(new_n657), .ZN(new_n1199));
  OAI211_X1 g0999(.A(G213), .B(new_n1199), .C1(new_n1196), .C2(new_n1197), .ZN(G409));
  NOR2_X1   g1000(.A1(G393), .A2(G396), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n802), .B1(new_n1000), .B2(new_n1034), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n970), .A2(new_n993), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1203), .B1(G390), .B2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1038), .A2(new_n1059), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n993), .B2(new_n970), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n995), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n970), .A2(KEYINPUT114), .A3(new_n993), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n1206), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1207), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1203), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1208), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n657), .A2(G213), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1140), .A2(G378), .A3(new_n1162), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1121), .A2(new_n1131), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1161), .B1(new_n1218), .B2(new_n948), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1216), .B1(new_n1217), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT60), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1186), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1120), .A2(new_n1165), .A3(KEYINPUT60), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1223), .A2(new_n683), .A3(new_n1089), .A4(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1185), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G384), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1185), .A2(G384), .A3(new_n1225), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n657), .A2(G213), .A3(G2897), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1221), .A2(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1235), .B(new_n1216), .C1(new_n1217), .C2(new_n1220), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT62), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(KEYINPUT62), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT61), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1215), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1214), .B1(new_n1195), .B2(new_n1207), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1208), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT61), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1236), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(KEYINPUT63), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT63), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1221), .B2(new_n1233), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1244), .B(new_n1246), .C1(new_n1245), .C2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1241), .A2(new_n1249), .ZN(G405));
  NAND2_X1  g1050(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(G375), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1140), .A2(G378), .A3(new_n1162), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(new_n1235), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1235), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1215), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1215), .B1(new_n1256), .B2(new_n1255), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(G402));
endmodule


