//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  XOR2_X1   g000(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n187), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G143), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(KEYINPUT64), .A3(G146), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n195), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT0), .A2(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n197), .A2(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n194), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n200), .A2(new_n201), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT65), .A2(G134), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT65), .A2(G134), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G137), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT11), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n211), .B1(new_n209), .B2(new_n210), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n208), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g033(.A1(KEYINPUT65), .A2(G134), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT65), .A2(G134), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G137), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n214), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n217), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT65), .B(G134), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT11), .B1(new_n225), .B2(new_n211), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n224), .A2(new_n226), .A3(G131), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n207), .B1(new_n219), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n229));
  INV_X1    g043(.A(G116), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G119), .ZN(new_n231));
  INV_X1    g045(.A(G119), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G116), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(G116), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(G119), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT67), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n237), .ZN(new_n240));
  OR2_X1    g054(.A1(new_n240), .A2(new_n235), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(G137), .B1(new_n220), .B2(new_n221), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  OAI22_X1  g059(.A1(new_n244), .A2(new_n245), .B1(G134), .B2(new_n211), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n225), .A2(new_n245), .A3(new_n211), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(G131), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n215), .A2(new_n208), .A3(new_n218), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  OAI21_X1  g065(.A(G128), .B1(new_n195), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n206), .ZN(new_n253));
  INV_X1    g067(.A(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(KEYINPUT1), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n194), .A2(KEYINPUT64), .A3(G146), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT64), .B1(new_n194), .B2(G146), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n204), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n249), .A2(new_n250), .A3(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n228), .A2(new_n243), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n243), .B1(new_n228), .B2(new_n260), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT28), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n228), .A2(new_n243), .A3(new_n260), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n193), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n228), .A2(new_n268), .A3(new_n260), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n228), .B2(new_n260), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n242), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n193), .A3(new_n264), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n216), .A2(KEYINPUT66), .B1(new_n213), .B2(G137), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n208), .B1(new_n275), .B2(new_n247), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n253), .A2(new_n258), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n227), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n207), .ZN(new_n279));
  OAI21_X1  g093(.A(G131), .B1(new_n224), .B2(new_n226), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n250), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT30), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n228), .A2(new_n268), .A3(new_n260), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n261), .B1(new_n284), .B2(new_n242), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT31), .A3(new_n193), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n267), .B1(new_n274), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT69), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n267), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT31), .B1(new_n285), .B2(new_n193), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n243), .B1(new_n282), .B2(new_n283), .ZN(new_n293));
  INV_X1    g107(.A(new_n193), .ZN(new_n294));
  NOR4_X1   g108(.A1(new_n293), .A2(new_n273), .A3(new_n294), .A4(new_n261), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n291), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n288), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n290), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n294), .B1(new_n293), .B2(new_n261), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n263), .A2(new_n193), .A3(new_n266), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n263), .A2(KEYINPUT72), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n307), .B(KEYINPUT28), .C1(new_n261), .C2(new_n262), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n266), .B(KEYINPUT73), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n309), .A2(KEYINPUT29), .A3(new_n193), .A4(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n305), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n314));
  OAI21_X1  g128(.A(G472), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n296), .A2(KEYINPUT32), .A3(new_n288), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n300), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT74), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n300), .A2(new_n315), .A3(new_n319), .A4(new_n316), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT25), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT23), .B1(new_n254), .B2(G119), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT75), .B1(new_n254), .B2(G119), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G110), .ZN(new_n326));
  XOR2_X1   g140(.A(G119), .B(G128), .Z(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT24), .B(G110), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n329), .A2(KEYINPUT16), .A3(G140), .ZN(new_n330));
  XNOR2_X1  g144(.A(G125), .B(G140), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n332), .A2(G146), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(G146), .ZN(new_n334));
  OAI221_X1 g148(.A(new_n326), .B1(new_n327), .B2(new_n328), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n327), .A2(new_n328), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n325), .B2(G110), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n331), .A2(new_n197), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n332), .B2(G146), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n337), .A2(KEYINPUT76), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT76), .B1(new_n337), .B2(new_n339), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n335), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G137), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n343), .B(new_n344), .Z(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n335), .B(new_n345), .C1(new_n340), .C2(new_n341), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n322), .B1(new_n349), .B2(G902), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n347), .A2(KEYINPUT25), .A3(new_n312), .A4(new_n348), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G217), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(G234), .B2(new_n312), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(G902), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n355), .B1(new_n349), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G478), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(KEYINPUT15), .ZN(new_n361));
  XOR2_X1   g175(.A(G128), .B(G143), .Z(new_n362));
  INV_X1    g176(.A(KEYINPUT13), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n254), .A2(G143), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n213), .B1(new_n365), .B2(new_n363), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT98), .B(G122), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(new_n230), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n230), .A2(G122), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT99), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT99), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n373), .B(new_n370), .C1(new_n368), .C2(new_n230), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n372), .A2(G107), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(G107), .B1(new_n372), .B2(new_n374), .ZN(new_n376));
  OAI221_X1 g190(.A(new_n367), .B1(new_n225), .B2(new_n362), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n362), .B(new_n225), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n370), .B(KEYINPUT14), .ZN(new_n379));
  OAI21_X1  g193(.A(G107), .B1(new_n379), .B2(new_n369), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(KEYINPUT100), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT100), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n376), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n377), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT9), .B(G234), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n387), .A2(new_n353), .A3(G953), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n377), .B(new_n388), .C1(new_n383), .C2(new_n385), .ZN(new_n391));
  AOI21_X1  g205(.A(G902), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT101), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI211_X1 g208(.A(KEYINPUT101), .B(G902), .C1(new_n390), .C2(new_n391), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n361), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI22_X1  g210(.A1(new_n392), .A2(new_n393), .B1(KEYINPUT15), .B2(new_n360), .ZN(new_n397));
  INV_X1    g211(.A(G952), .ZN(new_n398));
  AOI211_X1 g212(.A(G953), .B(new_n398), .C1(G234), .C2(G237), .ZN(new_n399));
  AOI211_X1 g213(.A(new_n312), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT21), .B(G898), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n396), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G214), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n405), .A2(G237), .A3(G953), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT93), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT93), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n194), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT94), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(G143), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT94), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n408), .A2(new_n410), .A3(new_n414), .A4(new_n194), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT17), .A3(G131), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n333), .A2(new_n334), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT97), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(G131), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT17), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n412), .A2(new_n208), .A3(new_n413), .A4(new_n415), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n417), .A2(KEYINPUT97), .A3(new_n418), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G113), .B(G122), .ZN(new_n428));
  INV_X1    g242(.A(G104), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n416), .A2(KEYINPUT95), .ZN(new_n431));
  NAND2_X1  g245(.A1(KEYINPUT18), .A2(G131), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(KEYINPUT18), .B(G131), .C1(new_n416), .C2(KEYINPUT95), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n331), .B(new_n197), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n427), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n430), .B1(new_n427), .B2(new_n436), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n312), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G475), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n422), .A2(new_n424), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n331), .B(KEYINPUT19), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n333), .B1(new_n197), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n436), .A2(new_n445), .A3(KEYINPUT96), .ZN(new_n446));
  INV_X1    g260(.A(new_n430), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT96), .B1(new_n436), .B2(new_n445), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n437), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n451));
  NOR2_X1   g265(.A1(G475), .A2(G902), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n450), .B2(new_n452), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n441), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n404), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G221), .ZN(new_n457));
  INV_X1    g271(.A(new_n387), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(new_n312), .ZN(new_n459));
  INV_X1    g273(.A(G469), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(new_n312), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n462));
  INV_X1    g276(.A(G107), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(KEYINPUT78), .A3(G104), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n429), .A2(G107), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT78), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n429), .B2(G107), .ZN(new_n468));
  OAI211_X1 g282(.A(G101), .B(new_n464), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT3), .B1(new_n429), .B2(G107), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n463), .A3(G104), .ZN(new_n472));
  INV_X1    g286(.A(G101), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n470), .A2(new_n472), .A3(new_n473), .A4(new_n465), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n259), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n258), .A2(KEYINPUT79), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n254), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n200), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT80), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n198), .A2(new_n199), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT79), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n204), .A4(new_n255), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n474), .A3(new_n469), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n482), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n486), .A2(new_n474), .A3(new_n469), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n258), .B(KEYINPUT79), .C1(new_n200), .C2(new_n480), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT80), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n462), .B(new_n478), .C1(new_n488), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n250), .A2(new_n280), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n483), .B1(new_n482), .B2(new_n487), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(KEYINPUT80), .A3(new_n490), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n477), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT81), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n497), .A2(KEYINPUT82), .A3(KEYINPUT12), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n492), .B(new_n493), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n476), .A2(new_n259), .A3(KEYINPUT10), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n470), .A2(new_n472), .A3(new_n465), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G101), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(KEYINPUT4), .A3(new_n474), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n504), .A3(G101), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n207), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n494), .A2(new_n495), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT10), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n493), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n493), .A2(KEYINPUT81), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT12), .B1(new_n496), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n499), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n189), .A2(G227), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT77), .ZN(new_n517));
  XNOR2_X1  g331(.A(G110), .B(G140), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n493), .A2(KEYINPUT83), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n510), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n510), .A2(new_n522), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n519), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n461), .B1(new_n526), .B2(G469), .ZN(new_n527));
  INV_X1    g341(.A(new_n524), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n510), .A2(new_n522), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n520), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n492), .A2(new_n493), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n496), .A2(new_n498), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT84), .B(new_n514), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n520), .B1(new_n510), .B2(new_n511), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT84), .B1(new_n499), .B2(new_n514), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n460), .A3(new_n312), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n459), .B1(new_n527), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n456), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G214), .B1(G237), .B2(G902), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT85), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n207), .A2(new_n329), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n277), .A2(KEYINPUT89), .A3(new_n329), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n253), .A2(new_n258), .A3(new_n329), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT89), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G224), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(G953), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n545), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n545), .B2(new_n550), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT6), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n241), .A2(new_n474), .A3(new_n469), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n234), .A2(new_n238), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT5), .ZN(new_n561));
  OAI21_X1  g375(.A(G113), .B1(new_n236), .B2(KEYINPUT5), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n559), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n242), .A2(new_n503), .A3(new_n505), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT86), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT86), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n242), .A2(new_n503), .A3(new_n567), .A4(new_n505), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n564), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(G110), .B(G122), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n558), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n568), .ZN(new_n572));
  INV_X1    g386(.A(new_n564), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n570), .B1(new_n574), .B2(KEYINPUT87), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT87), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n571), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n570), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n569), .B2(new_n576), .ZN(new_n580));
  AOI211_X1 g394(.A(KEYINPUT87), .B(new_n564), .C1(new_n566), .C2(new_n568), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n580), .A2(new_n558), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n557), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G210), .B1(G237), .B2(G902), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n572), .A2(new_n573), .A3(new_n570), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT7), .B1(new_n553), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n586), .B2(new_n553), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n545), .A2(new_n550), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n570), .B(KEYINPUT8), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n561), .A2(new_n563), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n476), .B1(new_n591), .B2(new_n241), .ZN(new_n592));
  INV_X1    g406(.A(new_n240), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT90), .B1(new_n593), .B2(KEYINPUT5), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(new_n562), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(KEYINPUT90), .A3(KEYINPUT5), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n559), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n590), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n585), .A2(new_n589), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n550), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n546), .A2(KEYINPUT91), .A3(new_n549), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n545), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n553), .A2(KEYINPUT7), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n599), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n583), .A2(new_n584), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n584), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n585), .A2(KEYINPUT6), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n580), .B2(new_n581), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n574), .A2(KEYINPUT87), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n611), .A2(KEYINPUT6), .A3(new_n577), .A4(new_n579), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n556), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n605), .A2(new_n585), .A3(new_n598), .A4(new_n589), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n312), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n608), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n542), .B1(new_n607), .B2(new_n616), .ZN(new_n617));
  AND4_X1   g431(.A1(new_n321), .A2(new_n359), .A3(new_n540), .A4(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n473), .ZN(G3));
  AND2_X1   g433(.A1(new_n539), .A2(new_n359), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n290), .A2(new_n298), .ZN(new_n621));
  OAI21_X1  g435(.A(G472), .B1(new_n287), .B2(G902), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n622), .A2(KEYINPUT102), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(KEYINPUT102), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n617), .A2(new_n403), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n620), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n392), .A2(new_n360), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n360), .A2(new_n312), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n390), .A2(new_n391), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n632), .B1(G478), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n455), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n628), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n454), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(KEYINPUT103), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n453), .A2(new_n645), .B1(G475), .B2(new_n440), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n396), .A2(new_n397), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n628), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  INV_X1    g466(.A(new_n342), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n346), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT104), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n356), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n355), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n540), .A2(new_n617), .A3(new_n625), .A4(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  INV_X1    g476(.A(new_n539), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n318), .B2(new_n320), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n400), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n399), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n644), .A2(new_n646), .A3(new_n647), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n617), .A2(new_n659), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  XNOR2_X1  g487(.A(new_n668), .B(KEYINPUT39), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n539), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT40), .Z(new_n676));
  INV_X1    g490(.A(new_n659), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n285), .A2(new_n294), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n261), .A2(new_n262), .A3(new_n193), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(G902), .ZN(new_n680));
  OAI21_X1  g494(.A(G472), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n300), .A2(new_n316), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n607), .A2(new_n616), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT38), .ZN(new_n684));
  INV_X1    g498(.A(new_n542), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n455), .A2(new_n684), .A3(new_n647), .A4(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n676), .A2(new_n677), .A3(new_n682), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT105), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  NAND3_X1  g503(.A1(new_n455), .A2(new_n636), .A3(new_n668), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n670), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n664), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  AOI21_X1  g507(.A(new_n358), .B1(new_n318), .B2(new_n320), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n537), .A2(new_n312), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  INV_X1    g510(.A(new_n459), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n697), .A3(new_n538), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n626), .A3(new_n637), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NOR3_X1   g516(.A1(new_n648), .A2(new_n698), .A3(new_n626), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n694), .A2(KEYINPUT106), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT106), .B1(new_n694), .B2(new_n703), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NAND4_X1  g521(.A1(new_n617), .A2(new_n696), .A3(new_n697), .A4(new_n538), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n537), .A2(new_n460), .A3(new_n312), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n460), .B1(new_n537), .B2(new_n312), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(KEYINPUT107), .A3(new_n697), .A4(new_n617), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n321), .A2(new_n715), .A3(new_n456), .A4(new_n659), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  INV_X1    g531(.A(new_n455), .ZN(new_n718));
  INV_X1    g532(.A(new_n647), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n683), .A2(new_n685), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n711), .A2(new_n712), .A3(new_n459), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n292), .A2(new_n295), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n193), .B1(new_n309), .B2(new_n310), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n288), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n622), .A2(new_n725), .A3(new_n359), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n721), .A2(new_n403), .A3(new_n722), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  NAND3_X1  g542(.A1(new_n622), .A2(new_n725), .A3(new_n659), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n622), .A2(new_n725), .A3(new_n659), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n690), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT107), .B1(new_n722), .B2(new_n617), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n698), .A2(new_n709), .A3(new_n720), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n715), .A2(KEYINPUT109), .A3(new_n733), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT110), .B(G125), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G27));
  INV_X1    g556(.A(new_n683), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n459), .A2(new_n542), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n525), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n523), .A2(KEYINPUT111), .A3(new_n524), .A4(new_n519), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n521), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n460), .B1(new_n749), .B2(new_n312), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n711), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n690), .A2(new_n745), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT32), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n287), .B2(new_n289), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n316), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT112), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n316), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n315), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n359), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT42), .B1(new_n753), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n745), .A2(new_n751), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n690), .A2(KEYINPUT42), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n694), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n208), .ZN(G33));
  INV_X1    g581(.A(new_n669), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n321), .A2(new_n768), .A3(new_n359), .A4(new_n763), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  NAND2_X1  g584(.A1(new_n635), .A2(G478), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n629), .A3(new_n631), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n772), .A2(new_n455), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT114), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n636), .B(KEYINPUT113), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n773), .B1(new_n776), .B2(new_n455), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n625), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n659), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n779), .A4(new_n659), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n743), .A2(new_n685), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT115), .ZN(new_n787));
  OAI21_X1  g601(.A(G469), .B1(new_n526), .B2(KEYINPUT45), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n749), .A2(new_n789), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n788), .A2(new_n790), .B1(new_n460), .B2(new_n312), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n538), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n697), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n674), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n782), .A2(new_n799), .A3(new_n783), .A4(new_n785), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n787), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n796), .B(new_n803), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n321), .A2(new_n359), .A3(new_n690), .A4(new_n784), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT116), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n804), .A2(new_n808), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NAND3_X1  g625(.A1(new_n359), .A2(new_n636), .A3(new_n744), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n684), .A2(new_n455), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n682), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n713), .B(KEYINPUT49), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n667), .B1(new_n775), .B2(new_n777), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n784), .A2(new_n698), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n730), .A2(new_n732), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT122), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n817), .A2(new_n726), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(KEYINPUT121), .A3(new_n785), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n823), .B2(new_n784), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n711), .A2(new_n712), .A3(new_n697), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n825), .B(new_n827), .C1(new_n804), .C2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n684), .A2(new_n685), .A3(new_n698), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n824), .A2(KEYINPUT50), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT50), .ZN(new_n832));
  INV_X1    g646(.A(new_n830), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n823), .B2(new_n833), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n359), .A2(new_n814), .A3(new_n818), .A4(new_n399), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n718), .A2(new_n772), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n831), .A2(new_n834), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n822), .A2(new_n829), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  INV_X1    g656(.A(new_n761), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n819), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT48), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n835), .A2(new_n638), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(G952), .A3(new_n189), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n824), .B2(new_n715), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n841), .A2(new_n842), .A3(new_n845), .A4(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n637), .B1(new_n719), .B2(new_n455), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n620), .A2(new_n625), .A3(new_n850), .A4(new_n627), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n660), .A2(new_n851), .A3(new_n727), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n618), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n700), .A2(new_n716), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n853), .B(new_n854), .C1(new_n705), .C2(new_n704), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n644), .A2(new_n646), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n719), .A2(new_n659), .A3(new_n668), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n857), .A3(new_n784), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n664), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n752), .A2(new_n820), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n769), .A3(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(new_n766), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n321), .B(new_n539), .C1(new_n671), .C2(new_n691), .ZN(new_n864));
  INV_X1    g678(.A(new_n668), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n751), .A2(new_n459), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n721), .A3(new_n677), .A4(new_n682), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n715), .A2(KEYINPUT109), .A3(new_n733), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT109), .B1(new_n715), .B2(new_n733), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n864), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n740), .A2(KEYINPUT117), .A3(new_n864), .A4(new_n867), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n872), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n863), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  XOR2_X1   g695(.A(KEYINPUT118), .B(KEYINPUT52), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n872), .A2(new_n873), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n867), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n738), .B2(new_n739), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(KEYINPUT52), .A3(new_n864), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(KEYINPUT53), .A3(new_n863), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n879), .A2(new_n880), .A3(new_n881), .A4(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n861), .A2(new_n766), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(new_n706), .A3(new_n853), .A4(new_n854), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT117), .B1(new_n885), .B2(new_n864), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n870), .A2(new_n871), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT52), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n888), .B(new_n881), .C1(new_n896), .C2(KEYINPUT53), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT119), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n887), .A2(new_n863), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n878), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n863), .B(KEYINPUT53), .C1(new_n875), .C2(new_n876), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n881), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n889), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT120), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(new_n889), .C1(new_n898), .C2(new_n902), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n849), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(G952), .A2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n816), .B1(new_n907), .B2(new_n908), .ZN(G75));
  NAND2_X1  g723(.A1(new_n398), .A2(G953), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT123), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n312), .B1(new_n879), .B2(new_n888), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(G210), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n578), .A2(new_n582), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n556), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n583), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT55), .Z(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n911), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n915), .B2(new_n920), .ZN(G51));
  INV_X1    g736(.A(new_n911), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n461), .B(KEYINPUT57), .ZN(new_n924));
  INV_X1    g738(.A(new_n897), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n881), .B1(new_n879), .B2(new_n888), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n537), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n788), .A2(new_n790), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n912), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n923), .B1(new_n928), .B2(new_n930), .ZN(G54));
  NAND3_X1  g745(.A1(new_n912), .A2(KEYINPUT58), .A3(G475), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(new_n450), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n450), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n923), .B1(new_n933), .B2(new_n934), .ZN(G60));
  XNOR2_X1  g749(.A(new_n630), .B(KEYINPUT59), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n635), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n925), .B2(new_n926), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n911), .ZN(new_n939));
  INV_X1    g753(.A(new_n936), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n904), .A2(new_n906), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(new_n941), .B2(new_n635), .ZN(G63));
  NAND2_X1  g756(.A1(new_n879), .A2(new_n888), .ZN(new_n943));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT60), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n349), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n656), .A2(new_n657), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n947), .B(new_n911), .C1(new_n948), .C2(new_n946), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G66));
  OAI21_X1  g765(.A(G953), .B1(new_n401), .B2(new_n551), .ZN(new_n952));
  INV_X1    g766(.A(new_n855), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n916), .B1(G898), .B2(new_n189), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT124), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G69));
  AOI21_X1  g771(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n958));
  INV_X1    g772(.A(new_n766), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n798), .A2(new_n721), .A3(new_n843), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n810), .A2(new_n959), .A3(new_n769), .A4(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n740), .A2(new_n864), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n801), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n801), .A2(KEYINPUT127), .A3(new_n962), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n961), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n284), .B(new_n443), .Z(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n189), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n688), .A2(new_n962), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT62), .Z(new_n972));
  XOR2_X1   g786(.A(new_n850), .B(KEYINPUT125), .Z(new_n973));
  NOR2_X1   g787(.A1(new_n675), .A2(new_n784), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n694), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT126), .Z(new_n976));
  AND3_X1   g790(.A1(new_n801), .A2(new_n810), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(G953), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  OAI22_X1  g792(.A1(new_n967), .A2(new_n970), .B1(new_n978), .B2(new_n969), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n958), .B1(new_n979), .B2(new_n665), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n958), .B2(new_n979), .ZN(G72));
  NAND2_X1  g795(.A1(new_n967), .A2(new_n953), .ZN(new_n982));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n293), .A2(new_n193), .A3(new_n261), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n900), .A2(new_n901), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n301), .A2(new_n272), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n972), .A2(new_n977), .A3(new_n953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n984), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n923), .B1(new_n992), .B2(new_n678), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n987), .A2(new_n990), .A3(new_n993), .ZN(G57));
endmodule


