//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969;
  NOR2_X1   g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT90), .B(G36gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G29gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(KEYINPUT15), .A3(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n210), .A2(new_n204), .A3(new_n211), .A4(new_n206), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n209), .A2(KEYINPUT17), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT17), .B1(new_n209), .B2(new_n212), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(G1gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G1gat), .B2(new_n216), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(G8gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n215), .A2(KEYINPUT91), .A3(new_n221), .ZN(new_n222));
  NOR3_X1   g021(.A1(new_n213), .A2(new_n220), .A3(new_n214), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n209), .A2(new_n212), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT91), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n222), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT18), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n220), .B(new_n224), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n229), .B(KEYINPUT92), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT13), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n228), .A2(KEYINPUT18), .A3(new_n229), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n232), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT11), .B(G169gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(G197gat), .ZN(new_n241));
  XOR2_X1   g040(.A(G113gat), .B(G141gat), .Z(new_n242));
  XOR2_X1   g041(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g042(.A(new_n243), .B(KEYINPUT12), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n232), .A2(new_n244), .A3(new_n237), .A4(new_n238), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(KEYINPUT93), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT93), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(new_n246), .B2(new_n247), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT95), .ZN(new_n254));
  XNOR2_X1  g053(.A(G127gat), .B(G155gat), .ZN(new_n255));
  INV_X1    g054(.A(G211gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G71gat), .B(G78gat), .Z(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT9), .ZN(new_n260));
  INV_X1    g059(.A(G71gat), .ZN(new_n261));
  INV_X1    g060(.A(G78gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G57gat), .B(G64gat), .Z(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n263), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n258), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT94), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT21), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n221), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G183gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n273), .A3(new_n221), .ZN(new_n274));
  NAND2_X1  g073(.A1(G231gat), .A2(G233gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n276), .B1(new_n272), .B2(new_n274), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n257), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n279), .ZN(new_n281));
  INV_X1    g080(.A(new_n257), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n277), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n268), .A2(KEYINPUT21), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n280), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n286), .B1(new_n280), .B2(new_n283), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G85gat), .A2(G92gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT7), .ZN(new_n291));
  NAND2_X1  g090(.A1(G99gat), .A2(G106gat), .ZN(new_n292));
  INV_X1    g091(.A(G85gat), .ZN(new_n293));
  INV_X1    g092(.A(G92gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(KEYINPUT8), .A2(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G99gat), .B(G106gat), .Z(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n215), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n297), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n296), .B(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(G232gat), .A2(G233gat), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n301), .A2(new_n224), .B1(KEYINPUT41), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(G134gat), .B(G162gat), .Z(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n302), .A2(KEYINPUT41), .ZN(new_n307));
  XNOR2_X1  g106(.A(G190gat), .B(G218gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n306), .B(new_n309), .Z(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n254), .B1(new_n289), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(KEYINPUT95), .B(new_n310), .C1(new_n287), .C2(new_n288), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n269), .A2(KEYINPUT10), .A3(new_n301), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT98), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT96), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n298), .A2(new_n268), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n267), .A3(new_n265), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(KEYINPUT97), .B(KEYINPUT10), .Z(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n322), .ZN(new_n324));
  AOI211_X1 g123(.A(KEYINPUT98), .B(new_n324), .C1(new_n318), .C2(new_n320), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n314), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT99), .ZN(new_n327));
  NAND2_X1  g126(.A1(G230gat), .A2(G233gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n327), .B1(new_n326), .B2(new_n328), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n321), .A2(new_n328), .ZN(new_n333));
  XNOR2_X1  g132(.A(G120gat), .B(G148gat), .ZN(new_n334));
  INV_X1    g133(.A(G176gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G204gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n332), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n326), .A2(new_n328), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n338), .B1(new_n342), .B2(new_n333), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n312), .A2(new_n313), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G190gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n273), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT24), .A3(new_n349), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n349), .A2(KEYINPUT24), .ZN(new_n351));
  NAND2_X1  g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT65), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT25), .B1(new_n352), .B2(new_n353), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n358));
  INV_X1    g157(.A(G169gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n335), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n356), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n357), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n363), .A2(new_n350), .A3(new_n351), .A4(new_n352), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n347), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT66), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n373));
  NOR2_X1   g172(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT26), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(new_n359), .A3(new_n335), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n352), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n373), .A2(new_n374), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n370), .A2(new_n371), .A3(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n376), .A2(new_n349), .A3(new_n380), .A4(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT29), .B1(new_n367), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n385), .B(KEYINPUT72), .Z(new_n386));
  OAI21_X1  g185(.A(KEYINPUT73), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n388));
  INV_X1    g187(.A(new_n386), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n355), .A2(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n370), .A2(new_n371), .A3(new_n381), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n381), .B1(new_n370), .B2(new_n371), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n380), .A2(new_n349), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n388), .B(new_n389), .C1(new_n395), .C2(KEYINPUT29), .ZN(new_n396));
  XNOR2_X1  g195(.A(G211gat), .B(G218gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT22), .ZN(new_n398));
  INV_X1    g197(.A(G218gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(new_n256), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G197gat), .B(G204gat), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(new_n401), .A3(new_n400), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT74), .B1(new_n390), .B2(new_n394), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT74), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n367), .A2(new_n408), .A3(new_n383), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n409), .A3(new_n386), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n387), .A2(new_n396), .A3(new_n406), .A4(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n407), .A2(new_n409), .A3(new_n412), .A4(new_n389), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n386), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n405), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G8gat), .B(G36gat), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(G64gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(new_n294), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n411), .A2(new_n415), .A3(new_n419), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(KEYINPUT30), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(new_n424), .A3(new_n420), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT0), .B(G57gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(G85gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G127gat), .B(G134gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT68), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(G134gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n437));
  INV_X1    g236(.A(G120gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G113gat), .ZN(new_n439));
  INV_X1    g238(.A(G113gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G120gat), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n435), .B(new_n437), .C1(KEYINPUT1), .C2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT1), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT69), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n441), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT69), .B1(new_n438), .B2(G113gat), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n444), .B(new_n433), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G141gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G148gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT77), .ZN(new_n452));
  INV_X1    g251(.A(G148gat), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(G141gat), .B2(new_n453), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n450), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G155gat), .A2(G162gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n459), .B2(KEYINPUT2), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n453), .A2(G141gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n450), .A2(G148gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT76), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n457), .A2(KEYINPUT2), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n453), .A2(G141gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT76), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT75), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n459), .A2(new_n469), .A3(new_n457), .ZN(new_n470));
  INV_X1    g269(.A(new_n457), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT75), .B1(new_n471), .B2(new_n458), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AOI221_X4 g272(.A(KEYINPUT78), .B1(new_n456), .B2(new_n460), .C1(new_n468), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT78), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n468), .A2(new_n473), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n456), .A2(new_n460), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n449), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n451), .A2(new_n465), .A3(new_n466), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n466), .B1(new_n451), .B2(new_n465), .ZN(new_n481));
  INV_X1    g280(.A(new_n464), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n470), .A2(new_n472), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n477), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(new_n449), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n479), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G225gat), .A2(G233gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n489), .B(KEYINPUT79), .Z(new_n490));
  AOI21_X1  g289(.A(KEYINPUT83), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n492));
  INV_X1    g291(.A(new_n490), .ZN(new_n493));
  AOI211_X1 g292(.A(new_n492), .B(new_n493), .C1(new_n479), .C2(new_n487), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT5), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n449), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT4), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n468), .A2(new_n473), .B1(new_n456), .B2(new_n460), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT81), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT81), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n501), .A3(new_n497), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n485), .A2(KEYINPUT80), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT80), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n449), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n500), .B(new_n502), .C1(new_n506), .C2(new_n497), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT82), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT3), .B1(new_n474), .B2(new_n478), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT3), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n496), .B1(new_n510), .B2(new_n498), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n490), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n507), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n508), .B1(new_n507), .B2(new_n512), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n495), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n511), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n516), .B(new_n517), .C1(KEYINPUT4), .C2(new_n506), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n518), .A2(KEYINPUT5), .A3(new_n490), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n432), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT6), .ZN(new_n521));
  INV_X1    g320(.A(new_n519), .ZN(new_n522));
  INV_X1    g321(.A(new_n514), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n512), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n431), .B(new_n522), .C1(new_n525), .C2(new_n495), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  OAI211_X1 g326(.A(KEYINPUT6), .B(new_n432), .C1(new_n515), .C2(new_n519), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n427), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n496), .A2(new_n367), .A3(new_n383), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n449), .B1(new_n390), .B2(new_n394), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT34), .ZN(new_n532));
  NAND2_X1  g331(.A1(G227gat), .A2(G233gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT64), .Z(new_n534));
  NAND4_X1  g333(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT71), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n539));
  XOR2_X1   g338(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n530), .A2(new_n531), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT32), .B1(new_n543), .B2(new_n534), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n535), .B(KEYINPUT71), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n547), .A2(new_n544), .A3(new_n541), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G43gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(G71gat), .B(G99gat), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n550), .B(new_n551), .Z(new_n552));
  NOR2_X1   g351(.A1(new_n543), .A2(new_n534), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(KEYINPUT33), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n548), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G22gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n405), .A2(new_n412), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n510), .B1(new_n560), .B2(KEYINPUT84), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT84), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n405), .B2(new_n412), .ZN(new_n563));
  OAI22_X1  g362(.A1(new_n561), .A2(new_n563), .B1(new_n478), .B2(new_n474), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT85), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT29), .B1(new_n498), .B2(new_n510), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(KEYINPUT86), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(KEYINPUT86), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n406), .A3(new_n569), .ZN(new_n570));
  OAI221_X1 g369(.A(KEYINPUT85), .B1(new_n474), .B2(new_n478), .C1(new_n561), .C2(new_n563), .ZN(new_n571));
  INV_X1    g370(.A(G228gat), .ZN(new_n572));
  INV_X1    g371(.A(G233gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n566), .A2(new_n570), .A3(new_n571), .A4(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n504), .B1(new_n476), .B2(new_n477), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n476), .A2(new_n504), .A3(new_n477), .ZN(new_n577));
  AOI211_X1 g376(.A(new_n576), .B(new_n577), .C1(new_n510), .C2(new_n560), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n567), .A2(new_n405), .ZN(new_n579));
  OAI22_X1  g378(.A1(new_n578), .A2(new_n579), .B1(new_n572), .B2(new_n573), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n559), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n559), .A3(new_n580), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT87), .ZN(new_n583));
  XOR2_X1   g382(.A(G78gat), .B(G106gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT31), .ZN(new_n585));
  INV_X1    g384(.A(G50gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT88), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n582), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n581), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n581), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n582), .A2(new_n591), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n594), .B(new_n589), .C1(new_n595), .C2(new_n588), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n558), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n529), .A2(new_n597), .A3(KEYINPUT35), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT35), .B1(new_n529), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n593), .A2(new_n596), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n529), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n558), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n420), .B1(new_n416), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n413), .A2(new_n414), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n406), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n387), .A2(new_n396), .A3(new_n410), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n609), .B(KEYINPUT37), .C1(new_n610), .C2(new_n406), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n421), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n411), .A2(KEYINPUT37), .A3(new_n415), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n607), .B1(new_n606), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n527), .A2(new_n528), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT89), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n496), .B1(new_n577), .B2(new_n576), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n497), .A2(new_n619), .B1(new_n509), .B2(new_n511), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n493), .B1(new_n620), .B2(new_n517), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n432), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n518), .A2(new_n490), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n488), .A2(new_n490), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(KEYINPUT39), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n627), .A3(KEYINPUT40), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n513), .A2(new_n514), .ZN(new_n629));
  INV_X1    g428(.A(new_n495), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n519), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n628), .B1(new_n631), .B2(new_n431), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n621), .A2(new_n622), .A3(new_n625), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n518), .A2(new_n622), .A3(new_n490), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n431), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n633), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(new_n425), .A3(new_n423), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n618), .B1(new_n632), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT40), .B1(new_n623), .B2(new_n627), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n426), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n641), .A2(KEYINPUT89), .A3(new_n520), .A4(new_n628), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n617), .A2(new_n639), .A3(new_n601), .A4(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n602), .A2(new_n604), .A3(new_n643), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n253), .B(new_n346), .C1(new_n600), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n527), .A2(new_n528), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n427), .ZN(new_n650));
  AND2_X1   g449(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(G8gat), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n657), .A2(KEYINPUT100), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(KEYINPUT100), .ZN(new_n659));
  OAI22_X1  g458(.A1(new_n655), .A2(new_n656), .B1(new_n658), .B2(new_n659), .ZN(G1325gat));
  INV_X1    g459(.A(new_n558), .ZN(new_n661));
  AOI21_X1  g460(.A(G15gat), .B1(new_n645), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n604), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n663), .A2(G15gat), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n645), .B2(new_n664), .ZN(G1326gat));
  INV_X1    g464(.A(new_n601), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n645), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n670));
  AND4_X1   g469(.A1(new_n601), .A2(new_n617), .A3(new_n639), .A4(new_n642), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n604), .B1(new_n529), .B2(new_n601), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n602), .A2(new_n643), .A3(KEYINPUT101), .A4(new_n604), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n600), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n311), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n600), .A2(new_n644), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(KEYINPUT44), .A3(new_n311), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n289), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n344), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n248), .ZN(new_n685));
  OAI21_X1  g484(.A(G29gat), .B1(new_n685), .B2(new_n646), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n682), .A2(new_n344), .A3(new_n310), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n679), .A2(new_n252), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(G29gat), .A3(new_n646), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT45), .Z(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n691), .ZN(G1328gat));
  OAI21_X1  g491(.A(new_n205), .B1(new_n685), .B2(new_n426), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n689), .A2(new_n426), .A3(new_n205), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT46), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1329gat));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n663), .A3(new_n248), .A4(new_n683), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G43gat), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(G43gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n688), .A2(new_n702), .A3(new_n661), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT102), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n698), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1330gat));
  NAND4_X1  g506(.A1(new_n684), .A2(G50gat), .A3(new_n666), .A4(new_n248), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n586), .B1(new_n689), .B2(new_n601), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n708), .A2(KEYINPUT48), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT48), .B1(new_n708), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(G1331gat));
  INV_X1    g511(.A(new_n248), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n675), .A2(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n312), .A2(new_n313), .A3(new_n344), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n647), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g518(.A1(new_n716), .A2(new_n426), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  AND2_X1   g520(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n720), .B2(new_n721), .ZN(G1333gat));
  OAI21_X1  g523(.A(G71gat), .B1(new_n716), .B2(new_n604), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n714), .A2(new_n661), .A3(new_n715), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n726), .B1(new_n731), .B2(new_n261), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g532(.A1(new_n716), .A2(new_n601), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(new_n262), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n682), .A2(new_n248), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n344), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT105), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n681), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n646), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n740), .A2(KEYINPUT106), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(KEYINPUT106), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(G85gat), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n675), .A2(new_n311), .A3(new_n736), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n675), .A2(KEYINPUT51), .A3(new_n311), .A4(new_n736), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n748), .A2(new_n293), .A3(new_n647), .A4(new_n344), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n743), .A2(new_n749), .ZN(G1336gat));
  NAND3_X1  g549(.A1(new_n681), .A2(new_n427), .A3(new_n738), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n345), .A2(G92gat), .A3(new_n426), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT52), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n746), .A2(new_n747), .B1(new_n756), .B2(new_n753), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n751), .A2(G92gat), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(G1337gat));
  OAI21_X1  g560(.A(G99gat), .B1(new_n739), .B2(new_n604), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n345), .A2(G99gat), .A3(new_n558), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT108), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(G1338gat));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769));
  INV_X1    g568(.A(G106gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n666), .A2(new_n344), .A3(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT109), .Z(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n769), .B1(new_n748), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g573(.A(KEYINPUT110), .B(new_n772), .C1(new_n746), .C2(new_n747), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n678), .A2(new_n738), .A3(new_n666), .A4(new_n680), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n768), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n771), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n748), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n768), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n767), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n778), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n785), .A2(new_n774), .A3(new_n775), .ZN(new_n786));
  OAI211_X1 g585(.A(KEYINPUT111), .B(new_n782), .C1(new_n786), .C2(new_n768), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1339gat));
  INV_X1    g587(.A(new_n228), .ZN(new_n789));
  INV_X1    g588(.A(new_n229), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n789), .A2(new_n790), .B1(new_n234), .B2(new_n236), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n791), .A2(new_n243), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n247), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n340), .B2(new_n343), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n326), .A2(new_n328), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT54), .B(new_n797), .C1(new_n330), .C2(new_n331), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n338), .B1(new_n341), .B2(KEYINPUT54), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(KEYINPUT55), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n798), .B2(new_n800), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n248), .B(new_n340), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n795), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n310), .ZN(new_n807));
  INV_X1    g606(.A(new_n331), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n796), .B1(new_n808), .B2(new_n329), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n799), .B1(new_n809), .B2(KEYINPUT54), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n803), .ZN(new_n811));
  INV_X1    g610(.A(new_n804), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n339), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n793), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n311), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n682), .B1(new_n807), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n346), .A2(new_n248), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n647), .B(new_n597), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n597), .ZN(new_n821));
  INV_X1    g620(.A(new_n815), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n311), .B1(new_n795), .B2(new_n805), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n289), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n346), .A2(new_n248), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(KEYINPUT112), .A3(new_n647), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n820), .A2(new_n426), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n440), .A3(new_n248), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n818), .A2(new_n427), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831), .B2(new_n253), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(G1340gat));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n438), .A3(new_n344), .ZN(new_n834));
  OAI21_X1  g633(.A(G120gat), .B1(new_n831), .B2(new_n345), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1341gat));
  NAND3_X1  g635(.A1(new_n830), .A2(G127gat), .A3(new_n682), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT113), .ZN(new_n838));
  AOI21_X1  g637(.A(G127gat), .B1(new_n828), .B2(new_n682), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(G1342gat));
  NOR2_X1   g639(.A1(new_n310), .A2(new_n427), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT114), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n820), .A2(new_n827), .A3(new_n436), .A4(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n826), .A2(new_n647), .A3(new_n841), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n844), .A2(new_n845), .B1(G134gat), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT115), .B1(new_n844), .B2(new_n845), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n843), .A2(new_n849), .A3(KEYINPUT56), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT116), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1343gat));
  NAND2_X1  g654(.A1(new_n807), .A2(new_n815), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n817), .B1(new_n856), .B2(new_n289), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n604), .A2(new_n647), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n857), .A2(new_n601), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n426), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n450), .A3(new_n252), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n858), .A2(new_n427), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n864), .B(new_n666), .C1(new_n816), .C2(new_n817), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT55), .B1(new_n801), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT117), .B(new_n803), .C1(new_n798), .C2(new_n800), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n252), .B(new_n340), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n311), .B1(new_n869), .B2(new_n795), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n289), .B1(new_n870), .B2(new_n822), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n601), .B1(new_n871), .B2(new_n825), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n863), .B(new_n865), .C1(new_n872), .C2(new_n864), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n253), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n861), .A2(new_n862), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n861), .A2(KEYINPUT119), .A3(new_n862), .A4(new_n874), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n803), .B1(new_n810), .B2(KEYINPUT117), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n801), .A2(new_n866), .A3(KEYINPUT55), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n339), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n794), .B1(new_n881), .B2(new_n252), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n815), .B1(new_n882), .B2(new_n311), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n817), .B1(new_n883), .B2(new_n289), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT57), .B1(new_n884), .B2(new_n601), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n885), .A2(new_n248), .A3(new_n863), .A4(new_n865), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G141gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT118), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n886), .A2(new_n889), .A3(G141gat), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n888), .A2(new_n861), .A3(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n877), .B(new_n878), .C1(new_n891), .C2(new_n862), .ZN(G1344gat));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  INV_X1    g693(.A(new_n871), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n346), .A2(new_n252), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n864), .B(new_n666), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT57), .B1(new_n857), .B2(new_n601), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n863), .B(KEYINPUT121), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n897), .A2(new_n898), .A3(new_n344), .A4(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n894), .B1(new_n900), .B2(G148gat), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n453), .A2(KEYINPUT59), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n873), .B2(new_n345), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT120), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n885), .A2(new_n344), .A3(new_n863), .A4(new_n865), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n906), .A3(new_n902), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n901), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n860), .A2(new_n453), .A3(new_n344), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n893), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n900), .A2(G148gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT59), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n905), .A2(new_n906), .A3(new_n902), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n906), .B1(new_n905), .B2(new_n902), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(KEYINPUT122), .A3(new_n909), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n911), .A2(new_n917), .ZN(G1345gat));
  AOI21_X1  g717(.A(G155gat), .B1(new_n860), .B2(new_n682), .ZN(new_n919));
  INV_X1    g718(.A(new_n873), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n682), .A2(G155gat), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT123), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n873), .B2(new_n310), .ZN(new_n924));
  INV_X1    g723(.A(G162gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n859), .A2(new_n925), .A3(new_n842), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n647), .A2(new_n426), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n826), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n248), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n929), .A2(G169gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n252), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT124), .ZN(G1348gat));
  NAND2_X1  g732(.A1(new_n929), .A2(new_n344), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g734(.A1(new_n929), .A2(new_n682), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G183gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n368), .A2(new_n369), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n936), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g739(.A1(new_n929), .A2(new_n311), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n941), .A2(new_n942), .A3(new_n347), .ZN(new_n943));
  XOR2_X1   g742(.A(KEYINPUT61), .B(G190gat), .Z(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n941), .B2(new_n944), .ZN(G1351gat));
  XNOR2_X1  g744(.A(KEYINPUT125), .B(G197gat), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n604), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT126), .Z(new_n948));
  NAND3_X1  g747(.A1(new_n897), .A2(new_n898), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n949), .B2(new_n253), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n857), .A2(new_n601), .A3(new_n947), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n713), .A2(new_n946), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n953), .ZN(G1352gat));
  NAND3_X1  g753(.A1(new_n951), .A2(new_n337), .A3(new_n344), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT62), .Z(new_n956));
  NAND2_X1  g755(.A1(new_n897), .A2(new_n898), .ZN(new_n957));
  INV_X1    g756(.A(new_n948), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n957), .A2(new_n345), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n337), .B2(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n951), .A2(new_n256), .A3(new_n682), .ZN(new_n961));
  OR3_X1    g760(.A1(new_n957), .A2(new_n289), .A3(new_n947), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n951), .B2(new_n311), .ZN(new_n966));
  INV_X1    g765(.A(new_n949), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n310), .A2(new_n399), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT127), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n966), .B1(new_n967), .B2(new_n969), .ZN(G1355gat));
endmodule


