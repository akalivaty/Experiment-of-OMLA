

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750;

  BUF_X1 U374 ( .A(n529), .Z(n353) );
  XNOR2_X1 U375 ( .A(n520), .B(KEYINPUT105), .ZN(n749) );
  OR2_X1 U376 ( .A1(n354), .A2(n580), .ZN(n582) );
  NOR2_X1 U377 ( .A1(n538), .A2(n523), .ZN(n524) );
  XNOR2_X1 U378 ( .A(n395), .B(KEYINPUT39), .ZN(n399) );
  BUF_X1 U379 ( .A(n602), .Z(n354) );
  AND2_X1 U380 ( .A1(n545), .A2(n407), .ZN(n516) );
  AND2_X1 U381 ( .A1(n572), .A2(n394), .ZN(n393) );
  BUF_X1 U382 ( .A(n673), .Z(n355) );
  XNOR2_X1 U383 ( .A(n463), .B(n462), .ZN(n673) );
  NOR2_X1 U384 ( .A1(n401), .A2(G902), .ZN(n463) );
  XNOR2_X1 U385 ( .A(n356), .B(n357), .ZN(n455) );
  XNOR2_X1 U386 ( .A(n489), .B(n441), .ZN(n400) );
  XNOR2_X1 U387 ( .A(KEYINPUT77), .B(G110), .ZN(n421) );
  XNOR2_X1 U388 ( .A(n449), .B(n409), .ZN(n356) );
  XOR2_X2 U389 ( .A(G104), .B(G107), .Z(n422) );
  INV_X2 U390 ( .A(KEYINPUT69), .ZN(n364) );
  XNOR2_X1 U391 ( .A(G143), .B(G104), .ZN(n485) );
  AND2_X1 U392 ( .A1(n541), .A2(n540), .ZN(n658) );
  XNOR2_X2 U393 ( .A(n542), .B(KEYINPUT101), .ZN(n690) );
  XNOR2_X2 U394 ( .A(n364), .B(G131), .ZN(n489) );
  OR2_X1 U395 ( .A1(n538), .A2(n519), .ZN(n520) );
  NOR2_X1 U396 ( .A1(n661), .A2(n648), .ZN(n550) );
  INV_X4 U397 ( .A(G953), .ZN(n451) );
  XNOR2_X1 U398 ( .A(n619), .B(KEYINPUT87), .ZN(n620) );
  NOR2_X1 U399 ( .A1(n645), .A2(n552), .ZN(n553) );
  AND2_X1 U400 ( .A1(n358), .A2(n748), .ZN(n376) );
  XNOR2_X1 U401 ( .A(n516), .B(n515), .ZN(n538) );
  NOR2_X1 U402 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U403 ( .A1(n690), .A2(KEYINPUT47), .ZN(n387) );
  INV_X1 U404 ( .A(n571), .ZN(n394) );
  NAND2_X1 U405 ( .A1(n411), .A2(n439), .ZN(n440) );
  XOR2_X1 U406 ( .A(G113), .B(G122), .Z(n488) );
  XNOR2_X2 U407 ( .A(n621), .B(KEYINPUT79), .ZN(n672) );
  XNOR2_X2 U408 ( .A(n476), .B(n381), .ZN(n712) );
  NOR2_X1 U409 ( .A1(n570), .A2(n406), .ZN(n391) );
  XNOR2_X1 U410 ( .A(n602), .B(n573), .ZN(n406) );
  NOR2_X1 U411 ( .A1(G237), .A2(G953), .ZN(n470) );
  NOR2_X1 U412 ( .A1(n513), .A2(n539), .ZN(n514) );
  XNOR2_X1 U413 ( .A(n383), .B(n480), .ZN(n668) );
  XNOR2_X1 U414 ( .A(n375), .B(n579), .ZN(n374) );
  XNOR2_X1 U415 ( .A(n468), .B(G113), .ZN(n396) );
  XNOR2_X1 U416 ( .A(n397), .B(G119), .ZN(n467) );
  XNOR2_X1 U417 ( .A(G116), .B(KEYINPUT3), .ZN(n397) );
  XNOR2_X1 U418 ( .A(n389), .B(n388), .ZN(n494) );
  NAND2_X1 U419 ( .A1(n673), .A2(n674), .ZN(n679) );
  XNOR2_X1 U420 ( .A(n478), .B(G472), .ZN(n568) );
  XNOR2_X1 U421 ( .A(n562), .B(KEYINPUT1), .ZN(n517) );
  XOR2_X1 U422 ( .A(G116), .B(G107), .Z(n499) );
  XNOR2_X1 U423 ( .A(G134), .B(G122), .ZN(n497) );
  XOR2_X1 U424 ( .A(KEYINPUT98), .B(KEYINPUT9), .Z(n498) );
  NAND2_X1 U425 ( .A1(n371), .A2(n368), .ZN(n689) );
  NAND2_X1 U426 ( .A1(n369), .A2(n359), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n403), .B(n402), .ZN(n564) );
  XNOR2_X1 U428 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n402) );
  BUF_X1 U429 ( .A(n517), .Z(n680) );
  NOR2_X1 U430 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U431 ( .A(KEYINPUT11), .B(KEYINPUT96), .ZN(n483) );
  INV_X1 U432 ( .A(n484), .ZN(n388) );
  INV_X1 U433 ( .A(KEYINPUT106), .ZN(n385) );
  INV_X1 U434 ( .A(G902), .ZN(n477) );
  NAND2_X1 U435 ( .A1(n370), .A2(n373), .ZN(n369) );
  NOR2_X1 U436 ( .A1(n406), .A2(n693), .ZN(n370) );
  NOR2_X1 U437 ( .A1(n560), .A2(n561), .ZN(n585) );
  NAND2_X1 U438 ( .A1(n585), .A2(n677), .ZN(n403) );
  OR2_X1 U439 ( .A1(G237), .A2(G902), .ZN(n433) );
  XNOR2_X1 U440 ( .A(G902), .B(KEYINPUT15), .ZN(n611) );
  XNOR2_X1 U441 ( .A(n496), .B(n495), .ZN(n539) );
  XNOR2_X1 U442 ( .A(n467), .B(n396), .ZN(n474) );
  XOR2_X1 U443 ( .A(KEYINPUT74), .B(KEYINPUT16), .Z(n418) );
  XNOR2_X1 U444 ( .A(n647), .B(KEYINPUT100), .ZN(n604) );
  INV_X1 U445 ( .A(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U446 ( .A(n366), .B(n365), .ZN(n686) );
  INV_X1 U447 ( .A(KEYINPUT95), .ZN(n365) );
  NOR2_X1 U448 ( .A1(n363), .A2(n547), .ZN(n366) );
  BUF_X1 U449 ( .A(n568), .Z(n677) );
  OR2_X1 U450 ( .A1(n541), .A2(n540), .ZN(n647) );
  XNOR2_X1 U451 ( .A(n539), .B(n390), .ZN(n541) );
  INV_X1 U452 ( .A(KEYINPUT97), .ZN(n390) );
  NOR2_X1 U453 ( .A1(n679), .A2(n562), .ZN(n546) );
  XNOR2_X1 U454 ( .A(n506), .B(n505), .ZN(n716) );
  XNOR2_X1 U455 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U456 ( .A(n501), .B(n500), .Z(n506) );
  BUF_X1 U457 ( .A(n709), .Z(n720) );
  NOR2_X1 U458 ( .A1(n451), .A2(G952), .ZN(n725) );
  NOR2_X1 U459 ( .A1(n689), .A2(n576), .ZN(n578) );
  XNOR2_X1 U460 ( .A(n574), .B(KEYINPUT40), .ZN(n750) );
  NAND2_X1 U461 ( .A1(n592), .A2(n591), .ZN(n664) );
  INV_X1 U462 ( .A(n647), .ZN(n660) );
  XNOR2_X1 U463 ( .A(n514), .B(KEYINPUT103), .ZN(n575) );
  XOR2_X1 U464 ( .A(KEYINPUT92), .B(G110), .Z(n357) );
  AND2_X1 U465 ( .A1(n664), .A2(n593), .ZN(n358) );
  XOR2_X1 U466 ( .A(KEYINPUT112), .B(KEYINPUT41), .Z(n359) );
  NOR2_X1 U467 ( .A1(n575), .A2(n406), .ZN(n360) );
  OR2_X1 U468 ( .A1(n693), .A2(n359), .ZN(n361) );
  XOR2_X1 U469 ( .A(n635), .B(KEYINPUT60), .Z(n362) );
  OR2_X1 U470 ( .A1(n517), .A2(n679), .ZN(n363) );
  OR2_X2 U471 ( .A1(n517), .A2(n679), .ZN(n543) );
  NAND2_X1 U472 ( .A1(n750), .A2(n404), .ZN(n375) );
  NAND2_X1 U473 ( .A1(n391), .A2(n393), .ZN(n395) );
  NAND2_X1 U474 ( .A1(n376), .A2(n374), .ZN(n596) );
  XNOR2_X1 U475 ( .A(n543), .B(n385), .ZN(n384) );
  NAND2_X1 U476 ( .A1(n509), .A2(n414), .ZN(n512) );
  XNOR2_X1 U477 ( .A(n482), .B(n481), .ZN(n509) );
  NAND2_X1 U478 ( .A1(n545), .A2(n668), .ZN(n482) );
  XNOR2_X1 U479 ( .A(n557), .B(n556), .ZN(n616) );
  NAND2_X1 U480 ( .A1(n712), .A2(n477), .ZN(n380) );
  XNOR2_X1 U481 ( .A(n367), .B(n362), .ZN(G60) );
  NAND2_X1 U482 ( .A1(n634), .A2(n633), .ZN(n367) );
  NOR2_X1 U483 ( .A1(n530), .A2(n749), .ZN(n531) );
  XNOR2_X1 U484 ( .A(n434), .B(n410), .ZN(n565) );
  NAND2_X1 U485 ( .A1(n372), .A2(n373), .ZN(n371) );
  NOR2_X1 U486 ( .A1(n406), .A2(n361), .ZN(n372) );
  INV_X1 U487 ( .A(n575), .ZN(n373) );
  XNOR2_X1 U488 ( .A(n583), .B(KEYINPUT109), .ZN(n748) );
  NOR2_X1 U489 ( .A1(n377), .A2(n749), .ZN(n525) );
  INV_X1 U490 ( .A(n529), .ZN(n377) );
  XNOR2_X1 U491 ( .A(n353), .B(G119), .ZN(G21) );
  XNOR2_X2 U492 ( .A(n524), .B(n378), .ZN(n529) );
  INV_X1 U493 ( .A(KEYINPUT32), .ZN(n378) );
  XNOR2_X2 U494 ( .A(n379), .B(KEYINPUT0), .ZN(n545) );
  NOR2_X2 U495 ( .A1(n565), .A2(n440), .ZN(n379) );
  XNOR2_X2 U496 ( .A(n380), .B(n448), .ZN(n562) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n381) );
  XNOR2_X2 U498 ( .A(n740), .B(G146), .ZN(n476) );
  XNOR2_X2 U499 ( .A(n382), .B(KEYINPUT4), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n382), .B(n499), .ZN(n500) );
  XNOR2_X2 U501 ( .A(G143), .B(G128), .ZN(n382) );
  NAND2_X1 U502 ( .A1(n384), .A2(n535), .ZN(n383) );
  XNOR2_X2 U503 ( .A(n422), .B(n421), .ZN(n732) );
  XNOR2_X1 U504 ( .A(n417), .B(n415), .ZN(n405) );
  XNOR2_X1 U505 ( .A(n405), .B(n442), .ZN(n420) );
  NAND2_X1 U506 ( .A1(n386), .A2(n656), .ZN(n594) );
  XNOR2_X1 U507 ( .A(n387), .B(KEYINPUT76), .ZN(n386) );
  XNOR2_X1 U508 ( .A(n456), .B(KEYINPUT10), .ZN(n484) );
  XNOR2_X2 U509 ( .A(G146), .B(G125), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n487), .B(n483), .ZN(n389) );
  INV_X1 U511 ( .A(n658), .ZN(n584) );
  NAND2_X1 U512 ( .A1(n658), .A2(n585), .ZN(n586) );
  XNOR2_X1 U513 ( .A(n546), .B(KEYINPUT94), .ZN(n572) );
  NAND2_X1 U514 ( .A1(n392), .A2(n393), .ZN(n580) );
  INV_X1 U515 ( .A(n570), .ZN(n392) );
  NAND2_X1 U516 ( .A1(n399), .A2(n658), .ZN(n574) );
  AND2_X1 U517 ( .A1(n399), .A2(n398), .ZN(n666) );
  INV_X1 U518 ( .A(n604), .ZN(n398) );
  XNOR2_X2 U519 ( .A(n400), .B(n442), .ZN(n740) );
  XNOR2_X1 U520 ( .A(n401), .B(n721), .ZN(n722) );
  XNOR2_X1 U521 ( .A(n458), .B(n739), .ZN(n401) );
  XNOR2_X1 U522 ( .A(n404), .B(G137), .ZN(G39) );
  XNOR2_X1 U523 ( .A(n578), .B(n577), .ZN(n404) );
  NOR2_X1 U524 ( .A1(n690), .A2(n406), .ZN(n691) );
  BUF_X1 U525 ( .A(n617), .Z(n741) );
  NOR2_X2 U526 ( .A1(n616), .A2(n741), .ZN(n670) );
  XNOR2_X2 U527 ( .A(n544), .B(KEYINPUT31), .ZN(n661) );
  NOR2_X1 U528 ( .A1(n602), .A2(n693), .ZN(n434) );
  AND2_X1 U529 ( .A1(n373), .A2(n674), .ZN(n407) );
  XOR2_X1 U530 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n408) );
  XNOR2_X1 U531 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n409) );
  XNOR2_X1 U532 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n410) );
  AND2_X1 U533 ( .A1(n701), .A2(n438), .ZN(n411) );
  AND2_X1 U534 ( .A1(KEYINPUT44), .A2(KEYINPUT68), .ZN(n412) );
  XOR2_X1 U535 ( .A(n631), .B(n630), .Z(n413) );
  XOR2_X1 U536 ( .A(n581), .B(n508), .Z(n414) );
  INV_X1 U537 ( .A(n690), .ZN(n566) );
  INV_X1 U538 ( .A(G137), .ZN(n468) );
  XNOR2_X1 U539 ( .A(n492), .B(n491), .ZN(n493) );
  BUF_X1 U540 ( .A(n446), .Z(n426) );
  XNOR2_X1 U541 ( .A(n461), .B(KEYINPUT25), .ZN(n462) );
  XNOR2_X1 U542 ( .A(n455), .B(n454), .ZN(n458) );
  INV_X1 U543 ( .A(n725), .ZN(n633) );
  XNOR2_X1 U544 ( .A(n723), .B(n722), .ZN(n724) );
  XOR2_X1 U545 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n415) );
  NAND2_X1 U546 ( .A1(G224), .A2(n451), .ZN(n416) );
  XNOR2_X1 U547 ( .A(n416), .B(n456), .ZN(n417) );
  XNOR2_X1 U548 ( .A(n488), .B(n418), .ZN(n419) );
  XNOR2_X1 U549 ( .A(n419), .B(n467), .ZN(n731) );
  XNOR2_X1 U550 ( .A(n420), .B(n731), .ZN(n428) );
  INV_X1 U551 ( .A(n428), .ZN(n425) );
  XOR2_X2 U552 ( .A(KEYINPUT67), .B(G101), .Z(n469) );
  INV_X1 U553 ( .A(KEYINPUT72), .ZN(n423) );
  XNOR2_X1 U554 ( .A(n469), .B(n423), .ZN(n424) );
  XNOR2_X1 U555 ( .A(n732), .B(n424), .ZN(n446) );
  NAND2_X1 U556 ( .A1(n425), .A2(n426), .ZN(n430) );
  INV_X1 U557 ( .A(n426), .ZN(n427) );
  NAND2_X1 U558 ( .A1(n428), .A2(n427), .ZN(n429) );
  NAND2_X1 U559 ( .A1(n430), .A2(n429), .ZN(n624) );
  NAND2_X1 U560 ( .A1(n624), .A2(n611), .ZN(n432) );
  NAND2_X1 U561 ( .A1(G210), .A2(n433), .ZN(n431) );
  XNOR2_X2 U562 ( .A(n432), .B(n431), .ZN(n602) );
  NAND2_X1 U563 ( .A1(G214), .A2(n433), .ZN(n588) );
  INV_X1 U564 ( .A(n588), .ZN(n693) );
  NAND2_X1 U565 ( .A1(G234), .A2(G237), .ZN(n435) );
  XNOR2_X1 U566 ( .A(n435), .B(KEYINPUT14), .ZN(n701) );
  NOR2_X1 U567 ( .A1(G902), .A2(n451), .ZN(n437) );
  NOR2_X1 U568 ( .A1(G953), .A2(G952), .ZN(n436) );
  NOR2_X1 U569 ( .A1(n437), .A2(n436), .ZN(n438) );
  NAND2_X1 U570 ( .A1(G953), .A2(G898), .ZN(n439) );
  INV_X1 U571 ( .A(G134), .ZN(n441) );
  XOR2_X1 U572 ( .A(G137), .B(G140), .Z(n457) );
  NAND2_X1 U573 ( .A1(n451), .A2(G227), .ZN(n443) );
  XNOR2_X1 U574 ( .A(n443), .B(KEYINPUT81), .ZN(n444) );
  XNOR2_X1 U575 ( .A(n457), .B(n444), .ZN(n445) );
  XNOR2_X1 U576 ( .A(KEYINPUT71), .B(G469), .ZN(n447) );
  XNOR2_X1 U577 ( .A(n447), .B(KEYINPUT70), .ZN(n448) );
  XNOR2_X1 U578 ( .A(G128), .B(G119), .ZN(n449) );
  XOR2_X1 U579 ( .A(KEYINPUT86), .B(KEYINPUT8), .Z(n453) );
  NAND2_X1 U580 ( .A1(G234), .A2(n451), .ZN(n452) );
  XNOR2_X1 U581 ( .A(n453), .B(n452), .ZN(n502) );
  NAND2_X1 U582 ( .A1(n502), .A2(G221), .ZN(n454) );
  XNOR2_X1 U583 ( .A(n457), .B(n484), .ZN(n739) );
  XOR2_X1 U584 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n460) );
  NAND2_X1 U585 ( .A1(G234), .A2(n611), .ZN(n459) );
  XNOR2_X1 U586 ( .A(n460), .B(n459), .ZN(n464) );
  NAND2_X1 U587 ( .A1(G217), .A2(n464), .ZN(n461) );
  NAND2_X1 U588 ( .A1(n464), .A2(G221), .ZN(n466) );
  INV_X1 U589 ( .A(KEYINPUT21), .ZN(n465) );
  XNOR2_X1 U590 ( .A(n466), .B(n465), .ZN(n674) );
  XOR2_X1 U591 ( .A(n469), .B(KEYINPUT5), .Z(n472) );
  XNOR2_X1 U592 ( .A(n470), .B(KEYINPUT78), .ZN(n490) );
  NAND2_X1 U593 ( .A1(G210), .A2(n490), .ZN(n471) );
  XNOR2_X1 U594 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U595 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U596 ( .A(n476), .B(n475), .ZN(n639) );
  NAND2_X1 U597 ( .A1(n639), .A2(n477), .ZN(n478) );
  INV_X1 U598 ( .A(KEYINPUT6), .ZN(n479) );
  XNOR2_X1 U599 ( .A(n568), .B(n479), .ZN(n535) );
  INV_X1 U600 ( .A(n535), .ZN(n587) );
  XNOR2_X1 U601 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n480) );
  XNOR2_X1 U602 ( .A(KEYINPUT13), .B(G475), .ZN(n496) );
  XOR2_X1 U603 ( .A(KEYINPUT12), .B(G140), .Z(n486) );
  XNOR2_X1 U604 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U605 ( .A(n489), .B(n488), .ZN(n492) );
  NAND2_X1 U606 ( .A1(n490), .A2(G214), .ZN(n491) );
  XNOR2_X1 U607 ( .A(n494), .B(n493), .ZN(n629) );
  NOR2_X1 U608 ( .A1(G902), .A2(n629), .ZN(n495) );
  XNOR2_X1 U609 ( .A(n498), .B(n497), .ZN(n501) );
  NAND2_X1 U610 ( .A1(G217), .A2(n502), .ZN(n504) );
  XNOR2_X1 U611 ( .A(KEYINPUT7), .B(KEYINPUT99), .ZN(n503) );
  NOR2_X1 U612 ( .A1(G902), .A2(n716), .ZN(n507) );
  XNOR2_X1 U613 ( .A(G478), .B(n507), .ZN(n540) );
  INV_X1 U614 ( .A(n540), .ZN(n513) );
  NAND2_X1 U615 ( .A1(n539), .A2(n513), .ZN(n581) );
  INV_X1 U616 ( .A(KEYINPUT83), .ZN(n508) );
  INV_X1 U617 ( .A(KEYINPUT82), .ZN(n510) );
  XNOR2_X1 U618 ( .A(n510), .B(KEYINPUT35), .ZN(n511) );
  XNOR2_X2 U619 ( .A(n512), .B(n511), .ZN(n636) );
  XNOR2_X1 U620 ( .A(n636), .B(KEYINPUT68), .ZN(n526) );
  XNOR2_X1 U621 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n515) );
  NOR2_X1 U622 ( .A1(n355), .A2(n677), .ZN(n518) );
  NAND2_X1 U623 ( .A1(n680), .A2(n518), .ZN(n519) );
  INV_X1 U624 ( .A(n355), .ZN(n534) );
  NAND2_X1 U625 ( .A1(n587), .A2(n534), .ZN(n521) );
  NOR2_X1 U626 ( .A1(n521), .A2(n680), .ZN(n522) );
  XOR2_X1 U627 ( .A(KEYINPUT84), .B(n522), .Z(n523) );
  NAND2_X1 U628 ( .A1(n526), .A2(n525), .ZN(n528) );
  INV_X1 U629 ( .A(KEYINPUT44), .ZN(n527) );
  NAND2_X1 U630 ( .A1(n528), .A2(n527), .ZN(n533) );
  NAND2_X1 U631 ( .A1(n529), .A2(n412), .ZN(n530) );
  NAND2_X1 U632 ( .A1(n531), .A2(n636), .ZN(n532) );
  NAND2_X1 U633 ( .A1(n533), .A2(n532), .ZN(n555) );
  NOR2_X1 U634 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U635 ( .A1(n536), .A2(n680), .ZN(n537) );
  NOR2_X1 U636 ( .A1(n538), .A2(n537), .ZN(n645) );
  NAND2_X1 U637 ( .A1(n584), .A2(n604), .ZN(n542) );
  INV_X1 U638 ( .A(n677), .ZN(n547) );
  NAND2_X1 U639 ( .A1(n545), .A2(n686), .ZN(n544) );
  INV_X1 U640 ( .A(n545), .ZN(n549) );
  NAND2_X1 U641 ( .A1(n547), .A2(n572), .ZN(n548) );
  NOR2_X1 U642 ( .A1(n549), .A2(n548), .ZN(n648) );
  NOR2_X1 U643 ( .A1(n690), .A2(n550), .ZN(n551) );
  XNOR2_X1 U644 ( .A(n551), .B(KEYINPUT102), .ZN(n552) );
  XNOR2_X1 U645 ( .A(n553), .B(KEYINPUT104), .ZN(n554) );
  NAND2_X1 U646 ( .A1(n555), .A2(n554), .ZN(n557) );
  INV_X1 U647 ( .A(KEYINPUT45), .ZN(n556) );
  INV_X1 U648 ( .A(n674), .ZN(n561) );
  NAND2_X1 U649 ( .A1(G953), .A2(G900), .ZN(n558) );
  NAND2_X1 U650 ( .A1(n411), .A2(n558), .ZN(n559) );
  XOR2_X1 U651 ( .A(KEYINPUT85), .B(n559), .Z(n571) );
  OR2_X1 U652 ( .A1(n673), .A2(n571), .ZN(n560) );
  XOR2_X1 U653 ( .A(KEYINPUT110), .B(n562), .Z(n563) );
  NAND2_X1 U654 ( .A1(n564), .A2(n563), .ZN(n576) );
  NOR2_X1 U655 ( .A1(n565), .A2(n576), .ZN(n656) );
  NAND2_X1 U656 ( .A1(n566), .A2(n656), .ZN(n567) );
  NAND2_X1 U657 ( .A1(n567), .A2(KEYINPUT47), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n568), .A2(n588), .ZN(n569) );
  XNOR2_X1 U659 ( .A(KEYINPUT30), .B(n569), .ZN(n570) );
  INV_X1 U660 ( .A(KEYINPUT38), .ZN(n573) );
  XNOR2_X1 U661 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n577) );
  INV_X1 U662 ( .A(KEYINPUT46), .ZN(n579) );
  NOR2_X1 U663 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n598) );
  NOR2_X1 U665 ( .A1(n598), .A2(n354), .ZN(n590) );
  XNOR2_X1 U666 ( .A(KEYINPUT36), .B(n590), .ZN(n592) );
  INV_X1 U667 ( .A(n680), .ZN(n591) );
  XNOR2_X1 U668 ( .A(n594), .B(KEYINPUT75), .ZN(n595) );
  XNOR2_X1 U669 ( .A(n597), .B(KEYINPUT48), .ZN(n607) );
  XNOR2_X1 U670 ( .A(n598), .B(KEYINPUT107), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n599), .A2(n680), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n600), .B(KEYINPUT43), .ZN(n601) );
  XNOR2_X1 U673 ( .A(KEYINPUT108), .B(n601), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n603), .A2(n354), .ZN(n667) );
  INV_X1 U675 ( .A(n667), .ZN(n605) );
  NOR2_X1 U676 ( .A1(n605), .A2(n666), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n617) );
  INV_X1 U678 ( .A(KEYINPUT2), .ZN(n608) );
  NOR2_X1 U679 ( .A1(n608), .A2(KEYINPUT65), .ZN(n609) );
  NOR2_X1 U680 ( .A1(n670), .A2(n609), .ZN(n610) );
  NOR2_X1 U681 ( .A1(n610), .A2(n611), .ZN(n615) );
  INV_X1 U682 ( .A(n611), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n612), .A2(KEYINPUT2), .ZN(n613) );
  AND2_X1 U684 ( .A1(n613), .A2(KEYINPUT65), .ZN(n614) );
  NOR2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n622) );
  INV_X1 U686 ( .A(n616), .ZN(n726) );
  INV_X1 U687 ( .A(n617), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n618), .A2(KEYINPUT2), .ZN(n619) );
  NAND2_X1 U689 ( .A1(n726), .A2(n620), .ZN(n621) );
  NOR2_X2 U690 ( .A1(n622), .A2(n672), .ZN(n709) );
  NAND2_X1 U691 ( .A1(n709), .A2(G210), .ZN(n626) );
  XOR2_X1 U692 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n623) );
  XNOR2_X1 U693 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U694 ( .A(n626), .B(n625), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n627), .A2(n633), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n628), .B(n408), .ZN(G51) );
  NAND2_X1 U697 ( .A1(n709), .A2(G475), .ZN(n632) );
  XOR2_X1 U698 ( .A(KEYINPUT59), .B(KEYINPUT64), .Z(n631) );
  XNOR2_X1 U699 ( .A(n629), .B(KEYINPUT90), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n632), .B(n413), .ZN(n634) );
  XNOR2_X1 U701 ( .A(KEYINPUT66), .B(KEYINPUT122), .ZN(n635) );
  XNOR2_X1 U702 ( .A(G122), .B(KEYINPUT127), .ZN(n637) );
  XOR2_X1 U703 ( .A(n637), .B(n636), .Z(G24) );
  NAND2_X1 U704 ( .A1(n709), .A2(G472), .ZN(n641) );
  XNOR2_X1 U705 ( .A(KEYINPUT89), .B(KEYINPUT62), .ZN(n638) );
  XNOR2_X1 U706 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U707 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X2 U708 ( .A1(n642), .A2(n725), .ZN(n644) );
  XNOR2_X1 U709 ( .A(KEYINPUT91), .B(KEYINPUT63), .ZN(n643) );
  XNOR2_X1 U710 ( .A(n644), .B(n643), .ZN(G57) );
  XOR2_X1 U711 ( .A(G101), .B(n645), .Z(G3) );
  NAND2_X1 U712 ( .A1(n648), .A2(n658), .ZN(n646) );
  XNOR2_X1 U713 ( .A(n646), .B(G104), .ZN(G6) );
  XOR2_X1 U714 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n650) );
  NAND2_X1 U715 ( .A1(n648), .A2(n660), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U717 ( .A(G107), .B(n651), .ZN(G9) );
  XOR2_X1 U718 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n653) );
  NAND2_X1 U719 ( .A1(n656), .A2(n660), .ZN(n652) );
  XNOR2_X1 U720 ( .A(n653), .B(n652), .ZN(n655) );
  XOR2_X1 U721 ( .A(G128), .B(KEYINPUT114), .Z(n654) );
  XNOR2_X1 U722 ( .A(n655), .B(n654), .ZN(G30) );
  NAND2_X1 U723 ( .A1(n656), .A2(n658), .ZN(n657) );
  XNOR2_X1 U724 ( .A(n657), .B(G146), .ZN(G48) );
  NAND2_X1 U725 ( .A1(n661), .A2(n658), .ZN(n659) );
  XNOR2_X1 U726 ( .A(n659), .B(G113), .ZN(G15) );
  NAND2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U728 ( .A(n662), .B(G116), .ZN(G18) );
  XOR2_X1 U729 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n663) );
  XNOR2_X1 U730 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U731 ( .A(G125), .B(n665), .ZN(G27) );
  XOR2_X1 U732 ( .A(G134), .B(n666), .Z(G36) );
  XNOR2_X1 U733 ( .A(G140), .B(n667), .ZN(G42) );
  INV_X1 U734 ( .A(n668), .ZN(n695) );
  NOR2_X1 U735 ( .A1(n689), .A2(n695), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n669), .A2(G953), .ZN(n707) );
  NOR2_X1 U737 ( .A1(n670), .A2(KEYINPUT2), .ZN(n671) );
  NOR2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n705) );
  NOR2_X1 U739 ( .A1(n674), .A2(n355), .ZN(n675) );
  XOR2_X1 U740 ( .A(KEYINPUT49), .B(n675), .Z(n676) );
  NOR2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U742 ( .A(KEYINPUT117), .B(n678), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U744 ( .A(KEYINPUT50), .B(n681), .Z(n682) );
  NOR2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U746 ( .A(n684), .B(KEYINPUT118), .ZN(n685) );
  NOR2_X1 U747 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U748 ( .A(KEYINPUT51), .B(n687), .Z(n688) );
  NOR2_X1 U749 ( .A1(n689), .A2(n688), .ZN(n698) );
  NOR2_X1 U750 ( .A1(n373), .A2(n691), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U752 ( .A1(n360), .A2(n694), .ZN(n696) );
  NOR2_X1 U753 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U754 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U755 ( .A(n699), .B(KEYINPUT119), .Z(n700) );
  XNOR2_X1 U756 ( .A(KEYINPUT52), .B(n700), .ZN(n703) );
  NAND2_X1 U757 ( .A1(n701), .A2(G952), .ZN(n702) );
  NOR2_X1 U758 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U759 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U760 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U761 ( .A(KEYINPUT53), .B(n708), .Z(G75) );
  NAND2_X1 U762 ( .A1(n720), .A2(G469), .ZN(n714) );
  XNOR2_X1 U763 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n710) );
  XOR2_X1 U764 ( .A(n710), .B(KEYINPUT57), .Z(n711) );
  XNOR2_X1 U765 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U766 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U767 ( .A1(n725), .A2(n715), .ZN(G54) );
  NAND2_X1 U768 ( .A1(n720), .A2(G478), .ZN(n718) );
  XOR2_X1 U769 ( .A(n716), .B(KEYINPUT123), .Z(n717) );
  XNOR2_X1 U770 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n725), .A2(n719), .ZN(G63) );
  NAND2_X1 U772 ( .A1(n720), .A2(G217), .ZN(n723) );
  XOR2_X1 U773 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n721) );
  NOR2_X1 U774 ( .A1(n725), .A2(n724), .ZN(G66) );
  NAND2_X1 U775 ( .A1(n726), .A2(n451), .ZN(n730) );
  NAND2_X1 U776 ( .A1(G953), .A2(G224), .ZN(n727) );
  XNOR2_X1 U777 ( .A(KEYINPUT61), .B(n727), .ZN(n728) );
  NAND2_X1 U778 ( .A1(n728), .A2(G898), .ZN(n729) );
  NAND2_X1 U779 ( .A1(n730), .A2(n729), .ZN(n738) );
  XNOR2_X1 U780 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U781 ( .A(n733), .B(KEYINPUT126), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n734), .B(G101), .ZN(n736) );
  NOR2_X1 U783 ( .A1(n451), .A2(G898), .ZN(n735) );
  NOR2_X1 U784 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U785 ( .A(n738), .B(n737), .ZN(G69) );
  XOR2_X1 U786 ( .A(n740), .B(n739), .Z(n743) );
  XNOR2_X1 U787 ( .A(n741), .B(n743), .ZN(n742) );
  NAND2_X1 U788 ( .A1(n742), .A2(n451), .ZN(n747) );
  XNOR2_X1 U789 ( .A(n743), .B(G227), .ZN(n744) );
  NAND2_X1 U790 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U791 ( .A1(n745), .A2(G953), .ZN(n746) );
  NAND2_X1 U792 ( .A1(n747), .A2(n746), .ZN(G72) );
  XNOR2_X1 U793 ( .A(n748), .B(G143), .ZN(G45) );
  XOR2_X1 U794 ( .A(G110), .B(n749), .Z(G12) );
  XNOR2_X1 U795 ( .A(n750), .B(G131), .ZN(G33) );
endmodule

