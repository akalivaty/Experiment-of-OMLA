//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G902), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT24), .B(G110), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT64), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT64), .A2(G119), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(G128), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n192), .A2(new_n196), .A3(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n200), .B(KEYINPUT70), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT71), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(KEYINPUT71), .A3(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(KEYINPUT16), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n203), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n214), .A3(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT64), .A2(G119), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(new_n193), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n219), .B2(G128), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n198), .B1(new_n219), .B2(G128), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(new_n217), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G110), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n201), .A2(new_n216), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT72), .B(G110), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n220), .B(new_n225), .C1(new_n221), .C2(new_n217), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n196), .A2(new_n199), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n191), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT73), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n203), .A2(new_n205), .A3(new_n214), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(new_n212), .B2(G146), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n229), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n230), .B1(new_n229), .B2(new_n233), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n224), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT22), .B(G137), .ZN(new_n237));
  INV_X1    g051(.A(G953), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n238), .A2(G221), .A3(G234), .ZN(new_n239));
  XOR2_X1   g053(.A(new_n237), .B(new_n239), .Z(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n224), .B(new_n240), .C1(new_n234), .C2(new_n235), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n242), .A2(KEYINPUT75), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT75), .B1(new_n242), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n190), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT76), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT76), .B(new_n190), .C1(new_n244), .C2(new_n245), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n242), .A2(new_n188), .A3(new_n243), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT25), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n242), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n243), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(KEYINPUT74), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n250), .A2(new_n256), .A3(new_n251), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n189), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n248), .B(new_n249), .C1(new_n255), .C2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT1), .B1(new_n260), .B2(G146), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(G146), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n214), .A2(G143), .ZN(new_n263));
  OAI211_X1 g077(.A(G128), .B(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n214), .A2(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(G146), .ZN(new_n266));
  INV_X1    g080(.A(G128), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n265), .B(new_n266), .C1(KEYINPUT1), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT11), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(G137), .ZN(new_n274));
  INV_X1    g088(.A(G137), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT11), .A3(G134), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(G137), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n274), .A2(new_n276), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n273), .A2(G137), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n275), .A2(G134), .ZN(new_n281));
  OAI21_X1  g095(.A(G131), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n264), .A2(KEYINPUT65), .A3(new_n268), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n271), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT0), .A4(G128), .ZN(new_n288));
  XNOR2_X1  g102(.A(G143), .B(G146), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT0), .B(G128), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n274), .A2(new_n276), .A3(new_n278), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G131), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n279), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n271), .A2(KEYINPUT66), .A3(new_n283), .A4(new_n284), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n287), .A2(KEYINPUT30), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n283), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n296), .B1(new_n299), .B2(new_n269), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT30), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT2), .B(G113), .ZN(new_n302));
  INV_X1    g116(.A(G116), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n218), .A2(new_n193), .A3(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n197), .A2(G116), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n304), .ZN(new_n307));
  INV_X1    g121(.A(new_n305), .ZN(new_n308));
  INV_X1    g122(.A(new_n302), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n300), .A2(new_n301), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n298), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n291), .B1(new_n279), .B2(new_n294), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n306), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n287), .A2(new_n315), .A3(new_n297), .ZN(new_n316));
  INV_X1    g130(.A(G237), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT67), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G237), .ZN(new_n320));
  AOI21_X1  g134(.A(G953), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G210), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G101), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n324), .B(new_n325), .Z(new_n326));
  NAND3_X1  g140(.A1(new_n312), .A2(new_n316), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT31), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n312), .A2(KEYINPUT31), .A3(new_n316), .A4(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT28), .B1(new_n315), .B2(new_n285), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n300), .A2(new_n314), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n316), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n333), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n326), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT32), .ZN(new_n341));
  NOR2_X1   g155(.A1(G472), .A2(G902), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n329), .A2(new_n330), .B1(new_n337), .B2(new_n338), .ZN(new_n344));
  INV_X1    g158(.A(new_n342), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT32), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n287), .A2(new_n297), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n315), .A2(new_n349), .B1(new_n298), .B2(new_n311), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n348), .B1(new_n350), .B2(new_n326), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n336), .B1(new_n316), .B2(new_n334), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n352), .A2(new_n338), .A3(new_n332), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT69), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n333), .B(new_n326), .C1(new_n335), .C2(new_n336), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n312), .A2(new_n316), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n338), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT69), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n355), .A2(new_n357), .A3(new_n358), .A4(new_n348), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n287), .A2(new_n296), .A3(new_n297), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n314), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n316), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n332), .B1(new_n362), .B2(KEYINPUT28), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n338), .A2(new_n348), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n354), .A2(new_n359), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G472), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n259), .B1(new_n347), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT9), .B(G234), .ZN(new_n369));
  OAI21_X1  g183(.A(G221), .B1(new_n369), .B2(G902), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT82), .B(G469), .ZN(new_n371));
  XNOR2_X1  g185(.A(G110), .B(G140), .ZN(new_n372));
  INV_X1    g186(.A(G227), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G953), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n372), .B(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n264), .A2(new_n268), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT77), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(KEYINPUT77), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G104), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G107), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n377), .A2(new_n380), .A3(KEYINPUT77), .A4(G104), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n382), .A2(new_n383), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G104), .B(G107), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G101), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT81), .B1(new_n388), .B2(new_n383), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n376), .A2(new_n387), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n271), .A2(new_n284), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n387), .A2(new_n391), .A3(KEYINPUT10), .A4(new_n392), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT77), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(KEYINPUT3), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n384), .A2(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(KEYINPUT3), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n386), .A2(new_n385), .ZN(new_n404));
  OAI211_X1 g218(.A(KEYINPUT78), .B(G101), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT4), .A3(new_n387), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT78), .B1(new_n407), .B2(G101), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n292), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n410), .B(G101), .C1(new_n403), .C2(new_n404), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n407), .A2(KEYINPUT79), .A3(new_n410), .A4(G101), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT80), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G101), .B1(new_n403), .B2(new_n404), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT78), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n419), .A2(KEYINPUT4), .A3(new_n405), .A4(new_n387), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(new_n414), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT80), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n420), .A2(new_n421), .A3(new_n422), .A4(new_n292), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n398), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n295), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n295), .B(new_n398), .C1(new_n416), .C2(new_n423), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n375), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n387), .A2(new_n391), .A3(new_n392), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n269), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n393), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT12), .B1(new_n431), .B2(new_n295), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT12), .ZN(new_n433));
  AOI211_X1 g247(.A(new_n433), .B(new_n425), .C1(new_n430), .C2(new_n393), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT83), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n416), .A2(new_n423), .ZN(new_n438));
  INV_X1    g252(.A(new_n398), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n425), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n375), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT83), .B1(new_n432), .B2(new_n434), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n437), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  AOI211_X1 g257(.A(G902), .B(new_n371), .C1(new_n428), .C2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G469), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n441), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n435), .B1(new_n424), .B2(new_n425), .ZN(new_n447));
  OAI22_X1  g261(.A1(new_n446), .A2(new_n426), .B1(new_n447), .B2(new_n441), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n445), .B1(new_n448), .B2(new_n188), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n370), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G210), .B1(G237), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n292), .A2(G125), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(G125), .B2(new_n269), .ZN(new_n456));
  INV_X1    g270(.A(G224), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G953), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT87), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n456), .B(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT84), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT86), .B(KEYINPUT6), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n420), .A2(new_n314), .A3(new_n421), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n307), .A2(KEYINPUT5), .A3(new_n308), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n304), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n467), .A3(G113), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n391), .A2(new_n392), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n468), .A2(new_n310), .A3(new_n469), .A4(new_n387), .ZN(new_n470));
  AOI211_X1 g284(.A(new_n462), .B(new_n463), .C1(new_n464), .C2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n314), .B1(new_n406), .B2(new_n408), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n461), .B(new_n470), .C1(new_n472), .C2(new_n415), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n476), .A3(KEYINPUT6), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n464), .A2(new_n470), .ZN(new_n478));
  INV_X1    g292(.A(new_n462), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n460), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(new_n457), .B2(G953), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n456), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n455), .B(new_n483), .C1(G125), .C2(new_n269), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n468), .A2(new_n310), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n429), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n470), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n461), .B(KEYINPUT8), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n473), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n188), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n454), .B1(new_n482), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(G902), .B1(new_n492), .B2(new_n473), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n474), .A2(new_n471), .B1(new_n477), .B2(new_n480), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n496), .B(new_n453), .C1(new_n497), .C2(new_n460), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n452), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n450), .A2(new_n500), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n369), .A2(new_n187), .A3(G953), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n260), .A2(G128), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT93), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n260), .A2(G128), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n273), .A3(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(G116), .B(G122), .Z(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT92), .B(G107), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n510), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(new_n506), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n505), .A2(new_n514), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n517), .A2(KEYINPUT95), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(KEYINPUT95), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n513), .B1(new_n520), .B2(G134), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n505), .A2(new_n507), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G134), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n508), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n303), .A2(G122), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n380), .B1(new_n525), .B2(KEYINPUT14), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n526), .A2(new_n509), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n509), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n503), .B1(new_n521), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n517), .B(KEYINPUT95), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n273), .B1(new_n532), .B2(new_n516), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n529), .B(new_n502), .C1(new_n533), .C2(new_n513), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n188), .ZN(new_n536));
  INV_X1    g350(.A(G478), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(KEYINPUT15), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n531), .B2(new_n534), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(KEYINPUT15), .B2(new_n537), .ZN(new_n541));
  INV_X1    g355(.A(G952), .ZN(new_n542));
  AOI211_X1 g356(.A(G953), .B(new_n542), .C1(G234), .C2(G237), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT21), .B(G898), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT96), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AOI211_X1 g360(.A(new_n188), .B(new_n238), .C1(G234), .C2(G237), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n539), .A2(new_n541), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT91), .ZN(new_n551));
  NOR2_X1   g365(.A1(G475), .A2(G902), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n207), .A2(new_n208), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n231), .B1(new_n554), .B2(new_n214), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n319), .A2(G237), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n317), .A2(KEYINPUT67), .ZN(new_n557));
  OAI211_X1 g371(.A(G214), .B(new_n238), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n260), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n321), .A2(G143), .A3(G214), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT88), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT18), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n559), .B(new_n560), .C1(new_n277), .C2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n558), .A2(new_n260), .ZN(new_n564));
  AOI21_X1  g378(.A(G143), .B1(new_n321), .B2(G214), .ZN(new_n565));
  OAI21_X1  g379(.A(G131), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n555), .B(new_n563), .C1(new_n566), .C2(new_n562), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n559), .A2(new_n277), .A3(new_n560), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n277), .B1(new_n559), .B2(new_n560), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n213), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT19), .B1(new_n203), .B2(new_n205), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(new_n554), .B2(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT89), .B1(new_n572), .B2(G146), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT89), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT19), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n207), .B2(new_n208), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n574), .B(new_n214), .C1(new_n576), .C2(new_n571), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n567), .B1(new_n570), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(G113), .B(G122), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(new_n384), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT17), .ZN(new_n584));
  OAI211_X1 g398(.A(KEYINPUT17), .B(G131), .C1(new_n564), .C2(new_n565), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n213), .A3(new_n215), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n581), .B(new_n567), .C1(new_n584), .C2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n553), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT20), .B1(new_n588), .B2(KEYINPUT90), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT90), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n590), .B(new_n553), .C1(new_n583), .C2(new_n587), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n587), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n559), .A2(new_n277), .A3(new_n560), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n566), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n595), .A2(new_n213), .A3(new_n573), .A4(new_n577), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n581), .B1(new_n596), .B2(new_n567), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n552), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT20), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n590), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n566), .A2(new_n601), .A3(new_n594), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n602), .A2(new_n213), .A3(new_n215), .A4(new_n585), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n581), .B1(new_n603), .B2(new_n567), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n188), .B1(new_n593), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G475), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n551), .B1(new_n592), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n583), .A2(new_n587), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT90), .B1(new_n609), .B2(new_n552), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n610), .A2(new_n599), .B1(G475), .B2(new_n605), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n598), .A2(new_n590), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n588), .A2(KEYINPUT90), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(KEYINPUT20), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n614), .A3(KEYINPUT91), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n550), .B1(new_n608), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n368), .A2(new_n501), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  NAND2_X1  g432(.A1(new_n535), .A2(KEYINPUT33), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n531), .A2(new_n620), .A3(new_n534), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(G478), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n537), .A2(new_n188), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n540), .B2(new_n537), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n608), .A2(new_n615), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n475), .A2(new_n481), .ZN(new_n627));
  INV_X1    g441(.A(new_n460), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n453), .B1(new_n629), .B2(new_n496), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n482), .A2(new_n494), .A3(new_n454), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n549), .B(new_n451), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n633), .A2(KEYINPUT97), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(KEYINPUT97), .ZN(new_n635));
  INV_X1    g449(.A(new_n259), .ZN(new_n636));
  INV_X1    g450(.A(new_n370), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n440), .B1(new_n434), .B2(new_n432), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n424), .A2(new_n425), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n375), .B1(new_n424), .B2(new_n425), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n638), .A2(new_n375), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(G469), .B1(new_n641), .B2(G902), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n428), .A2(new_n443), .ZN(new_n643));
  INV_X1    g457(.A(new_n371), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n188), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n637), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n331), .B2(new_n339), .ZN(new_n647));
  INV_X1    g461(.A(G472), .ZN(new_n648));
  OAI22_X1  g462(.A1(new_n647), .A2(new_n648), .B1(new_n345), .B2(new_n344), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n636), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n634), .A2(new_n635), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G104), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  NAND2_X1  g470(.A1(new_n611), .A2(new_n614), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n539), .A2(new_n541), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n499), .A2(new_n658), .A3(new_n549), .A4(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT35), .B(G107), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  OR3_X1    g477(.A1(new_n236), .A2(KEYINPUT36), .A3(new_n241), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n236), .B1(KEYINPUT36), .B2(new_n241), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n664), .A2(new_n190), .A3(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n257), .A2(new_n189), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n666), .B1(new_n667), .B2(new_n254), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(new_n616), .A3(new_n646), .A4(new_n499), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NAND2_X1  g486(.A1(new_n347), .A2(new_n367), .ZN(new_n673));
  INV_X1    g487(.A(new_n668), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n673), .A2(new_n646), .A3(new_n499), .A4(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n543), .B1(new_n547), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n659), .A2(new_n614), .A3(new_n611), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT99), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n267), .ZN(G30));
  NAND2_X1  g496(.A1(new_n495), .A2(new_n498), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n608), .A2(new_n615), .ZN(new_n690));
  INV_X1    g504(.A(new_n659), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n674), .A2(new_n690), .A3(new_n691), .A4(new_n452), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n688), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n689), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n677), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n646), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n356), .A2(new_n326), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n698), .B(new_n188), .C1(new_n326), .C2(new_n362), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n343), .A2(new_n346), .B1(G472), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT101), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n694), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n260), .ZN(G45));
  AND4_X1   g518(.A1(new_n673), .A2(new_n646), .A3(new_n499), .A4(new_n674), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n608), .A2(new_n615), .A3(new_n625), .A4(new_n678), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  NAND3_X1  g523(.A1(new_n643), .A2(KEYINPUT103), .A3(new_n188), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  AOI21_X1  g525(.A(G902), .B1(new_n428), .B2(new_n443), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(KEYINPUT103), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n370), .B(new_n645), .C1(new_n711), .C2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n634), .A2(new_n635), .A3(new_n715), .A4(new_n368), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND2_X1  g532(.A1(new_n673), .A2(new_n636), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n719), .A2(new_n714), .A3(new_n660), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n303), .ZN(G18));
  OR2_X1    g535(.A1(new_n712), .A2(KEYINPUT103), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n445), .B1(new_n712), .B2(KEYINPUT103), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n444), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n370), .A3(new_n499), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n673), .A2(new_n616), .A3(new_n674), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n197), .ZN(G21));
  OAI21_X1  g542(.A(new_n331), .B1(new_n326), .B2(new_n363), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n342), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n340), .A2(new_n188), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n731), .B1(new_n732), .B2(G472), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n647), .A2(KEYINPUT104), .A3(new_n648), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n259), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n667), .A2(new_n254), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(KEYINPUT105), .A3(new_n248), .A4(new_n249), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n735), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n608), .A2(new_n615), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n548), .B(new_n452), .C1(new_n495), .C2(new_n498), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n659), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n714), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  NAND3_X1  g560(.A1(new_n732), .A2(new_n731), .A3(G472), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT104), .B1(new_n647), .B2(new_n648), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n707), .A2(new_n674), .A3(new_n730), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n725), .ZN(new_n751));
  XOR2_X1   g565(.A(KEYINPUT106), .B(G125), .Z(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G27));
  NAND2_X1  g567(.A1(new_n737), .A2(new_n739), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n673), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n683), .A2(new_n452), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n646), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n758), .A2(new_n759), .A3(new_n706), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n719), .A2(new_n758), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT107), .B1(new_n762), .B2(new_n707), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n684), .A2(new_n451), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n450), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(new_n368), .A3(KEYINPUT107), .A4(new_n707), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n759), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n761), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n765), .A2(new_n368), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(new_n772), .B2(new_n706), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n759), .A3(new_n766), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT108), .B1(new_n774), .B2(new_n761), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NOR2_X1   g591(.A1(new_n772), .A2(new_n680), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT109), .B(G134), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G36));
  NAND2_X1  g594(.A1(new_n690), .A2(new_n625), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT43), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n690), .A2(new_n783), .A3(new_n625), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n650), .A2(new_n668), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n785), .A2(KEYINPUT44), .A3(new_n786), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n757), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n445), .B1(new_n448), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n641), .A2(KEYINPUT45), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n793), .A2(new_n794), .B1(G469), .B2(G902), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n795), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT110), .B1(new_n795), .B2(KEYINPUT46), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n444), .B1(new_n795), .B2(KEYINPUT46), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n370), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n695), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n791), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(new_n275), .ZN(G39));
  NAND2_X1  g617(.A1(new_n799), .A2(new_n370), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n804), .B1(new_n805), .B2(KEYINPUT47), .ZN(new_n806));
  XNOR2_X1  g620(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n799), .A2(new_n370), .A3(new_n808), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n673), .A2(new_n636), .A3(new_n764), .A4(new_n706), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  XNOR2_X1  g626(.A(new_n659), .B(KEYINPUT113), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n742), .A3(new_n690), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n670), .B1(new_n651), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n720), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n714), .A2(new_n500), .ZN(new_n817));
  INV_X1    g631(.A(new_n726), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n740), .A2(new_n744), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n816), .A2(new_n819), .A3(new_n716), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n450), .A2(new_n259), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n633), .A3(new_n650), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n617), .A2(new_n822), .A3(KEYINPUT112), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT112), .B1(new_n617), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n768), .A2(new_n769), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n774), .A2(KEYINPUT108), .A3(new_n761), .ZN(new_n828));
  INV_X1    g642(.A(new_n813), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n658), .A3(new_n678), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n673), .A2(new_n674), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n750), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n778), .B1(new_n765), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n826), .A2(new_n827), .A3(new_n828), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n735), .A2(new_n668), .A3(new_n706), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n679), .B(KEYINPUT99), .Z(new_n837));
  AOI22_X1  g651(.A1(new_n836), .A2(new_n817), .B1(new_n705), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n699), .A2(G472), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n347), .A2(new_n839), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n666), .B(new_n677), .C1(new_n667), .C2(new_n254), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n840), .A2(new_n646), .A3(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n500), .A2(new_n690), .A3(new_n691), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n705), .A2(new_n707), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n835), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  OAI22_X1  g659(.A1(new_n750), .A2(new_n725), .B1(new_n675), .B2(new_n680), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n840), .A2(new_n646), .A3(new_n841), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n741), .A2(new_n659), .A3(new_n499), .ZN(new_n848));
  OAI22_X1  g662(.A1(new_n675), .A2(new_n706), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n846), .A2(new_n849), .A3(KEYINPUT52), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT114), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n838), .A2(new_n844), .A3(new_n835), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT52), .B1(new_n846), .B2(new_n849), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT53), .B1(new_n834), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n832), .A2(new_n765), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n820), .A2(new_n825), .A3(new_n858), .A4(new_n778), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n845), .A2(new_n850), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n859), .A2(new_n776), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n857), .A2(KEYINPUT54), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n860), .B1(new_n834), .B2(new_n856), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n768), .A4(new_n861), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n782), .A2(new_n543), .A3(new_n784), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n714), .A2(new_n764), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n756), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT48), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n817), .A3(new_n740), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n542), .A2(G953), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n626), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n636), .A2(new_n543), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n701), .A2(new_n869), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n872), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n878), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n871), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n735), .A2(new_n668), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n868), .A2(new_n882), .A3(new_n869), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n741), .A2(new_n625), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n701), .A2(new_n869), .A3(new_n877), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n452), .B1(new_n686), .B2(new_n687), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n714), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n868), .A3(new_n740), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT50), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n888), .A2(new_n868), .A3(KEYINPUT50), .A4(new_n740), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n806), .A2(new_n809), .B1(new_n637), .B2(new_n724), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n868), .A2(new_n740), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT115), .B1(new_n895), .B2(new_n764), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n868), .A2(new_n897), .A3(new_n740), .A4(new_n757), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n893), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT51), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT51), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n893), .B(new_n902), .C1(new_n894), .C2(new_n899), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n881), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n863), .A2(new_n867), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n542), .A2(new_n238), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n688), .ZN(new_n908));
  NOR4_X1   g722(.A1(new_n908), .A2(new_n637), .A3(new_n452), .A4(new_n781), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n724), .B(KEYINPUT49), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n909), .A2(new_n701), .A3(new_n754), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT117), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n907), .A2(new_n914), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n238), .A2(G952), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n188), .B1(new_n864), .B2(new_n866), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(G210), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n497), .A2(new_n460), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n629), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT55), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n917), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT118), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n918), .A2(KEYINPUT118), .A3(G210), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n924), .A2(KEYINPUT56), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n925), .A2(new_n930), .ZN(G51));
  NAND2_X1  g745(.A1(G469), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT57), .Z(new_n933));
  INV_X1    g747(.A(new_n867), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n643), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n918), .A2(new_n794), .A3(new_n793), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n917), .B1(new_n937), .B2(new_n938), .ZN(G54));
  NAND3_X1  g753(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n940));
  INV_X1    g754(.A(new_n609), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n917), .ZN(G60));
  NAND2_X1  g758(.A1(new_n619), .A2(new_n621), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n623), .B(KEYINPUT59), .Z(new_n946));
  OAI211_X1 g760(.A(new_n945), .B(new_n946), .C1(new_n934), .C2(new_n935), .ZN(new_n947));
  INV_X1    g761(.A(new_n917), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n863), .A2(new_n867), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n950), .B2(new_n946), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(G63));
  OAI21_X1  g766(.A(new_n948), .B1(KEYINPUT120), .B2(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n864), .A2(new_n866), .ZN(new_n954));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT119), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n244), .A2(new_n245), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n954), .A2(new_n664), .A3(new_n665), .A4(new_n957), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(G66));
  AOI21_X1  g779(.A(new_n238), .B1(new_n545), .B2(G224), .ZN(new_n966));
  INV_X1    g780(.A(new_n826), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(new_n238), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n497), .B1(G898), .B2(new_n238), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT121), .Z(new_n970));
  XNOR2_X1  g784(.A(new_n968), .B(new_n970), .ZN(G69));
  NAND2_X1  g785(.A1(new_n300), .A2(new_n301), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n298), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(new_n572), .Z(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n838), .A2(new_n708), .ZN(new_n976));
  OAI21_X1  g790(.A(KEYINPUT124), .B1(new_n802), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n978));
  INV_X1    g792(.A(new_n976), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n978), .B(new_n979), .C1(new_n791), .C2(new_n801), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n800), .A2(new_n695), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n755), .A2(new_n848), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n778), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n776), .A2(new_n984), .A3(new_n811), .ZN(new_n985));
  AOI21_X1  g799(.A(G953), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n676), .A2(G953), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT123), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n975), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n626), .B1(new_n829), .B2(new_n741), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n762), .A2(new_n695), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n802), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n979), .B(new_n994), .C1(new_n694), .C2(new_n702), .ZN(new_n995));
  OAI21_X1  g809(.A(KEYINPUT62), .B1(new_n703), .B2(new_n976), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n993), .A2(new_n811), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n238), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n974), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n990), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(G953), .B1(new_n373), .B2(new_n676), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT122), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1000), .B(new_n1003), .ZN(G72));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT63), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(new_n357), .B2(new_n327), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n857), .A2(new_n862), .A3(new_n1007), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1006), .B(KEYINPUT125), .Z(new_n1009));
  OAI21_X1  g823(.A(new_n1009), .B1(new_n997), .B2(new_n967), .ZN(new_n1010));
  INV_X1    g824(.A(new_n698), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n1010), .A2(KEYINPUT126), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(KEYINPUT126), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n948), .B(new_n1008), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n350), .A2(new_n338), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n981), .A2(new_n985), .A3(new_n826), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n1009), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(KEYINPUT127), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1016), .A2(new_n1019), .A3(new_n1009), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1015), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1014), .A2(new_n1021), .ZN(G57));
endmodule


