//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  INV_X1    g000(.A(G36gat), .ZN(new_n202));
  AND2_X1   g001(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n210));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n210), .A2(new_n211), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT17), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT91), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(G1gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT90), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n218), .B(new_n219), .C1(G1gat), .C2(new_n216), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(G8gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT17), .B1(new_n212), .B2(new_n213), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(KEYINPUT89), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(KEYINPUT89), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n215), .A2(new_n222), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n213), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT92), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n226), .A2(KEYINPUT18), .A3(new_n227), .A4(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n221), .A2(new_n228), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n227), .B(KEYINPUT13), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT11), .B(G169gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT12), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n231), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n227), .A3(new_n230), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT93), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT93), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n246), .A3(new_n243), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n241), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n240), .ZN(new_n249));
  INV_X1    g048(.A(new_n244), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT85), .ZN(new_n255));
  XNOR2_X1  g054(.A(G78gat), .B(G106gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G22gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G228gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT2), .ZN(new_n264));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(KEYINPUT80), .A3(new_n263), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n270));
  INV_X1    g069(.A(new_n263), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(new_n271), .B2(new_n267), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n266), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n271), .A2(new_n267), .ZN(new_n274));
  INV_X1    g073(.A(new_n265), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(new_n261), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n274), .A2(new_n276), .A3(KEYINPUT80), .A4(new_n264), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT22), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT74), .B(G211gat), .ZN(new_n282));
  INV_X1    g081(.A(G218gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285));
  XNOR2_X1  g084(.A(G197gat), .B(G204gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n280), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n289), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n287), .A3(new_n279), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT84), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT3), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n290), .A2(new_n292), .A3(KEYINPUT84), .A4(new_n293), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n278), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT3), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n278), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n290), .A2(new_n292), .B1(new_n293), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n260), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n278), .B1(new_n294), .B2(new_n299), .ZN(new_n303));
  OR3_X1    g102(.A1(new_n303), .A2(new_n301), .A3(new_n260), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT31), .B(G50gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n302), .B2(new_n304), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n258), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n302), .A2(new_n304), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n305), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n312), .A2(new_n257), .A3(new_n307), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G1gat), .B(G29gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT0), .ZN(new_n317));
  XNOR2_X1  g116(.A(G57gat), .B(G85gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT69), .B(G134gat), .Z(new_n323));
  INV_X1    g122(.A(G127gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(G127gat), .A2(G134gat), .ZN(new_n326));
  INV_X1    g125(.A(G113gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G120gat), .ZN(new_n328));
  INV_X1    g127(.A(G120gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G113gat), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT1), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n325), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n326), .ZN(new_n334));
  NAND2_X1  g133(.A1(G127gat), .A2(G134gat), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT1), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(KEYINPUT70), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G120gat), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT71), .A4(G113gat), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT72), .B1(new_n329), .B2(G113gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n327), .A3(G120gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT70), .B(G120gat), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT71), .B1(new_n345), .B2(G113gat), .ZN(new_n346));
  OAI211_X1 g145(.A(KEYINPUT73), .B(new_n336), .C1(new_n344), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n337), .A2(new_n339), .A3(G113gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n341), .A2(new_n343), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n340), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT73), .B1(new_n353), .B2(new_n336), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n333), .B(new_n278), .C1(new_n348), .C2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n336), .B1(new_n344), .B2(new_n346), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n332), .B1(new_n358), .B2(new_n347), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n273), .A2(new_n277), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT3), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n300), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n355), .B(KEYINPUT4), .C1(new_n359), .C2(new_n362), .ZN(new_n363));
  AOI211_X1 g162(.A(new_n332), .B(new_n360), .C1(new_n358), .C2(new_n347), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n322), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n333), .B1(new_n348), .B2(new_n354), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n360), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n321), .B1(new_n370), .B2(new_n355), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT5), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n347), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n278), .B1(new_n374), .B2(new_n333), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n322), .B1(new_n375), .B2(new_n364), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n367), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n367), .A2(new_n372), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(KEYINPUT6), .B(new_n320), .C1(new_n378), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT82), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n363), .A2(new_n366), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n321), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n371), .A2(new_n368), .A3(new_n372), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT81), .B1(new_n376), .B2(KEYINPUT5), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n379), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT6), .A4(new_n320), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT6), .B1(new_n388), .B2(new_n320), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n379), .A3(new_n319), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n382), .A2(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n290), .A2(new_n292), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT27), .B(G183gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT28), .ZN(new_n396));
  AOI21_X1  g195(.A(G190gat), .B1(new_n396), .B2(KEYINPUT67), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n396), .A2(KEYINPUT67), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(G169gat), .B2(G176gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(G169gat), .A2(G176gat), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n405), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT68), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n404), .A2(new_n406), .A3(KEYINPUT68), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n402), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n405), .A2(KEYINPUT23), .ZN(new_n413));
  NAND2_X1  g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT23), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(G169gat), .B2(G176gat), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G183gat), .A2(G190gat), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT24), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G183gat), .ZN(new_n422));
  INV_X1    g221(.A(G190gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT64), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT64), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(G183gat), .B2(G190gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n421), .A2(new_n424), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT25), .B1(new_n418), .B2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n413), .A2(KEYINPUT25), .A3(new_n416), .A4(new_n414), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n419), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n431));
  AND2_X1   g230(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n422), .A2(new_n423), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n434), .A2(new_n427), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n430), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n412), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n438), .B(KEYINPUT76), .Z(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT66), .B1(new_n429), .B2(new_n436), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n435), .B1(new_n432), .B2(new_n431), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT25), .A3(new_n418), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT25), .ZN(new_n444));
  AND4_X1   g243(.A1(new_n421), .A2(new_n424), .A3(new_n426), .A4(new_n427), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n417), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT66), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n441), .A2(new_n448), .B1(new_n411), .B2(new_n402), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n439), .A2(KEYINPUT29), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  OAI221_X1 g250(.A(new_n394), .B1(new_n437), .B2(new_n440), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n402), .A2(new_n411), .B1(new_n443), .B2(new_n446), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n440), .B1(new_n453), .B2(KEYINPUT29), .ZN(new_n454));
  INV_X1    g253(.A(new_n394), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n454), .B(new_n455), .C1(new_n449), .C2(new_n440), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G8gat), .B(G36gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT77), .ZN(new_n459));
  XOR2_X1   g258(.A(G64gat), .B(G92gat), .Z(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(KEYINPUT79), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n452), .A2(new_n456), .A3(new_n461), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT79), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n461), .B(KEYINPUT78), .Z(new_n468));
  NOR2_X1   g267(.A1(new_n457), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n464), .A2(new_n463), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT83), .B1(new_n393), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n390), .A2(new_n382), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n320), .B1(new_n378), .B2(new_n380), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n392), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n479));
  INV_X1    g278(.A(new_n472), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n315), .B1(new_n473), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483));
  XOR2_X1   g282(.A(G15gat), .B(G43gat), .Z(new_n484));
  XNOR2_X1  g283(.A(G71gat), .B(G99gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n441), .A2(new_n448), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n412), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n359), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n449), .A2(new_n369), .ZN(new_n491));
  AND2_X1   g290(.A1(G227gat), .A2(G233gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n492), .B1(new_n490), .B2(new_n491), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT34), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI211_X1 g298(.A(KEYINPUT34), .B(new_n492), .C1(new_n490), .C2(new_n491), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n493), .A2(KEYINPUT32), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n497), .A2(new_n498), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n495), .B1(new_n505), .B2(new_n500), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n504), .B1(new_n502), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n483), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n506), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n495), .A2(new_n505), .A3(new_n500), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n503), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(KEYINPUT36), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n255), .B1(new_n482), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n479), .B1(new_n478), .B2(new_n480), .ZN(new_n517));
  AOI211_X1 g316(.A(KEYINPUT83), .B(new_n472), .C1(new_n474), .C2(new_n477), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n314), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n509), .A2(new_n514), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(KEYINPUT85), .A3(new_n520), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n383), .A2(KEYINPUT39), .A3(new_n321), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(new_n320), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n370), .A2(new_n355), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT39), .B1(new_n524), .B2(new_n322), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT86), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n321), .B2(new_n383), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n525), .A2(new_n526), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n523), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT40), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n472), .A2(new_n475), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n468), .A2(KEYINPUT38), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n452), .A2(new_n456), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(KEYINPUT37), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n449), .A2(new_n451), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n437), .A2(new_n440), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n455), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(KEYINPUT87), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n454), .B1(new_n440), .B2(new_n449), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n394), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(KEYINPUT87), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n536), .B1(new_n544), .B2(KEYINPUT37), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT38), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n461), .B1(new_n457), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n535), .A2(KEYINPUT37), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n462), .A2(new_n466), .ZN(new_n551));
  OR3_X1    g350(.A1(new_n545), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n533), .B(new_n315), .C1(new_n478), .C2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n516), .A2(new_n521), .A3(new_n553), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n314), .A2(new_n507), .A3(new_n508), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n473), .A2(new_n481), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n507), .B2(new_n508), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n512), .A2(KEYINPUT88), .A3(new_n513), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n314), .A2(KEYINPUT35), .ZN(new_n562));
  AND4_X1   g361(.A1(new_n478), .A2(new_n561), .A3(new_n562), .A4(new_n480), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n254), .B1(new_n554), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G57gat), .B(G64gat), .Z(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(KEYINPUT94), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(KEYINPUT9), .B2(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI221_X1 g372(.A(new_n570), .B1(KEYINPUT9), .B2(new_n567), .C1(new_n569), .C2(KEYINPUT94), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(G127gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n221), .B1(KEYINPUT21), .B2(new_n575), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n578), .A2(G127gat), .ZN(new_n582));
  OR3_X1    g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n580), .B2(new_n582), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G155gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n585), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT96), .ZN(new_n592));
  AND2_X1   g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n593), .A2(KEYINPUT41), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT7), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n600), .B1(KEYINPUT8), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n598), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n215), .A2(new_n224), .A3(new_n225), .A4(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n604), .B(new_n605), .Z(new_n608));
  AOI22_X1  g407(.A1(new_n228), .A2(new_n608), .B1(KEYINPUT41), .B2(new_n593), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n591), .A2(KEYINPUT96), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n613), .B1(new_n610), .B2(new_n611), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n596), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(new_n595), .A3(new_n614), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n608), .A2(new_n575), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n574), .A3(new_n573), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n575), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n621), .A2(new_n623), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G120gat), .B(G148gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT98), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n630), .A2(new_n632), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n590), .A2(new_n620), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT99), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n393), .A2(KEYINPUT100), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n393), .A2(KEYINPUT100), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n566), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g449(.A1(new_n644), .A2(new_n480), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n566), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(G8gat), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n217), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n653), .B1(new_n566), .B2(new_n651), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT42), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(KEYINPUT42), .B2(new_n656), .ZN(G1325gat));
  NAND2_X1  g458(.A1(new_n566), .A2(new_n645), .ZN(new_n660));
  INV_X1    g459(.A(G15gat), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n520), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT103), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n660), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n561), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n661), .B1(new_n660), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT101), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT101), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n665), .B1(new_n668), .B2(new_n669), .ZN(G1326gat));
  NOR2_X1   g469(.A1(new_n660), .A2(new_n315), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT43), .B(G22gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  NOR3_X1   g472(.A1(new_n590), .A2(new_n620), .A3(new_n641), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n566), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n648), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n675), .A2(G29gat), .A3(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(KEYINPUT45), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n620), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n554), .B2(new_n565), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n519), .A2(new_n663), .A3(new_n553), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n565), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n617), .A2(new_n619), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT44), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n585), .B(new_n589), .Z(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n253), .A3(new_n642), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT104), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n682), .A2(new_n686), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n676), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT45), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n693), .A3(new_n694), .ZN(G1328gat));
  NOR3_X1   g494(.A1(new_n675), .A2(G36gat), .A3(new_n480), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n692), .B2(new_n480), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n697), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(G1329gat));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702));
  INV_X1    g501(.A(G43gat), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n663), .B(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(new_n691), .B2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n675), .A2(G43gat), .A3(new_n666), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n702), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n554), .A2(new_n565), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n680), .ZN(new_n710));
  INV_X1    g509(.A(new_n663), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n515), .A2(new_n662), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n520), .A2(KEYINPUT102), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n553), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n482), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n563), .B1(new_n556), .B2(KEYINPUT35), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n679), .B1(new_n717), .B2(new_n620), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n710), .A2(new_n711), .A3(new_n718), .A4(new_n689), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G43gat), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n709), .A2(new_n253), .A3(new_n674), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n666), .A2(G43gat), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n702), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n720), .A2(KEYINPUT105), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT105), .B1(new_n720), .B2(new_n723), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n708), .B1(new_n724), .B2(new_n725), .ZN(G1330gat));
  INV_X1    g525(.A(G50gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n721), .A2(new_n727), .A3(new_n314), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT48), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n710), .A2(new_n314), .A3(new_n718), .A4(new_n689), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G50gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n728), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n732), .B(new_n728), .C1(new_n729), .C2(KEYINPUT48), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1331gat));
  NAND4_X1  g535(.A1(new_n254), .A2(new_n590), .A3(new_n620), .A4(new_n641), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT107), .Z(new_n738));
  NAND2_X1  g537(.A1(new_n684), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT108), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n684), .A2(new_n741), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n676), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g544(.A1(new_n743), .A2(new_n480), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  AND2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n746), .B2(new_n747), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n743), .B2(new_n664), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n666), .A2(G71gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n740), .A2(new_n742), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n751), .A2(KEYINPUT50), .A3(new_n753), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1334gat));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n315), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(G78gat), .Z(G1335gat));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n590), .A2(new_n253), .A3(new_n642), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n710), .A2(new_n648), .A3(new_n718), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G85gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n590), .A2(new_n253), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n685), .B(new_n766), .C1(new_n715), .C2(new_n716), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n684), .A2(KEYINPUT51), .A3(new_n685), .A4(new_n766), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n767), .A2(KEYINPUT109), .A3(new_n768), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n676), .A2(G85gat), .A3(new_n642), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n761), .B1(new_n765), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n772), .A2(new_n773), .ZN(new_n777));
  INV_X1    g576(.A(new_n774), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n764), .B(KEYINPUT110), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1336gat));
  NAND4_X1  g579(.A1(new_n710), .A2(new_n472), .A3(new_n718), .A4(new_n762), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(new_n781), .B2(G92gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n480), .A2(G92gat), .A3(new_n642), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n777), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n770), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n781), .A2(G92gat), .B1(new_n787), .B2(new_n783), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n786), .B2(new_n788), .ZN(G1337gat));
  NAND4_X1  g588(.A1(new_n710), .A2(new_n705), .A3(new_n718), .A4(new_n762), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G99gat), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n666), .A2(G99gat), .A3(new_n642), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n777), .B2(new_n792), .ZN(G1338gat));
  NAND4_X1  g592(.A1(new_n710), .A2(new_n314), .A3(new_n718), .A4(new_n762), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT53), .B1(new_n794), .B2(G106gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n315), .A2(G106gat), .A3(new_n642), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n777), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n794), .A2(G106gat), .B1(new_n787), .B2(new_n796), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n233), .A2(new_n234), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n227), .B1(new_n226), .B2(new_n230), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n239), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n248), .A2(new_n641), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n624), .A2(new_n625), .A3(new_n628), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n630), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n637), .B1(new_n630), .B2(KEYINPUT54), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n810), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n813), .A3(new_n640), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n248), .B2(new_n252), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n620), .B1(new_n805), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n814), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n685), .A2(new_n248), .A3(new_n817), .A4(new_n804), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n590), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NOR4_X1   g618(.A1(new_n687), .A2(new_n685), .A3(new_n253), .A4(new_n641), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n314), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(new_n480), .A3(new_n561), .A4(new_n648), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n823), .A2(KEYINPUT111), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(KEYINPUT111), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n254), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n821), .A2(new_n676), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(new_n555), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n480), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n253), .A2(new_n327), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT112), .Z(new_n832));
  OAI21_X1  g631(.A(new_n827), .B1(new_n830), .B2(new_n832), .ZN(G1340gat));
  OAI21_X1  g632(.A(G120gat), .B1(new_n826), .B2(new_n642), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n641), .A2(new_n345), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n834), .B1(new_n830), .B2(new_n835), .ZN(G1341gat));
  NOR2_X1   g635(.A1(new_n687), .A2(new_n324), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n824), .A2(new_n825), .A3(new_n837), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n838), .A2(KEYINPUT113), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n324), .B1(new_n830), .B2(new_n687), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(KEYINPUT113), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(G1342gat));
  NAND2_X1  g641(.A1(new_n685), .A2(new_n480), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT114), .Z(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n323), .A3(new_n845), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT56), .Z(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n826), .B2(new_n620), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1343gat));
  NOR2_X1   g648(.A1(new_n705), .A2(new_n315), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n254), .A2(G141gat), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n850), .A2(new_n480), .A3(new_n828), .A4(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n663), .A2(new_n648), .A3(new_n480), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n315), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n805), .B2(new_n815), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n253), .A2(new_n817), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n248), .A2(new_n641), .A3(new_n804), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(KEYINPUT116), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n862), .A3(new_n620), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n590), .B1(new_n863), .B2(new_n818), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n857), .B1(new_n864), .B2(new_n820), .ZN(new_n865));
  XOR2_X1   g664(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n821), .B2(new_n315), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n254), .B(new_n855), .C1(new_n865), .C2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G141gat), .B1(new_n868), .B2(KEYINPUT117), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n855), .B1(new_n865), .B2(new_n867), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n870), .A2(KEYINPUT117), .A3(new_n253), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n854), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT118), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n854), .B(new_n874), .C1(new_n869), .C2(new_n871), .ZN(new_n875));
  INV_X1    g674(.A(G141gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n852), .B1(new_n868), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT58), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(new_n875), .A3(new_n878), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n850), .A2(new_n828), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n472), .ZN(new_n881));
  INV_X1    g680(.A(G148gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n641), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n819), .A2(new_n820), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n314), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n886), .A2(new_n866), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n644), .A2(new_n253), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n314), .B1(new_n888), .B2(new_n864), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n856), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n855), .A2(new_n642), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n884), .B1(new_n893), .B2(G148gat), .ZN(new_n894));
  AOI211_X1 g693(.A(KEYINPUT59), .B(new_n882), .C1(new_n870), .C2(new_n641), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n883), .B1(new_n894), .B2(new_n895), .ZN(G1345gat));
  NOR2_X1   g695(.A1(new_n687), .A2(G155gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n870), .A2(new_n590), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n881), .A2(new_n897), .B1(G155gat), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n899), .B(new_n900), .ZN(G1346gat));
  NOR3_X1   g700(.A1(new_n880), .A2(G162gat), .A3(new_n844), .ZN(new_n902));
  INV_X1    g701(.A(G162gat), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n903), .B1(new_n870), .B2(new_n685), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT120), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n648), .A2(new_n480), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n822), .A2(new_n561), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(G169gat), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(new_n909), .A3(new_n254), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n885), .A2(new_n676), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n555), .A2(new_n472), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT121), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n253), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n910), .B1(new_n915), .B2(new_n909), .ZN(G1348gat));
  NOR2_X1   g715(.A1(new_n642), .A2(G176gat), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G176gat), .B1(new_n908), .B2(new_n642), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(KEYINPUT122), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1349gat));
  AND2_X1   g723(.A1(new_n590), .A2(new_n395), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n913), .A2(new_n925), .B1(new_n926), .B2(KEYINPUT60), .ZN(new_n927));
  OAI21_X1  g726(.A(G183gat), .B1(new_n908), .B2(new_n687), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n926), .A2(KEYINPUT60), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n929), .B(new_n930), .Z(G1350gat));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n423), .A3(new_n685), .ZN(new_n932));
  OAI21_X1  g731(.A(G190gat), .B1(new_n908), .B2(new_n620), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(KEYINPUT61), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(KEYINPUT61), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(G1351gat));
  NOR3_X1   g735(.A1(new_n705), .A2(new_n480), .A3(new_n315), .ZN(new_n937));
  INV_X1    g736(.A(new_n911), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n253), .A3(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G197gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n664), .A2(new_n907), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n887), .B2(new_n890), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n254), .A2(new_n944), .ZN(new_n947));
  AOI22_X1  g746(.A1(new_n943), .A2(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n641), .ZN(new_n949));
  XOR2_X1   g748(.A(KEYINPUT125), .B(G204gat), .Z(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n642), .A2(new_n951), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n937), .A2(new_n938), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n938), .A3(new_n956), .ZN(new_n958));
  XOR2_X1   g757(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n952), .A2(KEYINPUT127), .A3(new_n957), .A4(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n957), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n950), .B1(new_n946), .B2(new_n641), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n961), .A2(new_n965), .ZN(G1353gat));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n590), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n967), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n941), .A2(new_n942), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n590), .A2(new_n282), .ZN(new_n971));
  OAI22_X1  g770(.A1(new_n968), .A2(new_n969), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  NAND2_X1  g771(.A1(new_n685), .A2(new_n283), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n946), .A2(new_n685), .ZN(new_n974));
  OAI22_X1  g773(.A1(new_n970), .A2(new_n973), .B1(new_n283), .B2(new_n974), .ZN(G1355gat));
endmodule


