//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018;
  XNOR2_X1  g000(.A(G71gat), .B(G78gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT97), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205));
  NOR3_X1   g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(KEYINPUT97), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g007(.A(KEYINPUT97), .B(new_n202), .C1(new_n205), .C2(new_n204), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT21), .ZN(new_n211));
  NAND2_X1  g010(.A1(G231gat), .A2(G233gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G183gat), .B(G211gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G1gat), .B2(new_n218), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(G8gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(KEYINPUT21), .B2(new_n210), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT98), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n224), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n217), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(G190gat), .B(G218gat), .Z(new_n230));
  NAND3_X1  g029(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT14), .ZN(new_n232));
  INV_X1    g031(.A(G29gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n235));
  AOI21_X1  g034(.A(G36gat), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G36gat), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n232), .A2(new_n237), .A3(G29gat), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G43gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G50gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT90), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT15), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G50gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G43gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n241), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n249), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n239), .A2(new_n251), .A3(new_n245), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n238), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n244), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G85gat), .A2(G92gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT7), .ZN(new_n257));
  XNOR2_X1  g056(.A(G99gat), .B(G106gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(G99gat), .A2(G106gat), .ZN(new_n259));
  INV_X1    g058(.A(G85gat), .ZN(new_n260));
  INV_X1    g059(.A(G92gat), .ZN(new_n261));
  AOI22_X1  g060(.A1(KEYINPUT8), .A2(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n257), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n257), .B2(new_n262), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n231), .B1(new_n255), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT100), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT17), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n250), .A2(new_n269), .A3(new_n252), .A4(new_n254), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n265), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT91), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n272), .B1(new_n255), .B2(KEYINPUT17), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n255), .A2(new_n272), .A3(KEYINPUT17), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n230), .B1(new_n268), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n266), .B(KEYINPUT100), .ZN(new_n278));
  INV_X1    g077(.A(new_n275), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n270), .B(new_n265), .C1(new_n279), .C2(new_n273), .ZN(new_n280));
  INV_X1    g079(.A(new_n230), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT99), .ZN(new_n284));
  XOR2_X1   g083(.A(G134gat), .B(G162gat), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT101), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n286), .A2(KEYINPUT101), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n277), .A2(new_n282), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n288), .B1(new_n277), .B2(new_n282), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G230gat), .ZN(new_n296));
  INV_X1    g095(.A(G233gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n263), .A2(new_n264), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n210), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n265), .A2(new_n209), .A3(new_n208), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT10), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n210), .A2(KEYINPUT10), .A3(new_n299), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n301), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n305), .B1(new_n306), .B2(new_n298), .ZN(new_n307));
  XNOR2_X1  g106(.A(G120gat), .B(G148gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(G176gat), .B(G204gat), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n308), .B(new_n309), .Z(new_n310));
  OR2_X1    g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n310), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n229), .A2(new_n295), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT96), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n317));
  XNOR2_X1  g116(.A(G113gat), .B(G120gat), .ZN(new_n318));
  OAI211_X1 g117(.A(KEYINPUT69), .B(G127gat), .C1(new_n318), .C2(KEYINPUT1), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  INV_X1    g119(.A(G113gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n321), .A2(G120gat), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(G113gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n320), .B(new_n214), .C1(new_n322), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G134gat), .ZN(new_n327));
  INV_X1    g126(.A(G134gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n319), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT27), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(G183gat), .ZN(new_n332));
  INV_X1    g131(.A(G183gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(KEYINPUT27), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT67), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(KEYINPUT27), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT67), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(G190gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n336), .A2(new_n337), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n340), .B1(new_n343), .B2(G190gat), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n342), .A2(KEYINPUT68), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT68), .B1(new_n342), .B2(new_n344), .ZN(new_n346));
  NOR2_X1   g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT26), .ZN(new_n348));
  NAND2_X1  g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT65), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT65), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(G169gat), .A3(G176gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n345), .A2(new_n346), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n347), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT64), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(KEYINPUT24), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT24), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(G183gat), .A3(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n353), .B(new_n361), .C1(new_n364), .C2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT66), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n350), .A2(new_n352), .A3(new_n372), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n361), .A2(new_n373), .A3(KEYINPUT25), .ZN(new_n374));
  INV_X1    g173(.A(new_n362), .ZN(new_n375));
  AOI22_X1  g174(.A1(KEYINPUT66), .A2(new_n353), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n370), .A2(new_n371), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n330), .B1(new_n357), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G227gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(new_n297), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT68), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n338), .B1(new_n336), .B2(new_n337), .ZN(new_n383));
  INV_X1    g182(.A(new_n341), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n344), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n381), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT68), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n354), .A2(new_n355), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n319), .A2(new_n325), .A3(new_n328), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n328), .B1(new_n319), .B2(new_n325), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n370), .A2(new_n371), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n376), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n390), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n380), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT70), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n378), .A2(KEYINPUT70), .A3(new_n380), .A4(new_n397), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT32), .ZN(new_n403));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n403), .B1(new_n407), .B2(KEYINPUT33), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n317), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n408), .ZN(new_n410));
  AOI211_X1 g209(.A(KEYINPUT71), .B(new_n410), .C1(new_n400), .C2(new_n401), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n400), .A2(new_n401), .B1(new_n403), .B2(KEYINPUT33), .ZN(new_n412));
  OAI22_X1  g211(.A1(new_n409), .A2(new_n411), .B1(new_n412), .B2(new_n406), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT34), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n378), .A2(new_n397), .ZN(new_n415));
  INV_X1    g214(.A(new_n380), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT72), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI211_X1 g218(.A(KEYINPUT72), .B(KEYINPUT34), .C1(new_n415), .C2(new_n416), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n413), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n403), .A2(KEYINPUT33), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n390), .A2(new_n393), .A3(new_n396), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n393), .B1(new_n390), .B2(new_n396), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT70), .B1(new_n427), .B2(new_n380), .ZN(new_n428));
  INV_X1    g227(.A(new_n401), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n407), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n421), .C1(new_n409), .C2(new_n411), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n423), .A2(KEYINPUT36), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT36), .B1(new_n423), .B2(new_n432), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G8gat), .B(G36gat), .Z(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT75), .ZN(new_n437));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  NAND2_X1  g238(.A1(new_n390), .A2(new_n396), .ZN(new_n440));
  INV_X1    g239(.A(G226gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(new_n297), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT29), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  OR2_X1    g245(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n447));
  NAND2_X1  g246(.A1(G211gat), .A2(G218gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G211gat), .ZN(new_n451));
  INV_X1    g250(.A(G218gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(KEYINPUT74), .A3(new_n448), .ZN(new_n454));
  XNOR2_X1  g253(.A(G197gat), .B(G204gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT74), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(new_n448), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n457), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n460), .A2(new_n450), .A3(new_n454), .A4(new_n455), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n444), .A2(new_n446), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n346), .A2(new_n356), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n377), .B1(new_n465), .B2(new_n388), .ZN(new_n466));
  OAI22_X1  g265(.A1(new_n466), .A2(KEYINPUT29), .B1(new_n441), .B2(new_n297), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n462), .B1(new_n467), .B2(new_n443), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n439), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n463), .B1(new_n444), .B2(new_n446), .ZN(new_n470));
  INV_X1    g269(.A(new_n439), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n462), .A3(new_n443), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(KEYINPUT30), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n475), .B(new_n439), .C1(new_n464), .C2(new_n468), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT78), .ZN(new_n481));
  AND2_X1   g280(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n483));
  INV_X1    g282(.A(G148gat), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G141gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(G148gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n481), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n487), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT77), .B(G141gat), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT78), .B(new_n489), .C1(new_n490), .C2(new_n484), .ZN(new_n491));
  AND2_X1   g290(.A1(G155gat), .A2(G162gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(G155gat), .A2(G162gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G155gat), .A2(G162gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT2), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT79), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(KEYINPUT79), .A3(KEYINPUT2), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n494), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n488), .A2(new_n491), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G141gat), .B(G148gat), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n502), .A2(KEYINPUT76), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n496), .B1(new_n502), .B2(KEYINPUT76), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n494), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n501), .A2(new_n505), .A3(KEYINPUT80), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(KEYINPUT3), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT3), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n393), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n480), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT83), .B(KEYINPUT5), .Z(new_n516));
  INV_X1    g315(.A(KEYINPUT82), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n506), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n505), .A3(KEYINPUT82), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n520));
  NAND4_X1  g319(.A1(new_n518), .A2(new_n330), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT4), .B1(new_n393), .B2(new_n506), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n515), .A2(new_n516), .A3(new_n523), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n501), .A2(KEYINPUT80), .A3(new_n505), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT80), .B1(new_n501), .B2(new_n505), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n525), .A2(new_n526), .A3(new_n511), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n479), .B1(new_n527), .B2(new_n513), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n393), .A2(new_n506), .A3(KEYINPUT4), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n518), .A2(new_n330), .A3(new_n519), .ZN(new_n530));
  INV_X1    g329(.A(new_n520), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n525), .A2(new_n526), .A3(new_n330), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n330), .A2(new_n505), .A3(new_n501), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n480), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n516), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n524), .B1(new_n533), .B2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G1gat), .B(G29gat), .Z(new_n541));
  XNOR2_X1  g340(.A(G57gat), .B(G85gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n510), .A2(new_n514), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n479), .B1(new_n523), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n508), .A2(new_n509), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n479), .B(new_n535), .C1(new_n550), .C2(new_n330), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT39), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT39), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n545), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT40), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n553), .A2(KEYINPUT40), .A3(new_n555), .A4(new_n545), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n478), .A2(new_n547), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G228gat), .A2(G233gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n512), .A2(new_n445), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n462), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n511), .B1(new_n462), .B2(KEYINPUT29), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n508), .A3(new_n509), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G22gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n518), .A2(new_n519), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n568), .A2(new_n564), .B1(new_n462), .B2(new_n562), .ZN(new_n569));
  INV_X1    g368(.A(new_n561), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n566), .B(new_n567), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT86), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n501), .A2(KEYINPUT82), .A3(new_n505), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT82), .B1(new_n501), .B2(new_n505), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n564), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n562), .A2(new_n462), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n578), .A2(new_n561), .B1(new_n565), .B2(new_n563), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(KEYINPUT86), .A3(new_n567), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G22gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n573), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G78gat), .B(G106gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT31), .B(G50gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT85), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT87), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n579), .A2(KEYINPUT87), .A3(new_n567), .ZN(new_n591));
  INV_X1    g390(.A(new_n586), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n582), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT88), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT6), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n530), .A2(new_n531), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n515), .B1(new_n597), .B2(new_n529), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n535), .B1(new_n550), .B2(new_n330), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n516), .B1(new_n599), .B2(new_n480), .ZN(new_n600));
  AOI211_X1 g399(.A(new_n480), .B(new_n538), .C1(new_n510), .C2(new_n514), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n598), .A2(new_n600), .B1(new_n523), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n596), .B1(new_n602), .B2(new_n545), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n545), .B(new_n524), .C1(new_n533), .C2(new_n539), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n595), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n540), .A2(KEYINPUT6), .A3(new_n546), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n547), .A2(new_n604), .A3(KEYINPUT88), .A4(new_n596), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT37), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n470), .A2(new_n610), .A3(new_n472), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n470), .B2(new_n472), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n471), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT38), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT38), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n616), .B(new_n471), .C1(new_n612), .C2(new_n613), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n617), .A3(new_n469), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n560), .B(new_n594), .C1(new_n609), .C2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n547), .A2(new_n604), .A3(new_n596), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n607), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n477), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n590), .A2(new_n592), .A3(new_n582), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n623), .A2(new_n591), .B1(new_n583), .B2(new_n587), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n435), .A2(new_n619), .A3(new_n625), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n620), .A2(new_n607), .B1(new_n476), .B2(new_n474), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n410), .B1(new_n400), .B2(new_n401), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(new_n317), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n421), .B1(new_n629), .B2(new_n431), .ZN(new_n630));
  INV_X1    g429(.A(new_n432), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n594), .B(new_n627), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT35), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n624), .B1(new_n423), .B2(new_n432), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT35), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n609), .A4(new_n477), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n626), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G113gat), .B(G141gat), .ZN(new_n639));
  INV_X1    g438(.A(G197gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT11), .B(G169gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n221), .B(G8gat), .Z(new_n645));
  AND2_X1   g444(.A1(new_n645), .A2(new_n270), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n279), .B2(new_n273), .ZN(new_n647));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n255), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(KEYINPUT92), .A3(new_n222), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT92), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n645), .B2(new_n255), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n647), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT18), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n649), .B2(new_n222), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n645), .A2(KEYINPUT94), .A3(new_n255), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n648), .B(KEYINPUT13), .Z(new_n660));
  AOI22_X1  g459(.A1(new_n654), .A2(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n647), .A2(KEYINPUT18), .A3(new_n648), .A4(new_n653), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n662), .A2(KEYINPUT93), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(KEYINPUT93), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n644), .B(new_n661), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n662), .B(KEYINPUT93), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n668), .A2(KEYINPUT95), .A3(new_n644), .A4(new_n661), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n661), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n644), .B(KEYINPUT89), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n667), .A2(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n316), .B1(new_n638), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n558), .A2(new_n547), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n474), .A2(new_n559), .A3(new_n476), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n594), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n615), .A2(new_n617), .A3(new_n469), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n423), .A2(new_n432), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT36), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n423), .A2(KEYINPUT36), .A3(new_n432), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n625), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n637), .B1(new_n679), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n672), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(KEYINPUT96), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n315), .B1(new_n673), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n621), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n687), .ZN(new_n692));
  INV_X1    g491(.A(new_n315), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G8gat), .B1(new_n694), .B2(new_n477), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  NAND3_X1  g496(.A1(new_n688), .A2(new_n478), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n698), .A2(new_n699), .A3(new_n696), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n698), .B2(new_n696), .ZN(new_n701));
  OAI221_X1 g500(.A(new_n695), .B1(new_n696), .B2(new_n698), .C1(new_n700), .C2(new_n701), .ZN(G1325gat));
  OAI21_X1  g501(.A(G15gat), .B1(new_n694), .B2(new_n435), .ZN(new_n703));
  INV_X1    g502(.A(new_n680), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n704), .A2(G15gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n694), .B2(new_n705), .ZN(G1326gat));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n624), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT103), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  NOR2_X1   g509(.A1(new_n229), .A2(new_n313), .ZN(new_n711));
  INV_X1    g510(.A(new_n295), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n673), .B2(new_n687), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G29gat), .A3(new_n621), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(KEYINPUT45), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(KEYINPUT45), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT104), .B1(new_n684), .B2(new_n679), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n435), .A2(new_n619), .A3(new_n720), .A4(new_n625), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n633), .A2(new_n722), .A3(new_n636), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n633), .B2(new_n636), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n719), .B(new_n721), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT106), .B1(new_n293), .B2(new_n294), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n277), .A2(new_n282), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n728), .B(new_n292), .C1(new_n729), .C2(new_n288), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n725), .A2(new_n726), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n726), .B1(new_n685), .B2(new_n712), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n735), .A2(new_n686), .A3(new_n711), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(new_n689), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n717), .B(new_n718), .C1(new_n233), .C2(new_n737), .ZN(G1328gat));
  NOR3_X1   g537(.A1(new_n715), .A2(G36gat), .A3(new_n477), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n736), .A2(new_n478), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n741), .B(new_n742), .C1(new_n237), .C2(new_n743), .ZN(G1329gat));
  NOR2_X1   g543(.A1(new_n704), .A2(G43gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n714), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT47), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n435), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n736), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n746), .B(new_n749), .C1(new_n751), .C2(new_n240), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n240), .B1(new_n736), .B2(new_n750), .ZN(new_n753));
  INV_X1    g552(.A(new_n746), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n748), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(G1330gat));
  NAND3_X1  g555(.A1(new_n736), .A2(G50gat), .A3(new_n624), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n247), .B1(new_n715), .B2(new_n594), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT48), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n757), .A2(new_n761), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1331gat));
  INV_X1    g562(.A(new_n229), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n712), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n725), .A2(new_n672), .A3(new_n765), .A4(new_n313), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n621), .B(KEYINPUT108), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g570(.A1(new_n767), .A2(KEYINPUT109), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  AND2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n775), .B(new_n478), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n775), .A2(new_n478), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(new_n776), .ZN(G1333gat));
  NAND4_X1  g579(.A1(new_n772), .A2(G71gat), .A3(new_n750), .A4(new_n774), .ZN(new_n781));
  INV_X1    g580(.A(G71gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n766), .B2(new_n704), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g584(.A1(new_n775), .A2(new_n624), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT110), .B(G78gat), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n786), .B(new_n788), .ZN(G1335gat));
  NOR3_X1   g588(.A1(new_n686), .A2(new_n229), .A3(new_n295), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n725), .A2(KEYINPUT51), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT111), .ZN(new_n792));
  INV_X1    g591(.A(new_n790), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n719), .A2(new_n721), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n637), .A2(KEYINPUT105), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n633), .A2(new_n722), .A3(new_n636), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n793), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT112), .B1(new_n798), .B2(KEYINPUT51), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n725), .A2(new_n790), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n792), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n805), .A2(new_n260), .A3(new_n689), .A4(new_n313), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n686), .A2(new_n229), .A3(new_n314), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n735), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(new_n689), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n806), .B1(new_n260), .B2(new_n809), .ZN(G1336gat));
  NAND2_X1  g609(.A1(new_n731), .A2(new_n726), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n794), .B2(new_n797), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n478), .B(new_n807), .C1(new_n812), .C2(new_n733), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G92gat), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n800), .B(KEYINPUT51), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n478), .A2(new_n261), .A3(new_n313), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT113), .Z(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n817), .B1(new_n792), .B2(new_n804), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n820), .A2(KEYINPUT114), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824));
  INV_X1    g623(.A(new_n817), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n801), .B1(new_n800), .B2(new_n802), .ZN(new_n826));
  AOI211_X1 g625(.A(KEYINPUT112), .B(KEYINPUT51), .C1(new_n725), .C2(new_n790), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n798), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n791), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n825), .B1(new_n828), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(new_n813), .B2(G92gat), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n824), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n819), .B1(new_n823), .B2(new_n835), .ZN(G1337gat));
  NOR3_X1   g635(.A1(new_n704), .A2(G99gat), .A3(new_n314), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n805), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n808), .A2(new_n750), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G99gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(G1338gat));
  NAND3_X1  g640(.A1(new_n735), .A2(new_n624), .A3(new_n807), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G106gat), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n594), .A2(new_n314), .A3(G106gat), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT115), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n815), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n805), .A2(new_n844), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(G1339gat));
  NOR2_X1   g650(.A1(new_n315), .A2(new_n686), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n667), .A2(new_n669), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n647), .A2(new_n653), .ZN(new_n854));
  OAI22_X1  g653(.A1(new_n854), .A2(new_n648), .B1(new_n660), .B2(new_n659), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n643), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858));
  XOR2_X1   g657(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI211_X1 g659(.A(new_n298), .B(new_n860), .C1(new_n303), .C2(new_n304), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n858), .B1(new_n861), .B2(new_n310), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n305), .A2(new_n859), .ZN(new_n863));
  INV_X1    g662(.A(new_n310), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(KEYINPUT117), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n305), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n303), .A2(new_n304), .A3(new_n298), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(KEYINPUT54), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n866), .A2(KEYINPUT55), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n312), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT55), .B1(new_n866), .B2(new_n869), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n857), .A2(new_n314), .B1(new_n672), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n731), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n853), .A2(new_n731), .A3(new_n856), .A4(new_n873), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT118), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n667), .A2(new_n669), .B1(new_n643), .B2(new_n855), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n731), .A4(new_n873), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n852), .B1(new_n884), .B2(new_n764), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n768), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n477), .A3(new_n634), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n321), .A3(new_n686), .ZN(new_n889));
  INV_X1    g688(.A(new_n634), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n621), .A2(new_n478), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G113gat), .B1(new_n893), .B2(new_n672), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT119), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n889), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1340gat));
  NOR3_X1   g698(.A1(new_n893), .A2(new_n323), .A3(new_n314), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n888), .A2(new_n313), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n323), .ZN(G1341gat));
  OAI21_X1  g701(.A(G127gat), .B1(new_n893), .B2(new_n764), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n229), .A2(new_n214), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n887), .B2(new_n904), .ZN(G1342gat));
  NAND2_X1  g704(.A1(new_n712), .A2(new_n477), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT120), .ZN(new_n907));
  XNOR2_X1  g706(.A(KEYINPUT69), .B(G134gat), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n907), .A2(new_n890), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n886), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n886), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT122), .B1(new_n914), .B2(KEYINPUT56), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n911), .A2(new_n916), .A3(new_n917), .A4(new_n913), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n891), .A2(new_n712), .A3(new_n892), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n914), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1343gat));
  NAND2_X1  g721(.A1(new_n435), .A2(new_n892), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n852), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n876), .A2(new_n875), .B1(new_n879), .B2(new_n882), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n229), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT57), .B1(new_n927), .B2(new_n624), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n624), .A2(KEYINPUT57), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n875), .A2(new_n295), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n883), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n764), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n930), .B1(new_n933), .B2(new_n925), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n686), .B(new_n924), .C1(new_n928), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT123), .B1(new_n935), .B2(new_n490), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n750), .A2(new_n594), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n927), .A2(new_n769), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n686), .A2(new_n486), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n938), .A2(new_n478), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n935), .B2(new_n490), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n936), .A2(new_n941), .A3(KEYINPUT58), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT58), .ZN(new_n943));
  AOI221_X4 g742(.A(new_n940), .B1(KEYINPUT123), .B2(new_n943), .C1(new_n490), .C2(new_n935), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n942), .A2(new_n944), .ZN(G1344gat));
  NOR4_X1   g744(.A1(new_n938), .A2(G148gat), .A3(new_n478), .A4(new_n314), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT124), .Z(new_n947));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n857), .A2(new_n295), .A3(new_n874), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n949), .B1(new_n295), .B2(new_n875), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n925), .B1(new_n950), .B2(new_n229), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(new_n624), .ZN(new_n952));
  OAI22_X1  g751(.A1(new_n952), .A2(KEYINPUT57), .B1(new_n885), .B2(new_n930), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n313), .A3(new_n924), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n948), .B1(new_n954), .B2(G148gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n924), .B1(new_n928), .B2(new_n934), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(new_n314), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n957), .A2(KEYINPUT59), .A3(new_n484), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n947), .B1(new_n955), .B2(new_n958), .ZN(G1345gat));
  OAI21_X1  g758(.A(G155gat), .B1(new_n956), .B2(new_n764), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n886), .A2(new_n477), .A3(new_n937), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n229), .A2(new_n226), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(G1346gat));
  OAI21_X1  g762(.A(G162gat), .B1(new_n956), .B2(new_n876), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n907), .A2(G162gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n938), .B2(new_n965), .ZN(G1347gat));
  NOR2_X1   g765(.A1(new_n769), .A2(new_n477), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n891), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(G169gat), .B1(new_n968), .B2(new_n672), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n927), .A2(new_n621), .A3(new_n478), .A4(new_n634), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n970), .A2(G169gat), .A3(new_n672), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT125), .Z(G1348gat));
  OAI21_X1  g772(.A(G176gat), .B1(new_n968), .B2(new_n314), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n314), .A2(G176gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n970), .B2(new_n975), .ZN(G1349gat));
  NAND3_X1  g775(.A1(new_n229), .A2(new_n335), .A3(new_n339), .ZN(new_n977));
  OR3_X1    g776(.A1(new_n970), .A2(KEYINPUT126), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(KEYINPUT126), .B1(new_n970), .B2(new_n977), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(G183gat), .B1(new_n968), .B2(new_n764), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(KEYINPUT60), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT60), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n980), .A2(new_n984), .A3(new_n981), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(G1350gat));
  NAND3_X1  g785(.A1(new_n891), .A2(new_n712), .A3(new_n967), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n987), .A2(new_n988), .A3(G190gat), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n988), .B1(new_n987), .B2(G190gat), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n876), .A2(G190gat), .ZN(new_n992));
  OAI22_X1  g791(.A1(new_n990), .A2(new_n991), .B1(new_n970), .B2(new_n992), .ZN(G1351gat));
  NOR3_X1   g792(.A1(new_n769), .A2(new_n750), .A3(new_n477), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n953), .A2(new_n994), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n995), .A2(new_n640), .A3(new_n672), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n885), .A2(new_n689), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n750), .A2(new_n594), .A3(new_n477), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g799(.A(G197gat), .B1(new_n1000), .B2(new_n686), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n996), .A2(new_n1001), .ZN(G1352gat));
  OR3_X1    g801(.A1(new_n999), .A2(G204gat), .A3(new_n314), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  OAI21_X1  g803(.A(G204gat), .B1(new_n995), .B2(new_n314), .ZN(new_n1005));
  NOR3_X1   g804(.A1(new_n1003), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n1007));
  NOR3_X1   g806(.A1(new_n999), .A2(G204gat), .A3(new_n314), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g809(.A(new_n1004), .B(new_n1005), .C1(new_n1006), .C2(new_n1010), .ZN(G1353gat));
  NAND3_X1  g810(.A1(new_n1000), .A2(new_n451), .A3(new_n229), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n953), .A2(new_n229), .A3(new_n994), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n1013), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1014));
  AOI21_X1  g813(.A(KEYINPUT63), .B1(new_n1013), .B2(G211gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(G1354gat));
  OAI21_X1  g815(.A(G218gat), .B1(new_n995), .B2(new_n295), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n1000), .A2(new_n452), .A3(new_n731), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1017), .A2(new_n1018), .ZN(G1355gat));
endmodule


