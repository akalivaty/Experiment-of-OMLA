//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT0), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT0), .B(G128), .Z(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(new_n189), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G125), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  AND4_X1   g014(.A1(new_n196), .A2(new_n198), .A3(new_n200), .A4(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(KEYINPUT1), .A3(G146), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(G128), .B1(new_n198), .B2(new_n200), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n195), .B1(new_n205), .B2(G125), .ZN(new_n206));
  INV_X1    g020(.A(G953), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G224), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n206), .B(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT67), .B1(new_n210), .B2(G116), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n212));
  INV_X1    g026(.A(G116), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(G116), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT2), .B(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n218), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n215), .A3(new_n216), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT3), .B1(new_n223), .B2(G107), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  INV_X1    g039(.A(G107), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G104), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(G107), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G101), .ZN(new_n230));
  INV_X1    g044(.A(G101), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n224), .A2(new_n227), .A3(new_n231), .A4(new_n228), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(KEYINPUT4), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n229), .A2(new_n234), .A3(G101), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n222), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n215), .A2(KEYINPUT5), .A3(new_n216), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n237), .B(G113), .C1(KEYINPUT5), .C2(new_n216), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n226), .A2(G104), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n223), .A2(G107), .ZN(new_n240));
  OAI21_X1  g054(.A(G101), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n232), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n238), .A2(new_n221), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n236), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(G110), .B(G122), .Z(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OR2_X1    g060(.A1(new_n246), .A2(KEYINPUT6), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n248));
  INV_X1    g062(.A(new_n245), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n236), .B2(new_n243), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT87), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n236), .A2(new_n243), .A3(new_n249), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n253), .A2(KEYINPUT6), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n248), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n246), .A2(new_n251), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n250), .A2(KEYINPUT87), .ZN(new_n257));
  AND4_X1   g071(.A1(new_n248), .A2(new_n256), .A3(new_n254), .A4(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n209), .B(new_n247), .C1(new_n255), .C2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G902), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT7), .B1(new_n207), .B2(G224), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n209), .B(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n238), .A2(new_n221), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(new_n242), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n245), .B(KEYINPUT8), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n262), .B(new_n253), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n259), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(G210), .B1(G237), .B2(G902), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n259), .A2(new_n266), .A3(new_n260), .A4(new_n268), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n188), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G113), .B(G122), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(new_n223), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT78), .ZN(new_n276));
  INV_X1    g090(.A(G125), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT77), .A3(G140), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n280));
  XNOR2_X1  g094(.A(G125), .B(G140), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT16), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G140), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n285), .A3(G125), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(G125), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n277), .A2(G140), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n278), .B1(new_n289), .B2(KEYINPUT77), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT78), .A3(KEYINPUT16), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n284), .A2(G146), .A3(new_n286), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT91), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT19), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n281), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n197), .B(new_n295), .C1(new_n290), .C2(new_n294), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n292), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n293), .B1(new_n292), .B2(new_n296), .ZN(new_n298));
  INV_X1    g112(.A(G237), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n207), .A3(G214), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n300), .B(G143), .ZN(new_n301));
  INV_X1    g115(.A(G131), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n300), .B(new_n199), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G131), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT90), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT90), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n297), .A2(new_n298), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n304), .A2(KEYINPUT89), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT18), .A2(G131), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n289), .A2(G146), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT79), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n282), .A2(G146), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n275), .B1(new_n311), .B2(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n314), .A2(new_n318), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT17), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n305), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n305), .A2(new_n303), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(new_n322), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n284), .A2(new_n286), .A3(new_n291), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n197), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(new_n292), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n321), .A2(new_n328), .A3(new_n274), .ZN(new_n329));
  AOI21_X1  g143(.A(G475), .B1(new_n320), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT20), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n260), .ZN(new_n332));
  INV_X1    g146(.A(G475), .ZN(new_n333));
  INV_X1    g147(.A(new_n298), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n307), .A2(new_n309), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n292), .A2(new_n293), .A3(new_n296), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n274), .B1(new_n337), .B2(new_n321), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n321), .A2(new_n328), .A3(new_n274), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n333), .B(new_n260), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT20), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n274), .B1(new_n321), .B2(new_n328), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n260), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G475), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(G234), .A2(G237), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(G952), .A3(new_n207), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT21), .B(G898), .Z(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(G902), .A3(G953), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G122), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G116), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT92), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n353), .A2(G116), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n226), .A3(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n358), .A2(KEYINPUT93), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT14), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n355), .B1(new_n360), .B2(new_n356), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n213), .A3(G122), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n362), .B(KEYINPUT94), .Z(new_n363));
  OAI21_X1  g177(.A(G107), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G128), .B(G143), .ZN(new_n365));
  INV_X1    g179(.A(G134), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n358), .A2(KEYINPUT93), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n359), .A2(new_n364), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(KEYINPUT13), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n199), .A2(G128), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n370), .B(G134), .C1(KEYINPUT13), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n365), .A2(new_n366), .ZN(new_n373));
  INV_X1    g187(.A(new_n358), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n226), .B1(new_n355), .B2(new_n357), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n372), .B(new_n373), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT9), .B(G234), .Z(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(G217), .A3(new_n207), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n369), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n369), .B2(new_n376), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n260), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND2_X1   g196(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n383));
  NOR2_X1   g197(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n384));
  OAI21_X1  g198(.A(G478), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n382), .B(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n346), .A2(new_n352), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G469), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n233), .A2(new_n194), .A3(new_n235), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n198), .A2(new_n200), .A3(new_n196), .A4(G128), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n391), .B(new_n202), .C1(G128), .C2(new_n189), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n242), .A2(new_n392), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n393), .A2(KEYINPUT82), .A3(KEYINPUT10), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT10), .B1(new_n393), .B2(KEYINPUT82), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT11), .ZN(new_n397));
  OAI211_X1 g211(.A(KEYINPUT64), .B(new_n397), .C1(new_n366), .C2(G137), .ZN(new_n398));
  INV_X1    g212(.A(G137), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT64), .ZN(new_n400));
  OAI211_X1 g214(.A(G134), .B(new_n399), .C1(new_n400), .C2(KEYINPUT11), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(KEYINPUT11), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT65), .B1(new_n399), .B2(G134), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT65), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n366), .A3(G137), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G131), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n397), .A2(KEYINPUT64), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n366), .A2(G137), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n397), .A2(KEYINPUT64), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n404), .A2(new_n406), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n412), .A2(new_n302), .A3(new_n413), .A4(new_n398), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT68), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n408), .A2(KEYINPUT68), .A3(new_n414), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT83), .B1(new_n396), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n390), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n232), .A2(new_n241), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT82), .B1(new_n205), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT10), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n393), .A2(KEYINPUT82), .A3(KEYINPUT10), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n422), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n419), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n421), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(G110), .B(G140), .Z(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT81), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n207), .A2(G227), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n396), .A2(new_n420), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n431), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n205), .A2(new_n423), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n393), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n415), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT12), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n439), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n419), .A2(new_n443), .A3(KEYINPUT12), .ZN(new_n444));
  AOI211_X1 g258(.A(new_n442), .B(new_n444), .C1(new_n421), .C2(new_n430), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n437), .B1(new_n445), .B2(new_n435), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n389), .B1(new_n446), .B2(new_n260), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n396), .A2(new_n420), .A3(KEYINPUT83), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n429), .B1(new_n428), .B2(new_n419), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n436), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n435), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n444), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n431), .A2(new_n453), .A3(new_n441), .A4(new_n435), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT84), .B(G469), .Z(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n260), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT85), .ZN(new_n459));
  AOI21_X1  g273(.A(G902), .B1(new_n452), .B2(new_n454), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n457), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n447), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n464));
  INV_X1    g278(.A(G221), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n377), .B2(new_n260), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n447), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n460), .A2(new_n461), .A3(new_n457), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n461), .B1(new_n460), .B2(new_n457), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n466), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT86), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n272), .B(new_n388), .C1(new_n467), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT96), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT22), .B(G137), .ZN(new_n477));
  INV_X1    g291(.A(G234), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n465), .A2(new_n478), .A3(G953), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n477), .B(new_n479), .Z(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G110), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n191), .A2(G119), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT23), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n210), .A2(G128), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT23), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT75), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT75), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT23), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT76), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n485), .A2(new_n487), .A3(new_n489), .A4(KEYINPUT76), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI211_X1 g308(.A(new_n482), .B(new_n484), .C1(new_n494), .C2(new_n483), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT24), .B(G110), .Z(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n483), .A3(new_n485), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI211_X1 g312(.A(new_n495), .B(new_n498), .C1(new_n327), .C2(new_n292), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n496), .B1(new_n483), .B2(new_n485), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n483), .ZN(new_n501));
  INV_X1    g315(.A(new_n484), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n500), .B1(new_n503), .B2(new_n482), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n292), .A2(new_n316), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n481), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n506), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n327), .A2(new_n292), .ZN(new_n509));
  INV_X1    g323(.A(new_n495), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n497), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n511), .A3(new_n480), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(new_n512), .A3(new_n260), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT25), .ZN(new_n514));
  OAI21_X1  g328(.A(G217), .B1(new_n478), .B2(G902), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT74), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n507), .A2(new_n512), .A3(new_n517), .A4(new_n260), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT80), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT80), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n514), .A2(new_n521), .A3(new_n516), .A4(new_n518), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n513), .A2(new_n516), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n417), .A2(new_n418), .A3(new_n194), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n366), .A2(G137), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n399), .A2(G134), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n302), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT66), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n414), .A3(new_n392), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(KEYINPUT30), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n415), .A2(new_n194), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n530), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(new_n222), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n222), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n525), .A2(new_n537), .A3(new_n530), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n299), .A2(new_n207), .A3(G210), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(new_n231), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n541), .B(new_n542), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT69), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n525), .A2(KEYINPUT28), .A3(new_n537), .A4(new_n530), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n533), .A2(new_n222), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n548), .A2(new_n543), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT29), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT69), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n539), .A2(new_n554), .A3(new_n544), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n546), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT70), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n548), .A2(KEYINPUT71), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n525), .A2(new_n530), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n222), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n548), .A2(new_n560), .A3(KEYINPUT71), .A4(new_n549), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n544), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(G902), .B1(new_n562), .B2(KEYINPUT29), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT70), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n546), .A2(new_n553), .A3(new_n564), .A4(new_n555), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n557), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G472), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT72), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT72), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n569), .A3(G472), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n536), .A2(new_n543), .A3(new_n538), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n572), .A2(KEYINPUT31), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n544), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(KEYINPUT31), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G472), .A2(G902), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT73), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n578), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT32), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT73), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n577), .A2(new_n584), .A3(KEYINPUT32), .A4(new_n578), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n580), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n524), .B1(new_n571), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n270), .A2(new_n271), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n187), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n464), .B1(new_n463), .B2(new_n466), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n471), .A2(KEYINPUT86), .A3(new_n472), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(KEYINPUT96), .A3(new_n388), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n476), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  NAND2_X1  g409(.A1(new_n577), .A2(new_n260), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(new_n581), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n590), .B2(new_n591), .ZN(new_n600));
  INV_X1    g414(.A(new_n524), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n188), .B(new_n352), .C1(new_n270), .C2(new_n271), .ZN(new_n603));
  INV_X1    g417(.A(G478), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n382), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(new_n607));
  OR3_X1    g421(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT33), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT33), .B1(new_n380), .B2(new_n381), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(G478), .A3(new_n260), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n346), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n603), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n602), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT34), .B(G104), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  NAND2_X1  g432(.A1(new_n387), .A2(new_n345), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT98), .B1(new_n340), .B2(KEYINPUT20), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n330), .A2(new_n621), .A3(new_n331), .A4(new_n260), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n622), .A3(new_n341), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n620), .A2(new_n622), .A3(KEYINPUT99), .A4(new_n341), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n619), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n603), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n600), .A2(new_n601), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NAND2_X1  g445(.A1(new_n508), .A2(new_n511), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n481), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n516), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n260), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n520), .A2(new_n522), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n476), .A2(new_n593), .A3(new_n598), .A4(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT37), .B(G110), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  AND3_X1   g456(.A1(new_n566), .A2(new_n569), .A3(G472), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n569), .B1(new_n566), .B2(G472), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n586), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n348), .B(KEYINPUT101), .Z(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(G900), .B2(new_n350), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT102), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n627), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n592), .A2(new_n645), .A3(new_n639), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  NAND2_X1  g468(.A1(new_n346), .A2(new_n387), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n637), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n588), .B(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n560), .A2(new_n538), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n544), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n661), .A2(new_n572), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n662), .B2(G902), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n586), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n659), .A2(new_n665), .A3(new_n188), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n590), .A2(new_n591), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n649), .B(KEYINPUT39), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n656), .B(new_n666), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  NAND3_X1  g489(.A1(new_n346), .A2(new_n612), .A3(new_n650), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n592), .A2(new_n645), .A3(new_n639), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT104), .B(G146), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G48));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n589), .A2(new_n613), .A3(new_n352), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n459), .A2(new_n462), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n460), .A2(new_n389), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n466), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n587), .A2(new_n681), .A3(new_n682), .A4(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n645), .A2(new_n682), .A3(new_n601), .A4(new_n686), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT105), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT106), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n690), .B(new_n692), .ZN(G15));
  NAND4_X1  g507(.A1(new_n645), .A2(new_n628), .A3(new_n601), .A4(new_n686), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  AND4_X1   g509(.A1(new_n272), .A2(new_n472), .A3(new_n683), .A4(new_n684), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n645), .A2(new_n388), .A3(new_n639), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  XOR2_X1   g512(.A(new_n524), .B(KEYINPUT108), .Z(new_n699));
  NOR3_X1   g513(.A1(new_n589), .A2(new_n655), .A3(new_n352), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n558), .A2(new_n701), .A3(new_n561), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n544), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n701), .B1(new_n558), .B2(new_n561), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n576), .B(new_n573), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n578), .A2(new_n705), .B1(new_n596), .B2(G472), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n699), .A2(new_n700), .A3(new_n686), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  AND2_X1   g522(.A1(new_n706), .A2(new_n637), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n696), .A2(new_n677), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  OAI21_X1  g525(.A(KEYINPUT109), .B1(new_n445), .B2(new_n435), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n431), .A2(new_n453), .A3(new_n441), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n451), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n712), .A2(new_n437), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n260), .ZN(new_n717));
  AOI22_X1  g531(.A1(G469), .A2(new_n717), .B1(new_n459), .B2(new_n462), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n466), .A2(new_n188), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n718), .A2(new_n588), .A3(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n645), .A2(new_n721), .A3(new_n601), .A4(new_n677), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n571), .A2(new_n583), .A3(new_n579), .ZN(new_n725));
  NOR4_X1   g539(.A1(new_n718), .A2(new_n676), .A3(new_n588), .A4(new_n720), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(KEYINPUT42), .A3(new_n699), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  NAND2_X1  g543(.A1(new_n651), .A2(KEYINPUT110), .ZN(new_n730));
  AND4_X1   g544(.A1(new_n645), .A2(new_n730), .A3(new_n601), .A4(new_n721), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n651), .A2(KEYINPUT110), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  NAND3_X1  g548(.A1(new_n612), .A2(new_n342), .A3(new_n345), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT43), .Z(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n599), .A3(new_n637), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(KEYINPUT44), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n446), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(G469), .C1(new_n716), .C2(new_n740), .ZN(new_n742));
  NAND2_X1  g556(.A1(G469), .A2(G902), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(KEYINPUT111), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(KEYINPUT111), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n683), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n472), .A3(new_n669), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n739), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n270), .A2(new_n187), .A3(new_n271), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n738), .B2(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G137), .ZN(G39));
  NAND2_X1  g572(.A1(new_n749), .A2(new_n472), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n749), .A2(KEYINPUT47), .A3(new_n472), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n676), .B(new_n755), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n571), .A2(new_n586), .A3(new_n524), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  INV_X1    g581(.A(G952), .ZN(new_n768));
  INV_X1    g582(.A(new_n755), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n665), .A2(new_n686), .A3(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n770), .A2(new_n524), .A3(new_n348), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n768), .B(G953), .C1(new_n771), .C2(new_n614), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n725), .A2(new_n699), .ZN(new_n773));
  AND4_X1   g587(.A1(new_n646), .A2(new_n736), .A3(new_n686), .A4(new_n769), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n772), .B1(KEYINPUT48), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(KEYINPUT48), .B2(new_n775), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n646), .A2(new_n736), .A3(new_n699), .A4(new_n706), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n188), .A3(new_n659), .A4(new_n686), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(KEYINPUT118), .B2(new_n780), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n781), .A2(KEYINPUT118), .A3(new_n780), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n346), .A2(new_n612), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n771), .A2(new_n783), .B1(new_n709), .B2(new_n774), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(KEYINPUT118), .B2(new_n780), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n761), .A2(new_n762), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n685), .A2(new_n472), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n769), .B(new_n778), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n777), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n782), .A2(KEYINPUT119), .A3(new_n785), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT119), .B1(new_n782), .B2(new_n785), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n784), .B(new_n789), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n694), .A2(new_n697), .A3(new_n707), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n690), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n797), .B1(new_n690), .B2(new_n798), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n682), .A2(KEYINPUT114), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n346), .A2(new_n386), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n603), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n615), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n601), .A3(new_n600), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n594), .A2(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n724), .A2(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n755), .A2(new_n649), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n645), .A2(new_n812), .A3(new_n639), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n625), .A2(new_n626), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n345), .A3(new_n386), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n667), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n811), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n637), .B(KEYINPUT100), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n571), .B2(new_n586), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n815), .B1(new_n590), .B2(new_n591), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(KEYINPUT115), .A3(new_n821), .A4(new_n812), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n818), .A2(new_n822), .B1(new_n709), .B2(new_n726), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n809), .A2(new_n640), .A3(new_n810), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT116), .B1(new_n801), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n690), .A2(new_n798), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT113), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n690), .A2(new_n798), .A3(new_n797), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n818), .A2(new_n822), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n726), .A2(new_n709), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n733), .A3(new_n728), .A4(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n640), .A2(new_n594), .A3(new_n808), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n829), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n589), .A2(new_n655), .A3(new_n649), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n718), .A2(new_n637), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n664), .A3(new_n472), .A4(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n653), .A2(new_n678), .A3(new_n710), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n841), .A2(new_n842), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n837), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n653), .A2(new_n678), .A3(new_n710), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(KEYINPUT52), .A3(new_n840), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(KEYINPUT117), .A3(new_n843), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n825), .A2(new_n836), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n825), .A2(new_n836), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n844), .B2(new_n845), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n852), .B(KEYINPUT54), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n778), .A2(new_n696), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n844), .A2(new_n845), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n858), .A2(new_n824), .A3(new_n854), .A4(new_n826), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n851), .B2(new_n854), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n796), .A2(new_n856), .A3(new_n857), .A4(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(G952), .B2(G953), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n685), .B(KEYINPUT49), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n865), .A2(new_n664), .A3(new_n735), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n659), .A3(new_n699), .A4(new_n719), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n867), .ZN(G75));
  NAND2_X1  g682(.A1(new_n851), .A2(new_n854), .ZN(new_n869));
  INV_X1    g683(.A(new_n859), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(G210), .A3(G902), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n247), .B1(new_n255), .B2(new_n258), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n209), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT55), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n768), .A2(G953), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT121), .Z(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n860), .A2(new_n260), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT56), .B1(new_n882), .B2(G210), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n873), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n877), .B1(new_n883), .B2(new_n873), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(G51));
  INV_X1    g700(.A(new_n880), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n743), .B(KEYINPUT57), .Z(new_n888));
  INV_X1    g702(.A(new_n862), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n860), .A2(new_n861), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n455), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n860), .A2(new_n260), .A3(new_n742), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(G54));
  NAND3_X1  g708(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n320), .A2(new_n329), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n887), .B1(new_n897), .B2(new_n898), .ZN(G60));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT59), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n610), .B(new_n902), .C1(new_n889), .C2(new_n890), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n856), .B2(new_n862), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n903), .B(new_n880), .C1(new_n610), .C2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(G63));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT60), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n871), .A2(new_n634), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT61), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n507), .A2(new_n512), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n860), .B2(new_n908), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n880), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n912), .B(new_n915), .ZN(G66));
  AOI21_X1  g730(.A(new_n207), .B1(new_n349), .B2(G224), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n801), .A2(new_n833), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n919), .B2(new_n207), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n875), .B1(G898), .B2(new_n207), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n920), .B(new_n921), .Z(G69));
  INV_X1    g736(.A(G900), .ZN(new_n923));
  OAI21_X1  g737(.A(G953), .B1(new_n923), .B2(G227), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n754), .A2(new_n756), .B1(new_n763), .B2(new_n765), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n752), .A2(new_n753), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n589), .A2(new_n655), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n927), .A3(new_n773), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n810), .B(KEYINPUT124), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n925), .A2(new_n847), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n924), .B1(new_n930), .B2(G953), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n531), .A2(new_n535), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n295), .B1(new_n290), .B2(new_n294), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n587), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n671), .B(new_n769), .C1(new_n614), .C2(new_n803), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n757), .B(new_n207), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n674), .A2(new_n847), .ZN(new_n940));
  NAND2_X1  g754(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g756(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n943));
  OAI211_X1 g757(.A(new_n766), .B(new_n942), .C1(new_n940), .C2(new_n943), .ZN(new_n944));
  OAI22_X1  g758(.A1(new_n939), .A2(new_n944), .B1(new_n923), .B2(new_n924), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n936), .B1(new_n935), .B2(new_n945), .ZN(G72));
  XNOR2_X1  g760(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n947));
  NAND2_X1  g761(.A1(G472), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n930), .B2(new_n919), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n539), .B(KEYINPUT126), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n544), .A3(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n757), .B(new_n918), .C1(new_n937), .C2(new_n938), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n949), .B1(new_n953), .B2(new_n944), .ZN(new_n954));
  INV_X1    g768(.A(new_n951), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n543), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n952), .A2(new_n956), .A3(new_n880), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n852), .B1(new_n853), .B2(new_n855), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n546), .A2(new_n555), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n572), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n957), .B1(new_n960), .B2(new_n949), .ZN(G57));
endmodule


