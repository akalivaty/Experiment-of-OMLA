//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n451), .B(new_n452), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n464), .A2(G136), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n474), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  OR2_X1    g056(.A1(new_n461), .A2(new_n462), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n475), .ZN(new_n483));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT4), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n464), .A2(new_n486), .A3(G138), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(G114), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(G126), .B2(new_n476), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  OR2_X1    g069(.A1(KEYINPUT5), .A2(G543), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT5), .A2(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G88), .ZN(new_n502));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OAI21_X1  g080(.A(G543), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n501), .A2(new_n502), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n497), .A2(G62), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT69), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n508), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n507), .A2(new_n512), .ZN(G166));
  AOI22_X1  g088(.A1(new_n495), .A2(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT7), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(KEYINPUT7), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(G89), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n506), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g096(.A(KEYINPUT70), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G51), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n497), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n521), .B2(new_n522), .ZN(new_n529));
  INV_X1    g104(.A(new_n526), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT71), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n519), .B1(new_n527), .B2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(new_n523), .A2(G52), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  AND2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n539), .A2(G651), .B1(new_n514), .B2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n533), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  NAND3_X1  g117(.A1(new_n497), .A2(new_n500), .A3(G81), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n497), .B2(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n543), .B1(new_n546), .B2(new_n508), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n521), .B2(new_n522), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT72), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n544), .B1(new_n537), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G651), .B1(new_n514), .B2(G81), .ZN(new_n553));
  AOI21_X1  g128(.A(KEYINPUT70), .B1(new_n500), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n522), .ZN(new_n555));
  OAI21_X1  g130(.A(G43), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n553), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT73), .Z(G188));
  INV_X1    g140(.A(new_n506), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G53), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n568), .A2(new_n569), .B1(G91), .B2(new_n514), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n537), .B(KEYINPUT74), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g148(.A1(G78), .A2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n575), .ZN(G299));
  NAND2_X1  g151(.A1(new_n527), .A2(new_n531), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(new_n518), .ZN(G286));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n514), .A2(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n566), .A2(G49), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT75), .ZN(G288));
  AOI22_X1  g159(.A1(new_n497), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n508), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n501), .A2(new_n587), .B1(new_n588), .B2(new_n506), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n586), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n523), .A2(G47), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n514), .A2(G85), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(new_n508), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n571), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g172(.A1(G79), .A2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n523), .A2(G54), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n497), .A2(new_n500), .A3(G92), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT10), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n595), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n595), .B1(new_n604), .B2(G868), .ZN(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G280));
  INV_X1    g185(.A(G860), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n603), .B1(G559), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT76), .ZN(G148));
  NAND2_X1  g188(.A1(new_n550), .A2(new_n558), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n607), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n603), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n482), .A2(new_n466), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT77), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  AOI22_X1  g200(.A1(G123), .A2(new_n476), .B1(new_n464), .B2(G135), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(G111), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n627), .A2(KEYINPUT78), .B1(new_n628), .B2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(KEYINPUT78), .B2(new_n627), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND3_X1  g207(.A1(new_n624), .A2(new_n625), .A3(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(KEYINPUT14), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT79), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT80), .ZN(new_n648));
  OAI21_X1  g223(.A(G14), .B1(new_n645), .B2(new_n646), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(G401));
  INV_X1    g225(.A(KEYINPUT18), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2096), .B(G2100), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n654), .B2(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT81), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT20), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n665), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n665), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G33), .ZN(new_n682));
  NAND2_X1  g257(.A1(G115), .A2(G2104), .ZN(new_n683));
  INV_X1    g258(.A(G127), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n463), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n475), .B1(new_n685), .B2(KEYINPUT88), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(KEYINPUT88), .B2(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT25), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G139), .B2(new_n464), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT90), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n682), .B1(new_n695), .B2(new_n681), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n696), .A2(G2072), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT91), .Z(new_n698));
  NOR2_X1   g273(.A1(G4), .A2(G16), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n604), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT85), .B(G1348), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT82), .B(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G26), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  OAI21_X1  g280(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n706));
  INV_X1    g281(.A(G116), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G2105), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT86), .Z(new_n709));
  AOI22_X1  g284(.A1(G128), .A2(new_n476), .B1(new_n464), .B2(G140), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(G29), .ZN(new_n712));
  INV_X1    g287(.A(G2067), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G19), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n559), .B2(new_n715), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(G1341), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n702), .B(new_n718), .C1(G1341), .C2(new_n717), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n715), .A2(G20), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT23), .Z(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G299), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT96), .B(G1956), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT31), .B(G11), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT93), .B(G28), .Z(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n729), .B2(KEYINPUT30), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(KEYINPUT30), .B2(new_n729), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(new_n731), .C1(new_n631), .C2(new_n703), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G34), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n703), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT92), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G160), .B2(G29), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n732), .B1(new_n736), .B2(G2084), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n681), .A2(G32), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT26), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n466), .A2(G105), .ZN(new_n741));
  INV_X1    g316(.A(G141), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n483), .B2(new_n742), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n740), .B(new_n743), .C1(G129), .C2(new_n476), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n738), .B1(new_n744), .B2(new_n681), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n715), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n715), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n727), .A2(new_n737), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n736), .A2(G2084), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT94), .Z(new_n754));
  INV_X1    g329(.A(new_n703), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(G35), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G162), .B2(new_n755), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G2090), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n755), .A2(G27), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G164), .B2(new_n755), .ZN(new_n764));
  INV_X1    g339(.A(G2078), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n760), .B2(new_n759), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n715), .A2(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G168), .B2(new_n715), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1966), .ZN(new_n770));
  NOR4_X1   g345(.A1(new_n752), .A2(new_n762), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n696), .A2(G2072), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n721), .A2(new_n722), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  OR3_X1    g348(.A1(new_n698), .A2(KEYINPUT97), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(KEYINPUT97), .B1(new_n698), .B2(new_n773), .ZN(new_n775));
  MUX2_X1   g350(.A(G23), .B(new_n583), .S(G16), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT33), .ZN(new_n777));
  INV_X1    g352(.A(G1976), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G22), .ZN(new_n780));
  OR3_X1    g355(.A1(new_n780), .A2(KEYINPUT83), .A3(G16), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT83), .B1(new_n780), .B2(G16), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n781), .B(new_n782), .C1(G166), .C2(new_n715), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1971), .ZN(new_n784));
  NOR2_X1   g359(.A1(G6), .A2(G16), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n586), .A2(new_n589), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT32), .B(G1981), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n779), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n715), .A2(G24), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G290), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G1986), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n464), .A2(G131), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n476), .A2(G119), .ZN(new_n798));
  OR2_X1    g373(.A1(G95), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G25), .B(new_n801), .S(new_n755), .Z(new_n802));
  XOR2_X1   g377(.A(KEYINPUT35), .B(G1991), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n795), .A2(G1986), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n792), .A2(new_n796), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n790), .A2(new_n791), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT36), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT84), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n809), .A2(KEYINPUT84), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n774), .A2(new_n775), .B1(new_n811), .B2(new_n812), .ZN(G311));
  NAND2_X1  g388(.A1(new_n774), .A2(new_n775), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n812), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(G150));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  INV_X1    g392(.A(G67), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n537), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G651), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n821));
  OAI21_X1  g396(.A(G55), .B1(new_n554), .B2(new_n555), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT98), .B(G93), .Z(new_n823));
  AND3_X1   g398(.A1(new_n823), .A2(new_n497), .A3(new_n500), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n821), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G55), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n521), .B2(new_n522), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n828), .A2(KEYINPUT99), .A3(new_n824), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n820), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G860), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT101), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT37), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n604), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n553), .A2(new_n556), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n836), .B(new_n820), .C1(new_n826), .C2(new_n829), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n822), .A2(new_n825), .A3(new_n821), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT99), .B1(new_n828), .B2(new_n824), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n839), .A2(new_n840), .B1(G651), .B2(new_n819), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n837), .B(new_n838), .C1(new_n614), .C2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n830), .A2(new_n559), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n838), .B1(new_n844), .B2(new_n837), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n835), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n611), .B1(new_n848), .B2(KEYINPUT39), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n833), .B1(new_n849), .B2(new_n850), .ZN(G145));
  XNOR2_X1  g426(.A(new_n493), .B(new_n711), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n744), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n744), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n695), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n620), .B(new_n801), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n476), .A2(G130), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n464), .A2(G142), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n860), .A2(new_n475), .A3(G118), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n475), .B2(G118), .ZN(new_n862));
  OR2_X1    g437(.A1(G106), .A2(G2105), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(G2104), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n858), .B(new_n859), .C1(new_n861), .C2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n857), .B(new_n865), .Z(new_n866));
  NAND3_X1  g441(.A1(new_n853), .A2(new_n693), .A3(new_n854), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n856), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n856), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n472), .B(new_n480), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n631), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT104), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n868), .A2(new_n869), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT103), .B1(new_n875), .B2(new_n872), .ZN(new_n876));
  OAI211_X1 g451(.A(KEYINPUT103), .B(new_n872), .C1(new_n868), .C2(new_n869), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n874), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g455(.A(new_n846), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n616), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n602), .A2(new_n600), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n883), .A2(new_n575), .A3(new_n570), .A4(new_n599), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n603), .A2(G299), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT105), .B1(new_n886), .B2(KEYINPUT41), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n884), .A2(new_n885), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n888), .B(KEYINPUT107), .C1(new_n882), .C2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n583), .B(KEYINPUT108), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n786), .ZN(new_n900));
  XNOR2_X1  g475(.A(G290), .B(G166), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(KEYINPUT42), .Z(new_n903));
  OR3_X1    g478(.A1(new_n882), .A2(new_n897), .A3(KEYINPUT107), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n898), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n898), .B2(new_n904), .ZN(new_n906));
  OAI21_X1  g481(.A(G868), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(G868), .B2(new_n841), .ZN(G295));
  OAI21_X1  g483(.A(new_n907), .B1(G868), .B2(new_n841), .ZN(G331));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n910));
  NAND2_X1  g485(.A1(G301), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n533), .A2(new_n540), .A3(KEYINPUT109), .ZN(new_n912));
  AND3_X1   g487(.A1(G168), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(G168), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n843), .B2(new_n845), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n837), .B1(new_n841), .B2(new_n614), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT100), .ZN(new_n918));
  NAND3_X1  g493(.A1(G286), .A2(new_n910), .A3(G301), .ZN(new_n919));
  NAND3_X1  g494(.A1(G168), .A2(new_n911), .A3(new_n912), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n921), .A3(new_n842), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n916), .A2(new_n887), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT110), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n916), .A2(new_n922), .A3(new_n925), .A4(new_n887), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT41), .B1(new_n884), .B2(new_n885), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n887), .B2(new_n894), .ZN(new_n928));
  INV_X1    g503(.A(new_n922), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n921), .B1(new_n918), .B2(new_n842), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n924), .A2(new_n926), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n902), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n932), .A2(KEYINPUT111), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT111), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n896), .B1(new_n930), .B2(new_n929), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n902), .A3(new_n923), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n902), .B1(new_n937), .B2(new_n923), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n940), .A2(KEYINPUT43), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(KEYINPUT44), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n938), .A2(new_n945), .A3(new_n939), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n934), .B2(new_n935), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n940), .B2(new_n942), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT112), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n952));
  AOI211_X1 g527(.A(new_n952), .B(KEYINPUT44), .C1(new_n947), .C2(new_n948), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n944), .B1(new_n951), .B2(new_n953), .ZN(G397));
  INV_X1    g529(.A(KEYINPUT52), .ZN(new_n955));
  INV_X1    g530(.A(G8), .ZN(new_n956));
  AOI21_X1  g531(.A(G1384), .B1(new_n488), .B2(new_n492), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n467), .A2(new_n471), .A3(G40), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n583), .A2(new_n778), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT116), .ZN(new_n962));
  NOR2_X1   g537(.A1(G305), .A2(G1981), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT49), .ZN(new_n964));
  INV_X1    g539(.A(G1981), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n786), .A2(new_n965), .ZN(new_n966));
  OR3_X1    g541(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n964), .B1(new_n963), .B2(new_n966), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n959), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT52), .B1(G288), .B2(new_n778), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n970), .A2(new_n959), .A3(new_n960), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n962), .A2(new_n972), .A3(KEYINPUT117), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT117), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n959), .A2(new_n960), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT116), .B1(new_n975), .B2(KEYINPUT52), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n977), .B(new_n955), .C1(new_n959), .C2(new_n960), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n969), .A2(new_n971), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n974), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n973), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n958), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n493), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n957), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n760), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1971), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT113), .B(G1384), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n493), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n958), .B1(new_n957), .B2(KEYINPUT45), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G166), .B2(new_n956), .ZN(new_n1001));
  NAND4_X1  g576(.A1(G303), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n996), .A2(G8), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n996), .B2(G8), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n982), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n983), .B1(new_n985), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n957), .A2(KEYINPUT45), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(G2078), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n958), .B1(new_n957), .B2(new_n987), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n750), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT125), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1014), .A2(new_n1017), .A3(KEYINPUT125), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1010), .A2(new_n765), .A3(new_n992), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1012), .ZN(new_n1024));
  AOI21_X1  g599(.A(G301), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n493), .A2(new_n991), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n1009), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1027), .A2(new_n958), .A3(new_n992), .A4(new_n1013), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1017), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G171), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1008), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G2084), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n986), .A2(new_n1032), .A3(new_n988), .ZN(new_n1033));
  INV_X1    g608(.A(G1966), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1011), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(new_n994), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G8), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G168), .A2(new_n956), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT51), .B1(new_n1039), .B2(KEYINPUT123), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1041), .ZN(new_n1043));
  OAI211_X1 g618(.A(G8), .B(new_n1043), .C1(new_n1037), .C2(G286), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1029), .B2(G171), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1014), .A2(new_n1017), .A3(KEYINPUT125), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT125), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1050));
  OAI211_X1 g625(.A(G301), .B(new_n1024), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1045), .A2(new_n1046), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1007), .A2(new_n1031), .A3(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT56), .B(G2072), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1010), .A2(new_n992), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1956), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1010), .A2(KEYINPUT120), .A3(new_n992), .A4(new_n1054), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT119), .B1(new_n568), .B2(new_n569), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(KEYINPUT57), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(G299), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1057), .A2(new_n1064), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(KEYINPUT61), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n957), .A2(new_n958), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n957), .A2(KEYINPUT121), .A3(new_n958), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT58), .B(G1341), .Z(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1996), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1010), .A2(new_n1077), .A3(new_n992), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1070), .B1(new_n1079), .B2(new_n559), .ZN(new_n1080));
  AOI211_X1 g655(.A(KEYINPUT59), .B(new_n614), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1074), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT121), .B1(new_n957), .B2(new_n958), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n713), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1348), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n604), .A3(new_n1086), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1080), .A2(new_n1081), .B1(KEYINPUT60), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n603), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1090), .A2(KEYINPUT60), .A3(new_n1087), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1066), .A2(KEYINPUT61), .A3(new_n1068), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT122), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AND4_X1   g672(.A1(new_n1069), .A2(new_n1092), .A3(new_n1094), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1068), .A2(new_n604), .A3(new_n1089), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n1066), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1053), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1038), .A2(G286), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n982), .A2(new_n1006), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT118), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n979), .A2(new_n980), .A3(new_n1104), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1006), .A2(new_n1102), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1004), .A2(new_n962), .A3(new_n972), .ZN(new_n1112));
  NOR2_X1   g687(.A1(G288), .A2(G1976), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n969), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n959), .B1(new_n1114), .B2(new_n963), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n982), .A2(new_n1025), .A3(new_n1006), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1045), .A2(new_n1118), .A3(new_n1046), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1116), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1101), .A2(new_n1111), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1027), .A2(new_n983), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT114), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n744), .B(G1996), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n711), .B(new_n713), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n803), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n801), .A2(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n801), .A2(new_n1129), .ZN(new_n1131));
  OR3_X1    g706(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(G290), .B(G1986), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1125), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1123), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1125), .A2(new_n1077), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT46), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1127), .A2(new_n744), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1125), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT47), .Z(new_n1141));
  NOR2_X1   g716(.A1(G290), .A2(G1986), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1125), .A2(new_n1142), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1143), .A2(KEYINPUT127), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(KEYINPUT127), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1144), .A2(KEYINPUT48), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT48), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1132), .A2(new_n1125), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n711), .A2(G2067), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n1130), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1125), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1141), .A2(new_n1149), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1135), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g732(.A1(G401), .A2(G229), .A3(new_n459), .A4(G227), .ZN(new_n1159));
  NAND3_X1  g733(.A1(new_n879), .A2(new_n949), .A3(new_n1159), .ZN(G225));
  INV_X1    g734(.A(G225), .ZN(G308));
endmodule


