//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n566,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n598, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XOR2_X1   g020(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n463), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n468), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n471), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT3), .B(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G125), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n470), .B1(new_n484), .B2(new_n475), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT67), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n474), .B1(new_n482), .B2(new_n486), .ZN(G160));
  AND4_X1   g062(.A1(G2105), .A2(new_n468), .A3(new_n469), .A4(new_n471), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n470), .A2(G112), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n472), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(G136), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n468), .A2(new_n469), .A3(new_n497), .A4(new_n471), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(G138), .A3(new_n470), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(KEYINPUT4), .A2(new_n498), .B1(new_n502), .B2(new_n483), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G2105), .ZN(new_n508));
  NOR3_X1   g083(.A1(new_n470), .A2(KEYINPUT70), .A3(G114), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G126), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n468), .A2(new_n469), .A3(G2105), .A4(new_n471), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n503), .A2(new_n513), .ZN(G164));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n521), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(G89), .B1(new_n517), .B2(new_n518), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n516), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n528), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT72), .B(G52), .Z(new_n541));
  NOR2_X1   g116(.A1(new_n525), .A2(new_n541), .ZN(new_n542));
  AOI211_X1 g117(.A(new_n540), .B(new_n542), .C1(G90), .C2(new_n520), .ZN(G171));
  NAND2_X1  g118(.A1(new_n524), .A2(G43), .ZN(new_n544));
  INV_X1    g119(.A(new_n520), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT73), .B(G81), .Z(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n528), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n524), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n528), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n520), .A2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G299));
  XNOR2_X1  g140(.A(G171), .B(KEYINPUT75), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n520), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n524), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  AOI22_X1  g148(.A1(new_n520), .A2(G86), .B1(new_n524), .B2(G48), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n528), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G305));
  AND2_X1   g152(.A1(new_n515), .A2(G60), .ZN(new_n578));
  AND2_X1   g153(.A1(G72), .A2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(KEYINPUT76), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(KEYINPUT76), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n520), .A2(G85), .B1(new_n524), .B2(G47), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(new_n520), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT10), .Z(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n516), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n524), .B2(G54), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(G868), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n566), .B2(G868), .ZN(G284));
  AOI21_X1  g168(.A(new_n592), .B1(new_n566), .B2(G868), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n564), .B2(G868), .ZN(G297));
  OAI21_X1  g171(.A(new_n595), .B1(new_n564), .B2(G868), .ZN(G280));
  INV_X1    g172(.A(new_n591), .ZN(new_n598));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n483), .A2(new_n464), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT13), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(G2100), .ZN(new_n608));
  OR2_X1    g183(.A1(G99), .A2(G2105), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n609), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n610));
  INV_X1    g185(.A(G123), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n512), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G135), .B2(new_n493), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(G2096), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(G2096), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n608), .A2(new_n615), .A3(new_n616), .ZN(G156));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2435), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT77), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(G2427), .B(G2430), .Z(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(KEYINPUT14), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(G2451), .B(G2454), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n624), .B(new_n628), .Z(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(new_n632), .A3(G14), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT78), .Z(G401));
  XOR2_X1   g209(.A(G2072), .B(G2078), .Z(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT79), .Z(new_n636));
  XNOR2_X1  g211(.A(G2084), .B(G2090), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NOR3_X1   g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT18), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n636), .B(KEYINPUT17), .ZN(new_n642));
  INV_X1    g217(.A(new_n636), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n637), .B1(new_n643), .B2(new_n638), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n645));
  OAI22_X1  g220(.A1(new_n642), .A2(new_n639), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n637), .A2(new_n638), .ZN(new_n648));
  AOI211_X1 g223(.A(new_n641), .B(new_n647), .C1(new_n642), .C2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT82), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT81), .B(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n655), .A2(new_n658), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  AOI211_X1 g238(.A(new_n660), .B(new_n663), .C1(new_n655), .C2(new_n659), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G229));
  INV_X1    g245(.A(G29), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G26), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n488), .A2(G128), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n470), .A2(G116), .ZN(new_n675));
  OAI21_X1  g250(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G140), .B2(new_n493), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT91), .ZN(new_n679));
  AND3_X1   g254(.A1(new_n679), .A2(KEYINPUT92), .A3(G29), .ZN(new_n680));
  AOI21_X1  g255(.A(KEYINPUT92), .B1(new_n679), .B2(G29), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n673), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G2067), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NOR2_X1   g260(.A1(G171), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G5), .B2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1341), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n685), .A2(KEYINPUT85), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(KEYINPUT85), .ZN(new_n691));
  AND3_X1   g266(.A1(new_n690), .A2(G19), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n550), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n691), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n688), .A2(G1961), .B1(new_n689), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G1961), .ZN(new_n697));
  NOR2_X1   g272(.A1(G168), .A2(new_n685), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n685), .B2(G21), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n687), .A2(new_n697), .B1(G1966), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G1966), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n699), .A2(new_n702), .B1(G29), .B2(new_n613), .ZN(new_n703));
  INV_X1    g278(.A(G11), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT31), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT31), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT30), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(G28), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n671), .B1(new_n707), .B2(G28), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n705), .B(new_n706), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n695), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G1341), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n696), .A2(new_n701), .A3(new_n703), .A4(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT24), .ZN(new_n714));
  INV_X1    g289(.A(G34), .ZN(new_n715));
  AOI21_X1  g290(.A(G29), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n714), .B2(new_n715), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G160), .B2(new_n671), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G2084), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n671), .A2(G32), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT26), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n723), .A2(new_n724), .B1(G105), .B2(new_n464), .ZN(new_n725));
  INV_X1    g300(.A(G129), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n512), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G141), .B2(new_n493), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n720), .B1(new_n728), .B2(new_n671), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT27), .B(G1996), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT94), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n729), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n719), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G4), .A2(G16), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n598), .B2(G16), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT90), .B(G1348), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n690), .A2(G20), .A3(new_n691), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT23), .Z(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G299), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G1956), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR4_X1   g317(.A1(new_n713), .A2(new_n733), .A3(new_n737), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G29), .A2(G35), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G162), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT29), .ZN(new_n746));
  INV_X1    g321(.A(G2090), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT25), .Z(new_n750));
  AOI22_X1  g325(.A1(new_n483), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n470), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G139), .B2(new_n493), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G29), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G29), .B2(G33), .ZN(new_n756));
  INV_X1    g331(.A(G2072), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n671), .A2(G27), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G164), .B2(new_n671), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2078), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n758), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  AND4_X1   g338(.A1(new_n684), .A2(new_n743), .A3(new_n748), .A4(new_n763), .ZN(new_n764));
  MUX2_X1   g339(.A(G6), .B(G305), .S(G16), .Z(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT86), .Z(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT32), .B(G1981), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n768), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G23), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT87), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G288), .B2(new_n685), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT33), .B(G1976), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n694), .A2(G22), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G166), .B2(new_n694), .ZN(new_n777));
  INV_X1    g352(.A(G1971), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n769), .A2(new_n770), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT88), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT34), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n488), .A2(G119), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT84), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n788));
  INV_X1    g363(.A(G107), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G2105), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n493), .B2(G131), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G25), .B(new_n792), .S(G29), .Z(new_n793));
  XOR2_X1   g368(.A(KEYINPUT35), .B(G1991), .Z(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n793), .B(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G24), .B(G290), .S(new_n694), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G1986), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n797), .A2(G1986), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n796), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n784), .A2(new_n785), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n764), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(G311));
  XOR2_X1   g381(.A(G311), .B(KEYINPUT95), .Z(G150));
  NAND2_X1  g382(.A1(new_n598), .A2(G559), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n524), .A2(G55), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT96), .B(G93), .Z(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n545), .B2(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n528), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n550), .B(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n809), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT98), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT97), .B(G860), .Z(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n817), .B2(new_n818), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n821), .B1(new_n812), .B2(new_n814), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(G145));
  INV_X1    g401(.A(KEYINPUT100), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n754), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n728), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n792), .B(new_n606), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n503), .B2(new_n513), .ZN(new_n833));
  OAI21_X1  g408(.A(KEYINPUT70), .B1(new_n470), .B2(G114), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n506), .A2(new_n507), .A3(G2105), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n504), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n488), .B2(G126), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n502), .A2(new_n483), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n840), .A3(KEYINPUT99), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n833), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n679), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n488), .A2(G130), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n470), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G142), .B2(new_n493), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n843), .B(new_n848), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n831), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(G162), .B(new_n614), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G160), .ZN(new_n852));
  AOI21_X1  g427(.A(G37), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n850), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g430(.A(new_n591), .B1(KEYINPUT101), .B2(new_n564), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(KEYINPUT101), .B2(new_n564), .ZN(new_n857));
  OR3_X1    g432(.A1(new_n598), .A2(KEYINPUT101), .A3(new_n564), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(KEYINPUT41), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n601), .B(new_n816), .Z(new_n862));
  MUX2_X1   g437(.A(new_n860), .B(new_n861), .S(new_n862), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT42), .ZN(new_n864));
  XNOR2_X1  g439(.A(G290), .B(G305), .ZN(new_n865));
  XNOR2_X1  g440(.A(G166), .B(G288), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n864), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(G868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(G868), .B2(new_n815), .ZN(G295));
  OAI21_X1  g445(.A(new_n869), .B1(G868), .B2(new_n815), .ZN(G331));
  NOR2_X1   g446(.A1(G171), .A2(G168), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(new_n566), .B2(G168), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(new_n816), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n861), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n859), .B2(new_n874), .ZN(new_n876));
  AOI21_X1  g451(.A(G37), .B1(new_n876), .B2(new_n867), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n867), .B2(new_n876), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT43), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT102), .B1(new_n878), .B2(KEYINPUT43), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT44), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n879), .B(new_n881), .ZN(G397));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n883));
  INV_X1    g458(.A(G1384), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n842), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT45), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n883), .B1(new_n842), .B2(new_n884), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n474), .ZN(new_n890));
  AOI211_X1 g465(.A(new_n481), .B(new_n470), .C1(new_n484), .C2(new_n475), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT67), .B1(new_n479), .B2(G2105), .ZN(new_n892));
  OAI211_X1 g467(.A(G40), .B(new_n890), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n679), .B(new_n683), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(new_n728), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT127), .Z(new_n898));
  NOR2_X1   g473(.A1(new_n895), .A2(G1996), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT46), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(KEYINPUT47), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n728), .B(G1996), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n896), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n792), .B(new_n795), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT105), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n895), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT48), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n895), .A2(G1986), .A3(G290), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n904), .A2(new_n794), .A3(new_n787), .A4(new_n791), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(G2067), .B2(new_n679), .ZN(new_n913));
  INV_X1    g488(.A(new_n895), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n902), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n884), .B1(new_n503), .B2(new_n513), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT50), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT50), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(new_n884), .C1(new_n503), .C2(new_n513), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(KEYINPUT107), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n922), .A3(KEYINPUT50), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n893), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(KEYINPUT111), .B(G2084), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n893), .B1(new_n886), .B2(new_n917), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n837), .A2(new_n840), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(KEYINPUT45), .A3(new_n884), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n702), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(G8), .ZN(new_n933));
  INV_X1    g508(.A(G8), .ZN(new_n934));
  NOR2_X1   g509(.A1(G168), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(KEYINPUT51), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n938), .B(G8), .C1(new_n932), .C2(G286), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT118), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n932), .B2(new_n935), .ZN(new_n941));
  AOI211_X1 g516(.A(KEYINPUT118), .B(new_n936), .C1(new_n926), .C2(new_n931), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n937), .B(new_n939), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n921), .A2(new_n923), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n747), .A3(new_n894), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT108), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n945), .A2(new_n948), .A3(new_n747), .A4(new_n894), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n833), .A2(new_n841), .A3(KEYINPUT45), .A4(new_n884), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n917), .A2(new_n886), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n894), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n927), .A2(KEYINPUT106), .A3(new_n950), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n778), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n947), .A2(new_n949), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G303), .A2(G8), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT55), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(G8), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(G305), .A2(G1981), .ZN(new_n962));
  INV_X1    g537(.A(G1981), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n574), .A2(new_n963), .A3(new_n576), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT49), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n917), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n934), .B1(new_n894), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n962), .A2(KEYINPUT49), .A3(new_n964), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1976), .ZN(new_n972));
  OR2_X1    g547(.A1(G288), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT52), .B1(G288), .B2(new_n972), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n973), .B(G8), .C1(new_n917), .C2(new_n893), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT52), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n971), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n961), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n894), .A2(new_n918), .A3(new_n920), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n980), .A2(G2090), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n956), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n959), .B1(new_n982), .B2(new_n934), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n944), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G2078), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n952), .A2(new_n953), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT106), .B1(new_n927), .B2(new_n950), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT114), .B1(new_n945), .B2(new_n894), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n994), .B(new_n893), .C1(new_n921), .C2(new_n923), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT119), .B(G1961), .Z(new_n996));
  NOR3_X1   g571(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n986), .A2(KEYINPUT53), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n930), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT120), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n920), .A2(KEYINPUT107), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n919), .B1(new_n928), .B2(new_n884), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n923), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n894), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n994), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n924), .A2(KEYINPUT114), .ZN(new_n1007));
  INV_X1    g582(.A(new_n996), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n1010));
  INV_X1    g585(.A(new_n999), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n992), .B1(new_n1000), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT121), .B1(new_n1013), .B2(G301), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1010), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n991), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n566), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n985), .A2(new_n1020), .A3(KEYINPUT125), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT125), .B1(new_n985), .B2(new_n1020), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  AOI211_X1 g602(.A(new_n934), .B(G286), .C1(new_n926), .C2(new_n931), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n983), .A2(new_n961), .A3(new_n978), .A4(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n932), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n957), .A2(G8), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n959), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1027), .A2(new_n1029), .B1(new_n979), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n957), .A2(G8), .A3(new_n960), .A4(new_n978), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G288), .A2(G1976), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT109), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n971), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n964), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n969), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1034), .A2(new_n1035), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1035), .B1(new_n1034), .B2(new_n1040), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1026), .B1(new_n1033), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1029), .A2(new_n1027), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n979), .A2(new_n1032), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1042), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1034), .A2(new_n1035), .A3(new_n1040), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(KEYINPUT112), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1044), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G40), .ZN(new_n1053));
  NOR4_X1   g628(.A1(new_n485), .A2(new_n474), .A3(new_n1053), .A4(new_n998), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n950), .B(new_n1054), .C1(new_n887), .C2(new_n888), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n991), .A2(new_n1009), .A3(new_n1055), .A4(G301), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1014), .A2(new_n1019), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1348), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1006), .A2(new_n1062), .A3(new_n1007), .ZN(new_n1063));
  OR3_X1    g638(.A1(new_n893), .A2(KEYINPUT113), .A3(new_n917), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT113), .B1(new_n893), .B2(new_n917), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n683), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n559), .A2(KEYINPUT57), .A3(new_n563), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n1070));
  INV_X1    g645(.A(new_n563), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n558), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n980), .A2(new_n741), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n927), .A2(new_n950), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1077), .A2(new_n598), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1074), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1068), .A2(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1079), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1077), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1085), .A3(KEYINPUT61), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1082), .B(new_n1077), .C1(new_n1084), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1063), .A2(new_n1067), .A3(KEYINPUT60), .A4(new_n591), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT58), .B(G1341), .Z(new_n1091));
  NAND3_X1  g666(.A1(new_n1064), .A2(new_n1065), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1996), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n927), .A2(new_n1093), .A3(new_n950), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n693), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(KEYINPUT115), .A2(KEYINPUT59), .ZN(new_n1096));
  NAND2_X1  g671(.A1(KEYINPUT115), .A2(KEYINPUT59), .ZN(new_n1097));
  XOR2_X1   g672(.A(new_n1097), .B(KEYINPUT116), .Z(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  OR3_X1    g674(.A1(new_n1095), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1089), .A2(new_n1090), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1068), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1063), .A2(new_n1067), .A3(KEYINPUT60), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1105), .A2(new_n598), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1081), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n943), .A2(new_n979), .A3(new_n983), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(G301), .B(new_n991), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n991), .A2(new_n1009), .A3(new_n1055), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1060), .B1(new_n1112), .B2(G171), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1111), .A2(KEYINPUT123), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT123), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1108), .B(new_n1110), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1052), .B1(new_n1061), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT124), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1116), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1114), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1105), .A2(new_n598), .A3(new_n1106), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1123), .A2(new_n1090), .A3(new_n1102), .A4(new_n1089), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1109), .B1(new_n1124), .B2(new_n1081), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1120), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n1052), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1025), .B1(new_n1119), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n914), .A2(G1986), .A3(G290), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n909), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT104), .Z(new_n1133));
  NOR2_X1   g708(.A1(new_n1133), .A2(new_n907), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1129), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1025), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1126), .A2(new_n1127), .A3(new_n1052), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1127), .B1(new_n1126), .B2(new_n1052), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT126), .B1(new_n1140), .B2(new_n1134), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n916), .B1(new_n1136), .B2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g717(.A1(G227), .A2(G229), .A3(new_n461), .A4(G401), .ZN(new_n1144));
  NAND3_X1  g718(.A1(new_n879), .A2(new_n854), .A3(new_n1144), .ZN(G225));
  INV_X1    g719(.A(G225), .ZN(G308));
endmodule


