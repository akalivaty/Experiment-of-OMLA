

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742;

  XNOR2_X1 U368 ( .A(G116), .B(G113), .ZN(n422) );
  INV_X2 U369 ( .A(G953), .ZN(n729) );
  INV_X2 U370 ( .A(n522), .ZN(n348) );
  XNOR2_X2 U371 ( .A(n390), .B(n389), .ZN(n522) );
  OR2_X2 U372 ( .A1(n716), .A2(G902), .ZN(n390) );
  NAND2_X2 U373 ( .A1(n348), .A2(n524), .ZN(n374) );
  AND2_X2 U374 ( .A1(n360), .A2(n601), .ZN(n665) );
  NOR2_X2 U375 ( .A1(n544), .A2(n677), .ZN(n514) );
  INV_X2 U376 ( .A(G128), .ZN(n375) );
  XNOR2_X1 U377 ( .A(n367), .B(n488), .ZN(n566) );
  XNOR2_X1 U378 ( .A(n361), .B(KEYINPUT0), .ZN(n584) );
  OR2_X1 U379 ( .A1(n517), .A2(n370), .ZN(n692) );
  XNOR2_X1 U380 ( .A(n406), .B(n405), .ZN(n523) );
  XNOR2_X1 U381 ( .A(n366), .B(n362), .ZN(n625) );
  XNOR2_X1 U382 ( .A(n428), .B(n407), .ZN(n452) );
  XNOR2_X1 U383 ( .A(G101), .B(KEYINPUT69), .ZN(n421) );
  XNOR2_X1 U384 ( .A(KEYINPUT3), .B(G119), .ZN(n423) );
  OR2_X2 U385 ( .A1(n672), .A2(n671), .ZN(n575) );
  XNOR2_X1 U386 ( .A(n391), .B(n392), .ZN(n716) );
  NOR2_X1 U387 ( .A1(n739), .A2(n741), .ZN(n372) );
  AND2_X1 U388 ( .A1(n565), .A2(n566), .ZN(n567) );
  OR2_X1 U389 ( .A1(n619), .A2(n604), .ZN(n437) );
  NOR2_X1 U390 ( .A1(n625), .A2(G902), .ZN(n406) );
  NOR2_X1 U391 ( .A1(n712), .A2(G902), .ZN(n459) );
  INV_X1 U392 ( .A(KEYINPUT46), .ZN(n371) );
  INV_X1 U393 ( .A(KEYINPUT48), .ZN(n386) );
  XNOR2_X1 U394 ( .A(KEYINPUT15), .B(G902), .ZN(n561) );
  XNOR2_X1 U395 ( .A(n452), .B(n451), .ZN(n483) );
  XNOR2_X1 U396 ( .A(KEYINPUT4), .B(G131), .ZN(n451) );
  OR2_X1 U397 ( .A1(n575), .A2(n381), .ZN(n378) );
  NAND2_X1 U398 ( .A1(n382), .A2(KEYINPUT33), .ZN(n381) );
  INV_X1 U399 ( .A(n569), .ZN(n382) );
  XNOR2_X1 U400 ( .A(n350), .B(n471), .ZN(n675) );
  XNOR2_X1 U401 ( .A(n470), .B(KEYINPUT25), .ZN(n471) );
  XNOR2_X1 U402 ( .A(n441), .B(n440), .ZN(n537) );
  XNOR2_X1 U403 ( .A(n596), .B(KEYINPUT45), .ZN(n360) );
  XNOR2_X1 U404 ( .A(G128), .B(G119), .ZN(n460) );
  XNOR2_X1 U405 ( .A(n725), .B(n464), .ZN(n465) );
  XNOR2_X1 U406 ( .A(n395), .B(n393), .ZN(n467) );
  XNOR2_X1 U407 ( .A(KEYINPUT8), .B(KEYINPUT66), .ZN(n395) );
  NOR2_X1 U408 ( .A1(n394), .A2(G953), .ZN(n393) );
  INV_X1 U409 ( .A(G234), .ZN(n394) );
  INV_X1 U410 ( .A(KEYINPUT11), .ZN(n364) );
  XNOR2_X1 U411 ( .A(n399), .B(n401), .ZN(n365) );
  XOR2_X1 U412 ( .A(G140), .B(G113), .Z(n399) );
  XOR2_X1 U413 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n401) );
  XNOR2_X1 U414 ( .A(n483), .B(n463), .ZN(n724) );
  INV_X1 U415 ( .A(G110), .ZN(n419) );
  NAND2_X1 U416 ( .A1(G234), .A2(G237), .ZN(n445) );
  XNOR2_X1 U417 ( .A(n656), .B(n525), .ZN(n558) );
  NOR2_X1 U418 ( .A1(n547), .A2(n370), .ZN(n369) );
  INV_X1 U419 ( .A(G478), .ZN(n389) );
  BUF_X1 U420 ( .A(n675), .Z(n359) );
  NAND2_X1 U421 ( .A1(n584), .A2(n448), .ZN(n450) );
  NOR2_X1 U422 ( .A1(n519), .A2(n508), .ZN(n531) );
  XNOR2_X1 U423 ( .A(n536), .B(n535), .ZN(n539) );
  AND2_X2 U424 ( .A1(n558), .A2(n543), .ZN(n693) );
  AND2_X1 U425 ( .A1(n517), .A2(n370), .ZN(n690) );
  XOR2_X1 U426 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n474) );
  XNOR2_X1 U427 ( .A(G137), .B(G146), .ZN(n476) );
  INV_X1 U428 ( .A(n662), .ZN(n559) );
  XNOR2_X1 U429 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n427) );
  OR2_X1 U430 ( .A1(G237), .A2(G902), .ZN(n396) );
  INV_X1 U431 ( .A(G902), .ZN(n484) );
  BUF_X1 U432 ( .A(n600), .Z(n728) );
  OR2_X1 U433 ( .A1(n665), .A2(n605), .ZN(n606) );
  NOR2_X1 U434 ( .A1(n491), .A2(n377), .ZN(n376) );
  INV_X1 U435 ( .A(n384), .ZN(n377) );
  NOR2_X1 U436 ( .A1(n537), .A2(n447), .ZN(n361) );
  XNOR2_X1 U437 ( .A(KEYINPUT70), .B(KEYINPUT16), .ZN(n418) );
  XNOR2_X1 U438 ( .A(n468), .B(n355), .ZN(n720) );
  XNOR2_X1 U439 ( .A(n411), .B(n410), .ZN(n392) );
  XNOR2_X1 U440 ( .A(n365), .B(n363), .ZN(n362) );
  XNOR2_X1 U441 ( .A(n725), .B(n400), .ZN(n366) );
  XNOR2_X1 U442 ( .A(n402), .B(n364), .ZN(n363) );
  XNOR2_X1 U443 ( .A(n724), .B(n458), .ZN(n712) );
  XNOR2_X1 U444 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U445 ( .A(G101), .B(G146), .Z(n456) );
  XNOR2_X1 U446 ( .A(n613), .B(n612), .ZN(n723) );
  XNOR2_X1 U447 ( .A(n373), .B(n521), .ZN(n739) );
  OR2_X1 U448 ( .A1(n557), .A2(n543), .ZN(n373) );
  XNOR2_X1 U449 ( .A(n368), .B(n548), .ZN(n549) );
  XNOR2_X1 U450 ( .A(KEYINPUT36), .B(KEYINPUT90), .ZN(n548) );
  NAND2_X1 U451 ( .A1(n572), .A2(n354), .ZN(n367) );
  INV_X1 U452 ( .A(G143), .ZN(n509) );
  XOR2_X1 U453 ( .A(n497), .B(KEYINPUT30), .Z(n349) );
  NOR2_X1 U454 ( .A1(n720), .A2(G902), .ZN(n350) );
  XOR2_X1 U455 ( .A(KEYINPUT38), .B(KEYINPUT73), .Z(n351) );
  XOR2_X1 U456 ( .A(n372), .B(n371), .Z(n352) );
  AND2_X1 U457 ( .A1(n379), .A2(n378), .ZN(n353) );
  AND2_X1 U458 ( .A1(n487), .A2(n486), .ZN(n354) );
  AND2_X1 U459 ( .A1(G221), .A2(n467), .ZN(n355) );
  AND2_X1 U460 ( .A1(n510), .A2(n675), .ZN(n356) );
  OR2_X1 U461 ( .A1(n380), .A2(n383), .ZN(n357) );
  INV_X1 U462 ( .A(n689), .ZN(n370) );
  XNOR2_X2 U463 ( .A(n431), .B(KEYINPUT10), .ZN(n725) );
  NAND2_X1 U464 ( .A1(n608), .A2(n484), .ZN(n485) );
  XNOR2_X1 U465 ( .A(n482), .B(n483), .ZN(n608) );
  NOR2_X1 U466 ( .A1(n586), .A2(n693), .ZN(n587) );
  XNOR2_X2 U467 ( .A(n582), .B(KEYINPUT1), .ZN(n672) );
  NAND2_X1 U468 ( .A1(n358), .A2(n352), .ZN(n387) );
  XNOR2_X1 U469 ( .A(n551), .B(n388), .ZN(n358) );
  XNOR2_X1 U470 ( .A(n387), .B(n386), .ZN(n385) );
  NAND2_X1 U471 ( .A1(n385), .A2(n397), .ZN(n600) );
  NAND2_X1 U472 ( .A1(n349), .A2(n356), .ZN(n519) );
  NAND2_X1 U473 ( .A1(n360), .A2(n729), .ZN(n631) );
  NAND2_X1 U474 ( .A1(n597), .A2(n360), .ZN(n599) );
  NAND2_X1 U475 ( .A1(n552), .A2(n554), .ZN(n368) );
  AND2_X1 U476 ( .A1(n546), .A2(n369), .ZN(n552) );
  XNOR2_X1 U477 ( .A(n554), .B(n351), .ZN(n517) );
  XNOR2_X2 U478 ( .A(n374), .B(KEYINPUT99), .ZN(n656) );
  XNOR2_X2 U479 ( .A(n375), .B(G143), .ZN(n428) );
  INV_X1 U480 ( .A(n378), .ZN(n380) );
  NAND2_X1 U481 ( .A1(n379), .A2(n384), .ZN(n383) );
  NAND2_X1 U482 ( .A1(n353), .A2(n376), .ZN(n493) );
  NAND2_X1 U483 ( .A1(n575), .A2(n490), .ZN(n379) );
  NAND2_X1 U484 ( .A1(n569), .A2(n490), .ZN(n384) );
  INV_X1 U485 ( .A(KEYINPUT67), .ZN(n388) );
  XNOR2_X1 U486 ( .A(n452), .B(n412), .ZN(n391) );
  NOR2_X1 U487 ( .A1(n562), .A2(n561), .ZN(n597) );
  XNOR2_X1 U488 ( .A(n600), .B(n560), .ZN(n562) );
  NAND2_X2 U489 ( .A1(n607), .A2(n606), .ZN(n710) );
  AND2_X1 U490 ( .A1(n737), .A2(n559), .ZN(n397) );
  INV_X1 U491 ( .A(KEYINPUT72), .ZN(n535) );
  INV_X1 U492 ( .A(KEYINPUT5), .ZN(n475) );
  XNOR2_X1 U493 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U494 ( .A(n478), .B(n477), .ZN(n481) );
  INV_X1 U495 ( .A(n728), .ZN(n601) );
  XNOR2_X1 U496 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U497 ( .A(n481), .B(n480), .ZN(n482) );
  INV_X1 U498 ( .A(G134), .ZN(n407) );
  INV_X1 U499 ( .A(KEYINPUT100), .ZN(n525) );
  XNOR2_X1 U500 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n521) );
  XNOR2_X2 U501 ( .A(G122), .B(G104), .ZN(n417) );
  XNOR2_X1 U502 ( .A(G143), .B(G131), .ZN(n398) );
  XNOR2_X1 U503 ( .A(n417), .B(n398), .ZN(n400) );
  XNOR2_X2 U504 ( .A(G146), .B(G125), .ZN(n431) );
  NOR2_X2 U505 ( .A1(G953), .A2(G237), .ZN(n472) );
  NAND2_X1 U506 ( .A1(G214), .A2(n472), .ZN(n402) );
  XNOR2_X1 U507 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n404) );
  INV_X1 U508 ( .A(G475), .ZN(n403) );
  XOR2_X1 U509 ( .A(KEYINPUT7), .B(G122), .Z(n409) );
  XNOR2_X1 U510 ( .A(G116), .B(G107), .ZN(n408) );
  XNOR2_X1 U511 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U512 ( .A(KEYINPUT98), .B(KEYINPUT9), .Z(n412) );
  NAND2_X1 U513 ( .A1(G217), .A2(n467), .ZN(n411) );
  OR2_X1 U514 ( .A1(n523), .A2(n348), .ZN(n691) );
  NAND2_X1 U515 ( .A1(n561), .A2(G234), .ZN(n413) );
  XNOR2_X1 U516 ( .A(n413), .B(KEYINPUT20), .ZN(n469) );
  NAND2_X1 U517 ( .A1(G221), .A2(n469), .ZN(n414) );
  XOR2_X1 U518 ( .A(KEYINPUT21), .B(n414), .Z(n674) );
  INV_X1 U519 ( .A(n674), .ZN(n505) );
  NOR2_X1 U520 ( .A1(n691), .A2(n505), .ZN(n416) );
  INV_X1 U521 ( .A(KEYINPUT101), .ZN(n415) );
  XNOR2_X1 U522 ( .A(n416), .B(n415), .ZN(n448) );
  XNOR2_X1 U523 ( .A(n417), .B(n418), .ZN(n420) );
  XNOR2_X1 U524 ( .A(n419), .B(G107), .ZN(n455) );
  XNOR2_X1 U525 ( .A(n420), .B(n455), .ZN(n425) );
  XNOR2_X1 U526 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U527 ( .A(n424), .B(n423), .ZN(n479) );
  XNOR2_X1 U528 ( .A(n479), .B(n425), .ZN(n637) );
  NAND2_X1 U529 ( .A1(n729), .A2(G224), .ZN(n426) );
  XNOR2_X1 U530 ( .A(n427), .B(n426), .ZN(n429) );
  XNOR2_X1 U531 ( .A(n428), .B(n429), .ZN(n433) );
  XNOR2_X1 U532 ( .A(KEYINPUT79), .B(KEYINPUT4), .ZN(n430) );
  XNOR2_X1 U533 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U534 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U535 ( .A(n637), .B(n434), .ZN(n619) );
  INV_X1 U536 ( .A(n561), .ZN(n604) );
  XNOR2_X1 U537 ( .A(KEYINPUT74), .B(n396), .ZN(n438) );
  NAND2_X1 U538 ( .A1(n438), .A2(G210), .ZN(n435) );
  XNOR2_X1 U539 ( .A(n435), .B(KEYINPUT81), .ZN(n436) );
  XNOR2_X2 U540 ( .A(n437), .B(n436), .ZN(n554) );
  NAND2_X1 U541 ( .A1(n438), .A2(G214), .ZN(n689) );
  NAND2_X1 U542 ( .A1(n554), .A2(n689), .ZN(n441) );
  INV_X1 U543 ( .A(KEYINPUT78), .ZN(n439) );
  XNOR2_X1 U544 ( .A(n439), .B(KEYINPUT19), .ZN(n440) );
  NOR2_X1 U545 ( .A1(G898), .A2(n729), .ZN(n442) );
  XOR2_X1 U546 ( .A(KEYINPUT93), .B(n442), .Z(n636) );
  NAND2_X1 U547 ( .A1(n636), .A2(G902), .ZN(n443) );
  NAND2_X1 U548 ( .A1(n729), .A2(G952), .ZN(n499) );
  NAND2_X1 U549 ( .A1(n443), .A2(n499), .ZN(n446) );
  INV_X1 U550 ( .A(KEYINPUT14), .ZN(n444) );
  XNOR2_X1 U551 ( .A(n445), .B(n444), .ZN(n703) );
  INV_X1 U552 ( .A(n703), .ZN(n501) );
  NAND2_X1 U553 ( .A1(n446), .A2(n501), .ZN(n447) );
  INV_X1 U554 ( .A(KEYINPUT22), .ZN(n449) );
  XNOR2_X2 U555 ( .A(n450), .B(n449), .ZN(n572) );
  XNOR2_X1 U556 ( .A(G137), .B(G140), .ZN(n463) );
  NAND2_X1 U557 ( .A1(G227), .A2(n729), .ZN(n453) );
  XNOR2_X1 U558 ( .A(n453), .B(G104), .ZN(n454) );
  XOR2_X1 U559 ( .A(n455), .B(n454), .Z(n457) );
  XNOR2_X2 U560 ( .A(n459), .B(G469), .ZN(n582) );
  XOR2_X1 U561 ( .A(KEYINPUT23), .B(G110), .Z(n461) );
  XNOR2_X1 U562 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U563 ( .A(n462), .B(KEYINPUT24), .Z(n466) );
  INV_X1 U564 ( .A(n463), .ZN(n464) );
  XNOR2_X1 U565 ( .A(n466), .B(n465), .ZN(n468) );
  NAND2_X1 U566 ( .A1(n469), .A2(G217), .ZN(n470) );
  NOR2_X1 U567 ( .A1(n672), .A2(n359), .ZN(n487) );
  NAND2_X1 U568 ( .A1(n472), .A2(G210), .ZN(n473) );
  XNOR2_X1 U569 ( .A(n474), .B(n473), .ZN(n478) );
  INV_X1 U570 ( .A(n479), .ZN(n480) );
  XNOR2_X2 U571 ( .A(n485), .B(G472), .ZN(n513) );
  XNOR2_X1 U572 ( .A(n513), .B(KEYINPUT6), .ZN(n569) );
  XNOR2_X1 U573 ( .A(n569), .B(KEYINPUT80), .ZN(n486) );
  XNOR2_X1 U574 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n488) );
  XNOR2_X1 U575 ( .A(G119), .B(KEYINPUT126), .ZN(n489) );
  XNOR2_X1 U576 ( .A(n566), .B(n489), .ZN(G21) );
  NAND2_X1 U577 ( .A1(n675), .A2(n674), .ZN(n671) );
  INV_X1 U578 ( .A(KEYINPUT33), .ZN(n490) );
  INV_X1 U579 ( .A(n584), .ZN(n491) );
  INV_X1 U580 ( .A(KEYINPUT34), .ZN(n492) );
  XNOR2_X1 U581 ( .A(n493), .B(n492), .ZN(n494) );
  AND2_X1 U582 ( .A1(n523), .A2(n348), .ZN(n506) );
  NAND2_X1 U583 ( .A1(n494), .A2(n506), .ZN(n496) );
  XNOR2_X1 U584 ( .A(KEYINPUT87), .B(KEYINPUT35), .ZN(n495) );
  XNOR2_X1 U585 ( .A(n496), .B(n495), .ZN(n568) );
  XNOR2_X1 U586 ( .A(n568), .B(G122), .ZN(G24) );
  NAND2_X1 U587 ( .A1(n513), .A2(n689), .ZN(n497) );
  NOR2_X1 U588 ( .A1(G900), .A2(n729), .ZN(n498) );
  NAND2_X1 U589 ( .A1(n498), .A2(G902), .ZN(n500) );
  NAND2_X1 U590 ( .A1(n500), .A2(n499), .ZN(n502) );
  NAND2_X1 U591 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U592 ( .A(KEYINPUT82), .B(n503), .ZN(n504) );
  NOR2_X1 U593 ( .A1(n505), .A2(n504), .ZN(n510) );
  NAND2_X1 U594 ( .A1(n506), .A2(n554), .ZN(n507) );
  OR2_X1 U595 ( .A1(n507), .A2(n582), .ZN(n508) );
  XNOR2_X1 U596 ( .A(n531), .B(n509), .ZN(G45) );
  INV_X1 U597 ( .A(n675), .ZN(n512) );
  XNOR2_X1 U598 ( .A(KEYINPUT68), .B(n510), .ZN(n511) );
  NAND2_X1 U599 ( .A1(n512), .A2(n511), .ZN(n544) );
  BUF_X2 U600 ( .A(n513), .Z(n580) );
  INV_X1 U601 ( .A(n580), .ZN(n677) );
  XNOR2_X1 U602 ( .A(n514), .B(KEYINPUT28), .ZN(n527) );
  XOR2_X1 U603 ( .A(n582), .B(KEYINPUT106), .Z(n526) );
  NAND2_X1 U604 ( .A1(n527), .A2(n526), .ZN(n538) );
  NOR2_X1 U605 ( .A1(n691), .A2(n692), .ZN(n515) );
  XNOR2_X1 U606 ( .A(KEYINPUT41), .B(n515), .ZN(n687) );
  NOR2_X1 U607 ( .A1(n538), .A2(n687), .ZN(n516) );
  XNOR2_X1 U608 ( .A(n516), .B(KEYINPUT42), .ZN(n741) );
  OR2_X1 U609 ( .A1(n517), .A2(n582), .ZN(n518) );
  NOR2_X1 U610 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U611 ( .A(n520), .B(KEYINPUT39), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n523), .A2(n522), .ZN(n543) );
  INV_X1 U613 ( .A(n523), .ZN(n524) );
  NOR2_X1 U614 ( .A1(n693), .A2(n537), .ZN(n529) );
  AND2_X1 U615 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U616 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U617 ( .A1(n530), .A2(KEYINPUT47), .ZN(n533) );
  XNOR2_X1 U618 ( .A(n531), .B(KEYINPUT85), .ZN(n532) );
  NAND2_X1 U619 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U620 ( .A(n534), .B(KEYINPUT84), .ZN(n541) );
  NOR2_X1 U621 ( .A1(n693), .A2(KEYINPUT47), .ZN(n536) );
  OR2_X1 U622 ( .A1(n538), .A2(n537), .ZN(n647) );
  NOR2_X1 U623 ( .A1(n539), .A2(n647), .ZN(n540) );
  NOR2_X1 U624 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U625 ( .A(n542), .B(KEYINPUT71), .ZN(n550) );
  XNOR2_X1 U626 ( .A(n543), .B(KEYINPUT103), .ZN(n654) );
  INV_X1 U627 ( .A(n654), .ZN(n547) );
  NOR2_X1 U628 ( .A1(n569), .A2(n544), .ZN(n545) );
  XNOR2_X1 U629 ( .A(n545), .B(KEYINPUT104), .ZN(n546) );
  NOR2_X1 U630 ( .A1(n672), .A2(n549), .ZN(n659) );
  NOR2_X1 U631 ( .A1(n550), .A2(n659), .ZN(n551) );
  AND2_X1 U632 ( .A1(n672), .A2(n552), .ZN(n553) );
  XNOR2_X1 U633 ( .A(n553), .B(KEYINPUT43), .ZN(n555) );
  NOR2_X1 U634 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U635 ( .A(n556), .B(KEYINPUT105), .ZN(n737) );
  NOR2_X1 U636 ( .A1(n558), .A2(n557), .ZN(n662) );
  INV_X1 U637 ( .A(KEYINPUT77), .ZN(n560) );
  NOR2_X1 U638 ( .A1(n580), .A2(n359), .ZN(n563) );
  AND2_X1 U639 ( .A1(n672), .A2(n563), .ZN(n564) );
  AND2_X1 U640 ( .A1(n572), .A2(n564), .ZN(n646) );
  INV_X1 U641 ( .A(n646), .ZN(n565) );
  NAND2_X1 U642 ( .A1(n568), .A2(n567), .ZN(n591) );
  NAND2_X1 U643 ( .A1(n591), .A2(KEYINPUT44), .ZN(n589) );
  AND2_X1 U644 ( .A1(n569), .A2(n359), .ZN(n570) );
  AND2_X1 U645 ( .A1(n672), .A2(n570), .ZN(n571) );
  NAND2_X1 U646 ( .A1(n572), .A2(n571), .ZN(n574) );
  INV_X1 U647 ( .A(KEYINPUT102), .ZN(n573) );
  XNOR2_X1 U648 ( .A(n574), .B(n573), .ZN(n742) );
  INV_X1 U649 ( .A(n575), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n580), .A2(n576), .ZN(n682) );
  INV_X1 U651 ( .A(n682), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n584), .A2(n577), .ZN(n579) );
  XNOR2_X1 U653 ( .A(KEYINPUT94), .B(KEYINPUT31), .ZN(n578) );
  XNOR2_X1 U654 ( .A(n579), .B(n578), .ZN(n657) );
  OR2_X1 U655 ( .A1(n580), .A2(n671), .ZN(n581) );
  NOR2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  AND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n641) );
  OR2_X1 U658 ( .A1(n657), .A2(n641), .ZN(n585) );
  XNOR2_X1 U659 ( .A(n585), .B(KEYINPUT95), .ZN(n586) );
  NOR2_X1 U660 ( .A1(n742), .A2(n587), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n590), .B(KEYINPUT89), .ZN(n595) );
  INV_X1 U663 ( .A(n591), .ZN(n593) );
  INV_X1 U664 ( .A(KEYINPUT44), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U667 ( .A(KEYINPUT86), .ZN(n598) );
  XNOR2_X1 U668 ( .A(n599), .B(n598), .ZN(n603) );
  NAND2_X1 U669 ( .A1(n665), .A2(KEYINPUT2), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U671 ( .A1(n604), .A2(KEYINPUT2), .ZN(n605) );
  NAND2_X1 U672 ( .A1(n710), .A2(G472), .ZN(n610) );
  XOR2_X1 U673 ( .A(KEYINPUT62), .B(n608), .Z(n609) );
  XNOR2_X1 U674 ( .A(n610), .B(n609), .ZN(n614) );
  INV_X1 U675 ( .A(G952), .ZN(n611) );
  NAND2_X1 U676 ( .A1(n611), .A2(G953), .ZN(n613) );
  INV_X1 U677 ( .A(KEYINPUT92), .ZN(n612) );
  NOR2_X2 U678 ( .A1(n614), .A2(n723), .ZN(n616) );
  XOR2_X1 U679 ( .A(KEYINPUT108), .B(KEYINPUT63), .Z(n615) );
  XNOR2_X1 U680 ( .A(n616), .B(n615), .ZN(G57) );
  NAND2_X1 U681 ( .A1(n710), .A2(G210), .ZN(n621) );
  XNOR2_X1 U682 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n617) );
  XNOR2_X1 U683 ( .A(n617), .B(KEYINPUT55), .ZN(n618) );
  XNOR2_X1 U684 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U685 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X2 U686 ( .A1(n622), .A2(n723), .ZN(n624) );
  XNOR2_X1 U687 ( .A(KEYINPUT88), .B(KEYINPUT56), .ZN(n623) );
  XNOR2_X1 U688 ( .A(n624), .B(n623), .ZN(G51) );
  NAND2_X1 U689 ( .A1(n710), .A2(G475), .ZN(n628) );
  XNOR2_X1 U690 ( .A(KEYINPUT65), .B(KEYINPUT59), .ZN(n626) );
  XNOR2_X1 U691 ( .A(n625), .B(n626), .ZN(n627) );
  XNOR2_X1 U692 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X2 U693 ( .A1(n629), .A2(n723), .ZN(n630) );
  XNOR2_X1 U694 ( .A(n630), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U695 ( .A(n631), .B(KEYINPUT122), .ZN(n635) );
  NAND2_X1 U696 ( .A1(G953), .A2(G224), .ZN(n632) );
  XNOR2_X1 U697 ( .A(KEYINPUT61), .B(n632), .ZN(n633) );
  NAND2_X1 U698 ( .A1(n633), .A2(G898), .ZN(n634) );
  NAND2_X1 U699 ( .A1(n635), .A2(n634), .ZN(n639) );
  NOR2_X1 U700 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U701 ( .A(n639), .B(n638), .ZN(G69) );
  NAND2_X1 U702 ( .A1(n654), .A2(n641), .ZN(n640) );
  XNOR2_X1 U703 ( .A(n640), .B(G104), .ZN(G6) );
  XOR2_X1 U704 ( .A(KEYINPUT109), .B(KEYINPUT26), .Z(n643) );
  NAND2_X1 U705 ( .A1(n641), .A2(n656), .ZN(n642) );
  XNOR2_X1 U706 ( .A(n643), .B(n642), .ZN(n645) );
  XOR2_X1 U707 ( .A(G107), .B(KEYINPUT27), .Z(n644) );
  XNOR2_X1 U708 ( .A(n645), .B(n644), .ZN(G9) );
  XOR2_X1 U709 ( .A(G110), .B(n646), .Z(G12) );
  XOR2_X1 U710 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n649) );
  INV_X1 U711 ( .A(n647), .ZN(n651) );
  NAND2_X1 U712 ( .A1(n656), .A2(n651), .ZN(n648) );
  XNOR2_X1 U713 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U714 ( .A(G128), .B(n650), .ZN(G30) );
  XOR2_X1 U715 ( .A(G146), .B(KEYINPUT111), .Z(n653) );
  NAND2_X1 U716 ( .A1(n651), .A2(n654), .ZN(n652) );
  XNOR2_X1 U717 ( .A(n653), .B(n652), .ZN(G48) );
  NAND2_X1 U718 ( .A1(n657), .A2(n654), .ZN(n655) );
  XNOR2_X1 U719 ( .A(n655), .B(G113), .ZN(G15) );
  NAND2_X1 U720 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U721 ( .A(n658), .B(G116), .ZN(G18) );
  XNOR2_X1 U722 ( .A(n659), .B(KEYINPUT37), .ZN(n660) );
  XNOR2_X1 U723 ( .A(n660), .B(KEYINPUT112), .ZN(n661) );
  XNOR2_X1 U724 ( .A(G125), .B(n661), .ZN(G27) );
  XNOR2_X1 U725 ( .A(G134), .B(n662), .ZN(n663) );
  XNOR2_X1 U726 ( .A(n663), .B(KEYINPUT113), .ZN(G36) );
  NAND2_X1 U727 ( .A1(KEYINPUT2), .A2(KEYINPUT83), .ZN(n667) );
  NOR2_X1 U728 ( .A1(KEYINPUT2), .A2(KEYINPUT83), .ZN(n664) );
  XNOR2_X1 U729 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U730 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U731 ( .A1(n668), .A2(n729), .ZN(n708) );
  NOR2_X1 U732 ( .A1(n357), .A2(n687), .ZN(n669) );
  XNOR2_X1 U733 ( .A(n669), .B(KEYINPUT120), .ZN(n705) );
  XNOR2_X1 U734 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n670) );
  XNOR2_X1 U735 ( .A(n670), .B(KEYINPUT51), .ZN(n685) );
  NAND2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U737 ( .A(n673), .B(KEYINPUT50), .ZN(n681) );
  NOR2_X1 U738 ( .A1(n359), .A2(n674), .ZN(n676) );
  XNOR2_X1 U739 ( .A(n676), .B(KEYINPUT49), .ZN(n678) );
  NAND2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U741 ( .A(KEYINPUT115), .B(n679), .ZN(n680) );
  NAND2_X1 U742 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U744 ( .A(n685), .B(n684), .Z(n686) );
  NOR2_X1 U745 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U746 ( .A(KEYINPUT118), .B(n688), .Z(n699) );
  NOR2_X1 U747 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U749 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U750 ( .A1(n696), .A2(n357), .ZN(n697) );
  XNOR2_X1 U751 ( .A(KEYINPUT119), .B(n697), .ZN(n698) );
  NAND2_X1 U752 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U753 ( .A(KEYINPUT52), .B(n700), .ZN(n701) );
  NAND2_X1 U754 ( .A1(n701), .A2(G952), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U756 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U757 ( .A(n706), .B(KEYINPUT121), .ZN(n707) );
  NOR2_X1 U758 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U759 ( .A(KEYINPUT53), .B(n709), .ZN(G75) );
  BUF_X1 U760 ( .A(n710), .Z(n719) );
  NAND2_X1 U761 ( .A1(n719), .A2(G469), .ZN(n714) );
  XOR2_X1 U762 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n711) );
  XNOR2_X1 U763 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U764 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U765 ( .A1(n723), .A2(n715), .ZN(G54) );
  NAND2_X1 U766 ( .A1(n719), .A2(G478), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U768 ( .A1(n723), .A2(n718), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n719), .A2(G217), .ZN(n721) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U771 ( .A1(n723), .A2(n722), .ZN(G66) );
  XOR2_X1 U772 ( .A(n724), .B(n725), .Z(n726) );
  XOR2_X1 U773 ( .A(KEYINPUT123), .B(n726), .Z(n731) );
  XOR2_X1 U774 ( .A(KEYINPUT124), .B(n731), .Z(n727) );
  XOR2_X1 U775 ( .A(n728), .B(n727), .Z(n730) );
  NAND2_X1 U776 ( .A1(n730), .A2(n729), .ZN(n736) );
  XNOR2_X1 U777 ( .A(G227), .B(n731), .ZN(n732) );
  NAND2_X1 U778 ( .A1(n732), .A2(G900), .ZN(n733) );
  XOR2_X1 U779 ( .A(KEYINPUT125), .B(n733), .Z(n734) );
  NAND2_X1 U780 ( .A1(G953), .A2(n734), .ZN(n735) );
  NAND2_X1 U781 ( .A1(n736), .A2(n735), .ZN(G72) );
  XNOR2_X1 U782 ( .A(G140), .B(KEYINPUT114), .ZN(n738) );
  XNOR2_X1 U783 ( .A(n738), .B(n737), .ZN(G42) );
  XNOR2_X1 U784 ( .A(G131), .B(KEYINPUT127), .ZN(n740) );
  XNOR2_X1 U785 ( .A(n740), .B(n739), .ZN(G33) );
  XOR2_X1 U786 ( .A(G137), .B(n741), .Z(G39) );
  XOR2_X1 U787 ( .A(G101), .B(n742), .Z(G3) );
endmodule

