

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744;

  XNOR2_X1 U365 ( .A(n605), .B(n601), .ZN(n733) );
  OR2_X1 U366 ( .A1(n520), .A2(n519), .ZN(n521) );
  OR2_X1 U367 ( .A1(n506), .A2(n492), .ZN(n493) );
  XNOR2_X1 U368 ( .A(n503), .B(KEYINPUT31), .ZN(n668) );
  XNOR2_X1 U369 ( .A(n456), .B(KEYINPUT0), .ZN(n506) );
  OR2_X1 U370 ( .A1(n531), .A2(n681), .ZN(n372) );
  NOR2_X2 U371 ( .A1(n550), .A2(n490), .ZN(n366) );
  XNOR2_X1 U372 ( .A(n732), .B(G146), .ZN(n429) );
  XNOR2_X1 U373 ( .A(n459), .B(n424), .ZN(n731) );
  BUF_X1 U374 ( .A(G143), .Z(n343) );
  INV_X1 U375 ( .A(G143), .ZN(n370) );
  NOR2_X2 U376 ( .A1(n563), .A2(n682), .ZN(n543) );
  XNOR2_X2 U377 ( .A(n540), .B(KEYINPUT76), .ZN(n563) );
  AND2_X2 U378 ( .A1(n733), .A2(n604), .ZN(n345) );
  AND2_X2 U379 ( .A1(n631), .A2(n483), .ZN(n401) );
  XNOR2_X1 U380 ( .A(n576), .B(n449), .ZN(n580) );
  XOR2_X1 U381 ( .A(n443), .B(n442), .Z(n344) );
  OR2_X1 U382 ( .A1(n506), .A2(n689), .ZN(n503) );
  XNOR2_X2 U383 ( .A(n474), .B(n369), .ZN(n443) );
  XNOR2_X1 U384 ( .A(n436), .B(n355), .ZN(n356) );
  AND2_X1 U385 ( .A1(n518), .A2(n515), .ZN(n516) );
  OR2_X1 U386 ( .A1(n742), .A2(n488), .ZN(n498) );
  XNOR2_X1 U387 ( .A(n487), .B(n486), .ZN(n742) );
  XNOR2_X1 U388 ( .A(n432), .B(n431), .ZN(n715) );
  XNOR2_X1 U389 ( .A(n570), .B(KEYINPUT105), .ZN(n665) );
  OR2_X1 U390 ( .A1(n551), .A2(n502), .ZN(n689) );
  XNOR2_X1 U391 ( .A(n430), .B(G469), .ZN(n553) );
  XNOR2_X1 U392 ( .A(n443), .B(n368), .ZN(n732) );
  XNOR2_X1 U393 ( .A(G101), .B(KEYINPUT75), .ZN(n373) );
  NOR2_X2 U394 ( .A1(n653), .A2(n510), .ZN(n518) );
  NOR2_X1 U395 ( .A1(n715), .A2(n506), .ZN(n457) );
  XNOR2_X1 U396 ( .A(n372), .B(n371), .ZN(n539) );
  XNOR2_X2 U397 ( .A(n598), .B(n542), .ZN(n682) );
  NAND2_X1 U398 ( .A1(n528), .A2(n527), .ZN(n530) );
  INV_X1 U399 ( .A(G237), .ZN(n444) );
  XNOR2_X1 U400 ( .A(n553), .B(KEYINPUT1), .ZN(n494) );
  AND2_X1 U401 ( .A1(n348), .A2(n604), .ZN(n677) );
  AND2_X1 U402 ( .A1(n352), .A2(n680), .ZN(n510) );
  INV_X1 U403 ( .A(n349), .ZN(n354) );
  XNOR2_X1 U404 ( .A(n401), .B(G472), .ZN(n531) );
  XNOR2_X1 U405 ( .A(G101), .B(G137), .ZN(n391) );
  XOR2_X1 U406 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n392) );
  NOR2_X1 U407 ( .A1(G953), .A2(G237), .ZN(n461) );
  XNOR2_X1 U408 ( .A(n367), .B(n440), .ZN(n459) );
  XNOR2_X1 U409 ( .A(n351), .B(KEYINPUT69), .ZN(n403) );
  INV_X1 U410 ( .A(KEYINPUT10), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n458), .B(G134), .ZN(n368) );
  XNOR2_X1 U412 ( .A(G137), .B(KEYINPUT71), .ZN(n424) );
  OR2_X1 U413 ( .A1(n648), .A2(G902), .ZN(n430) );
  XNOR2_X1 U414 ( .A(n399), .B(n398), .ZN(n435) );
  XNOR2_X1 U415 ( .A(G119), .B(G116), .ZN(n396) );
  XNOR2_X1 U416 ( .A(KEYINPUT24), .B(KEYINPUT96), .ZN(n404) );
  XNOR2_X1 U417 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U418 ( .A(G128), .B(G119), .ZN(n407) );
  XOR2_X1 U419 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n411) );
  XNOR2_X1 U420 ( .A(n423), .B(n422), .ZN(n434) );
  XNOR2_X1 U421 ( .A(KEYINPUT90), .B(G110), .ZN(n422) );
  XNOR2_X1 U422 ( .A(n374), .B(n373), .ZN(n423) );
  XNOR2_X1 U423 ( .A(G107), .B(G104), .ZN(n374) );
  XNOR2_X1 U424 ( .A(n356), .B(n344), .ZN(n610) );
  BUF_X1 U425 ( .A(n541), .Z(n598) );
  NAND2_X1 U426 ( .A1(n375), .A2(n595), .ZN(n576) );
  BUF_X1 U427 ( .A(n494), .Z(n690) );
  XNOR2_X1 U428 ( .A(n493), .B(n350), .ZN(n361) );
  INV_X1 U429 ( .A(n677), .ZN(n606) );
  NAND2_X1 U430 ( .A1(n385), .A2(KEYINPUT81), .ZN(n384) );
  NOR2_X1 U431 ( .A1(n678), .A2(n677), .ZN(n382) );
  INV_X1 U432 ( .A(KEYINPUT82), .ZN(n381) );
  INV_X2 U433 ( .A(G953), .ZN(n737) );
  NAND2_X1 U434 ( .A1(G234), .A2(G237), .ZN(n450) );
  INV_X1 U435 ( .A(KEYINPUT30), .ZN(n371) );
  INV_X1 U436 ( .A(KEYINPUT72), .ZN(n395) );
  XNOR2_X1 U437 ( .A(KEYINPUT70), .B(G131), .ZN(n458) );
  XNOR2_X1 U438 ( .A(n343), .B(G113), .ZN(n466) );
  XOR2_X1 U439 ( .A(G122), .B(G104), .Z(n465) );
  XNOR2_X1 U440 ( .A(n378), .B(G146), .ZN(n440) );
  INV_X1 U441 ( .A(G125), .ZN(n378) );
  XNOR2_X1 U442 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n369) );
  XNOR2_X1 U443 ( .A(n429), .B(n383), .ZN(n631) );
  XNOR2_X1 U444 ( .A(n435), .B(n400), .ZN(n383) );
  INV_X1 U445 ( .A(KEYINPUT81), .ZN(n390) );
  NOR2_X1 U446 ( .A1(n573), .A2(n502), .ZN(n432) );
  XNOR2_X1 U447 ( .A(n357), .B(KEYINPUT41), .ZN(n705) );
  NAND2_X1 U448 ( .A1(n358), .A2(n557), .ZN(n357) );
  XNOR2_X1 U449 ( .A(n473), .B(n472), .ZN(n509) );
  BUF_X1 U450 ( .A(n550), .Z(n694) );
  INV_X1 U451 ( .A(n690), .ZN(n376) );
  INV_X1 U452 ( .A(n435), .ZN(n355) );
  XNOR2_X1 U453 ( .A(n434), .B(n433), .ZN(n436) );
  INV_X1 U454 ( .A(n377), .ZN(n723) );
  BUF_X1 U455 ( .A(n604), .Z(n377) );
  XNOR2_X1 U456 ( .A(n731), .B(n414), .ZN(n637) );
  XNOR2_X1 U457 ( .A(n409), .B(n408), .ZN(n413) );
  AND2_X1 U458 ( .A1(n606), .A2(G475), .ZN(n362) );
  AND2_X1 U459 ( .A1(n607), .A2(n606), .ZN(n645) );
  XNOR2_X1 U460 ( .A(n427), .B(n428), .ZN(n360) );
  AND2_X1 U461 ( .A1(n606), .A2(G210), .ZN(n363) );
  AND2_X1 U462 ( .A1(n578), .A2(n690), .ZN(n672) );
  NAND2_X1 U463 ( .A1(n607), .A2(n346), .ZN(n642) );
  AND2_X1 U464 ( .A1(n380), .A2(n379), .ZN(n720) );
  AND2_X1 U465 ( .A1(n719), .A2(n737), .ZN(n379) );
  XNOR2_X1 U466 ( .A(n382), .B(n381), .ZN(n380) );
  AND2_X1 U467 ( .A1(n606), .A2(G478), .ZN(n346) );
  AND2_X1 U468 ( .A1(n573), .A2(n511), .ZN(n347) );
  AND2_X1 U469 ( .A1(n605), .A2(KEYINPUT2), .ZN(n348) );
  NOR2_X1 U470 ( .A1(n506), .A2(n505), .ZN(n349) );
  XOR2_X1 U471 ( .A(KEYINPUT66), .B(KEYINPUT22), .Z(n350) );
  NAND2_X1 U472 ( .A1(n353), .A2(n354), .ZN(n352) );
  INV_X1 U473 ( .A(n668), .ZN(n353) );
  XNOR2_X1 U474 ( .A(n356), .B(KEYINPUT125), .ZN(n722) );
  INV_X1 U475 ( .A(n682), .ZN(n358) );
  XNOR2_X1 U476 ( .A(n429), .B(n359), .ZN(n648) );
  XNOR2_X1 U477 ( .A(n360), .B(n434), .ZN(n359) );
  NAND2_X1 U478 ( .A1(n361), .A2(n347), .ZN(n514) );
  NAND2_X1 U479 ( .A1(n361), .A2(n376), .ZN(n501) );
  NAND2_X1 U480 ( .A1(n607), .A2(n362), .ZN(n619) );
  NAND2_X1 U481 ( .A1(n607), .A2(n363), .ZN(n612) );
  NAND2_X1 U482 ( .A1(n607), .A2(n364), .ZN(n633) );
  AND2_X1 U483 ( .A1(n606), .A2(G472), .ZN(n364) );
  NAND2_X1 U484 ( .A1(n365), .A2(n389), .ZN(n388) );
  NAND2_X1 U485 ( .A1(n345), .A2(n390), .ZN(n365) );
  NAND2_X1 U486 ( .A1(n366), .A2(n553), .ZN(n537) );
  NAND2_X1 U487 ( .A1(n494), .A2(n366), .ZN(n502) );
  NOR2_X1 U488 ( .A1(n690), .A2(n366), .ZN(n692) );
  XNOR2_X1 U489 ( .A(n403), .B(G140), .ZN(n367) );
  XNOR2_X2 U490 ( .A(n551), .B(n402), .ZN(n573) );
  XNOR2_X2 U491 ( .A(n370), .B(G128), .ZN(n474) );
  NAND2_X1 U492 ( .A1(n580), .A2(n455), .ZN(n456) );
  INV_X1 U493 ( .A(n541), .ZN(n375) );
  XNOR2_X2 U494 ( .A(n446), .B(n445), .ZN(n541) );
  XNOR2_X2 U495 ( .A(n530), .B(n529), .ZN(n604) );
  NAND2_X2 U496 ( .A1(n387), .A2(n384), .ZN(n607) );
  NAND2_X1 U497 ( .A1(n386), .A2(n604), .ZN(n385) );
  AND2_X1 U498 ( .A1(n733), .A2(n603), .ZN(n386) );
  NAND2_X1 U499 ( .A1(n388), .A2(n603), .ZN(n387) );
  INV_X1 U500 ( .A(KEYINPUT2), .ZN(n389) );
  INV_X1 U501 ( .A(G110), .ZN(n406) );
  XNOR2_X1 U502 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n431) );
  INV_X1 U503 ( .A(KEYINPUT83), .ZN(n601) );
  XNOR2_X1 U504 ( .A(n471), .B(G475), .ZN(n472) );
  BUF_X1 U505 ( .A(n659), .Z(n662) );
  INV_X1 U506 ( .A(KEYINPUT60), .ZN(n621) );
  XNOR2_X1 U507 ( .A(n392), .B(n391), .ZN(n394) );
  AND2_X1 U508 ( .A1(n461), .A2(G210), .ZN(n393) );
  XNOR2_X1 U509 ( .A(n394), .B(n393), .ZN(n400) );
  XNOR2_X1 U510 ( .A(n395), .B(G113), .ZN(n397) );
  XNOR2_X1 U511 ( .A(n397), .B(n396), .ZN(n399) );
  XNOR2_X1 U512 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n398) );
  INV_X1 U513 ( .A(G902), .ZN(n483) );
  INV_X1 U514 ( .A(n531), .ZN(n700) );
  INV_X2 U515 ( .A(n700), .ZN(n551) );
  INV_X1 U516 ( .A(KEYINPUT6), .ZN(n402) );
  XOR2_X1 U517 ( .A(KEYINPUT95), .B(KEYINPUT23), .Z(n405) );
  XNOR2_X1 U518 ( .A(n405), .B(n404), .ZN(n409) );
  NAND2_X1 U519 ( .A1(G234), .A2(n737), .ZN(n410) );
  XNOR2_X1 U520 ( .A(n411), .B(n410), .ZN(n476) );
  NAND2_X1 U521 ( .A1(n476), .A2(G221), .ZN(n412) );
  XNOR2_X1 U522 ( .A(n413), .B(n412), .ZN(n414) );
  NAND2_X1 U523 ( .A1(n637), .A2(n483), .ZN(n418) );
  XNOR2_X1 U524 ( .A(G902), .B(KEYINPUT15), .ZN(n602) );
  NAND2_X1 U525 ( .A1(n602), .A2(G234), .ZN(n415) );
  XNOR2_X1 U526 ( .A(n415), .B(KEYINPUT20), .ZN(n419) );
  NAND2_X1 U527 ( .A1(n419), .A2(G217), .ZN(n416) );
  XNOR2_X1 U528 ( .A(n416), .B(KEYINPUT25), .ZN(n417) );
  XNOR2_X2 U529 ( .A(n418), .B(n417), .ZN(n550) );
  NAND2_X1 U530 ( .A1(n419), .A2(G221), .ZN(n421) );
  XOR2_X1 U531 ( .A(KEYINPUT97), .B(KEYINPUT21), .Z(n420) );
  XNOR2_X1 U532 ( .A(n421), .B(n420), .ZN(n693) );
  XNOR2_X1 U533 ( .A(n693), .B(KEYINPUT98), .ZN(n490) );
  INV_X1 U534 ( .A(n424), .ZN(n426) );
  NAND2_X1 U535 ( .A1(G227), .A2(n737), .ZN(n425) );
  XNOR2_X1 U536 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U537 ( .A(KEYINPUT94), .B(G140), .ZN(n428) );
  XNOR2_X1 U538 ( .A(KEYINPUT16), .B(G122), .ZN(n433) );
  NAND2_X1 U539 ( .A1(n737), .A2(G224), .ZN(n437) );
  XNOR2_X1 U540 ( .A(n437), .B(KEYINPUT91), .ZN(n439) );
  XNOR2_X1 U541 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n438) );
  XNOR2_X1 U542 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U543 ( .A(n441), .B(n440), .ZN(n442) );
  NAND2_X1 U544 ( .A1(n610), .A2(n602), .ZN(n446) );
  NAND2_X1 U545 ( .A1(n483), .A2(n444), .ZN(n447) );
  NAND2_X1 U546 ( .A1(n447), .A2(G210), .ZN(n445) );
  NAND2_X1 U547 ( .A1(n447), .A2(G214), .ZN(n595) );
  INV_X1 U548 ( .A(n595), .ZN(n681) );
  INV_X1 U549 ( .A(KEYINPUT67), .ZN(n448) );
  XNOR2_X1 U550 ( .A(n448), .B(KEYINPUT19), .ZN(n449) );
  XNOR2_X1 U551 ( .A(n450), .B(KEYINPUT14), .ZN(n451) );
  NAND2_X1 U552 ( .A1(G952), .A2(n451), .ZN(n712) );
  NOR2_X1 U553 ( .A1(n712), .A2(G953), .ZN(n535) );
  INV_X1 U554 ( .A(n535), .ZN(n454) );
  NAND2_X1 U555 ( .A1(G902), .A2(n451), .ZN(n532) );
  XOR2_X1 U556 ( .A(G898), .B(KEYINPUT92), .Z(n726) );
  NAND2_X1 U557 ( .A1(G953), .A2(n726), .ZN(n721) );
  NOR2_X1 U558 ( .A1(n532), .A2(n721), .ZN(n452) );
  XNOR2_X1 U559 ( .A(n452), .B(KEYINPUT93), .ZN(n453) );
  NAND2_X1 U560 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U561 ( .A(n457), .B(KEYINPUT34), .ZN(n485) );
  INV_X1 U562 ( .A(n458), .ZN(n460) );
  XNOR2_X1 U563 ( .A(n460), .B(n459), .ZN(n470) );
  XOR2_X1 U564 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n463) );
  NAND2_X1 U565 ( .A1(G214), .A2(n461), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U567 ( .A(n464), .B(KEYINPUT100), .Z(n468) );
  XNOR2_X1 U568 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U569 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U570 ( .A(n470), .B(n469), .ZN(n617) );
  NOR2_X1 U571 ( .A1(G902), .A2(n617), .ZN(n473) );
  XNOR2_X1 U572 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n474), .B(G134), .ZN(n475) );
  XNOR2_X1 U574 ( .A(n475), .B(G107), .ZN(n482) );
  XNOR2_X1 U575 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n480) );
  XNOR2_X1 U576 ( .A(G116), .B(G122), .ZN(n478) );
  NAND2_X1 U577 ( .A1(G217), .A2(n476), .ZN(n477) );
  XNOR2_X1 U578 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U579 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U580 ( .A(n482), .B(n481), .ZN(n643) );
  NAND2_X1 U581 ( .A1(n643), .A2(n483), .ZN(n484) );
  XNOR2_X1 U582 ( .A(n484), .B(G478), .ZN(n508) );
  INV_X1 U583 ( .A(n508), .ZN(n489) );
  NOR2_X1 U584 ( .A1(n509), .A2(n489), .ZN(n565) );
  NAND2_X1 U585 ( .A1(n485), .A2(n565), .ZN(n487) );
  INV_X1 U586 ( .A(KEYINPUT35), .ZN(n486) );
  INV_X1 U587 ( .A(KEYINPUT86), .ZN(n488) );
  AND2_X1 U588 ( .A1(n509), .A2(n489), .ZN(n683) );
  INV_X1 U589 ( .A(n490), .ZN(n491) );
  NAND2_X1 U590 ( .A1(n683), .A2(n491), .ZN(n492) );
  INV_X1 U591 ( .A(KEYINPUT104), .ZN(n495) );
  XNOR2_X1 U592 ( .A(n501), .B(n495), .ZN(n497) );
  AND2_X1 U593 ( .A1(n551), .A2(n694), .ZN(n496) );
  NAND2_X1 U594 ( .A1(n497), .A2(n496), .ZN(n628) );
  AND2_X1 U595 ( .A1(n498), .A2(n628), .ZN(n517) );
  INV_X1 U596 ( .A(n694), .ZN(n499) );
  NAND2_X1 U597 ( .A1(n573), .A2(n499), .ZN(n500) );
  NOR2_X1 U598 ( .A1(n501), .A2(n500), .ZN(n653) );
  INV_X1 U599 ( .A(n537), .ZN(n504) );
  NAND2_X1 U600 ( .A1(n551), .A2(n504), .ZN(n505) );
  NAND2_X1 U601 ( .A1(n508), .A2(n509), .ZN(n507) );
  XOR2_X1 U602 ( .A(KEYINPUT102), .B(n507), .Z(n669) );
  XNOR2_X1 U603 ( .A(n669), .B(KEYINPUT103), .ZN(n591) );
  OR2_X1 U604 ( .A1(n509), .A2(n508), .ZN(n570) );
  NAND2_X1 U605 ( .A1(n591), .A2(n570), .ZN(n680) );
  AND2_X1 U606 ( .A1(n694), .A2(n690), .ZN(n511) );
  INV_X1 U607 ( .A(KEYINPUT77), .ZN(n512) );
  XNOR2_X1 U608 ( .A(n512), .B(KEYINPUT32), .ZN(n513) );
  XNOR2_X2 U609 ( .A(n514), .B(n513), .ZN(n626) );
  AND2_X1 U610 ( .A1(n626), .A2(KEYINPUT44), .ZN(n515) );
  NAND2_X1 U611 ( .A1(n517), .A2(n516), .ZN(n522) );
  INV_X1 U612 ( .A(n518), .ZN(n520) );
  INV_X1 U613 ( .A(KEYINPUT44), .ZN(n523) );
  NAND2_X1 U614 ( .A1(n523), .A2(KEYINPUT86), .ZN(n519) );
  NAND2_X1 U615 ( .A1(n522), .A2(n521), .ZN(n528) );
  AND2_X1 U616 ( .A1(n626), .A2(n523), .ZN(n524) );
  NAND2_X1 U617 ( .A1(n524), .A2(n628), .ZN(n525) );
  NAND2_X1 U618 ( .A1(n525), .A2(KEYINPUT86), .ZN(n526) );
  NAND2_X1 U619 ( .A1(n526), .A2(n742), .ZN(n527) );
  XNOR2_X1 U620 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n529) );
  OR2_X1 U621 ( .A1(n737), .A2(n532), .ZN(n533) );
  NOR2_X1 U622 ( .A1(G900), .A2(n533), .ZN(n534) );
  NOR2_X1 U623 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U624 ( .A(KEYINPUT79), .B(n536), .Z(n548) );
  NOR2_X1 U625 ( .A1(n537), .A2(n548), .ZN(n538) );
  NAND2_X1 U626 ( .A1(n539), .A2(n538), .ZN(n540) );
  INV_X1 U627 ( .A(KEYINPUT38), .ZN(n542) );
  XNOR2_X1 U628 ( .A(n543), .B(KEYINPUT39), .ZN(n592) );
  INV_X1 U629 ( .A(n592), .ZN(n545) );
  INV_X1 U630 ( .A(n570), .ZN(n544) );
  NAND2_X1 U631 ( .A1(n545), .A2(n544), .ZN(n547) );
  INV_X1 U632 ( .A(KEYINPUT40), .ZN(n546) );
  XNOR2_X1 U633 ( .A(n547), .B(n546), .ZN(n743) );
  NOR2_X1 U634 ( .A1(n693), .A2(n548), .ZN(n549) );
  NAND2_X1 U635 ( .A1(n550), .A2(n549), .ZN(n572) );
  NOR2_X1 U636 ( .A1(n572), .A2(n551), .ZN(n552) );
  XNOR2_X1 U637 ( .A(KEYINPUT28), .B(n552), .ZN(n554) );
  AND2_X1 U638 ( .A1(n554), .A2(n553), .ZN(n556) );
  INV_X1 U639 ( .A(KEYINPUT107), .ZN(n555) );
  XNOR2_X1 U640 ( .A(n556), .B(n555), .ZN(n581) );
  AND2_X1 U641 ( .A1(n683), .A2(n595), .ZN(n557) );
  NAND2_X1 U642 ( .A1(n581), .A2(n705), .ZN(n560) );
  INV_X1 U643 ( .A(KEYINPUT108), .ZN(n558) );
  XNOR2_X1 U644 ( .A(n558), .B(KEYINPUT42), .ZN(n559) );
  XNOR2_X1 U645 ( .A(n560), .B(n559), .ZN(n623) );
  NOR2_X1 U646 ( .A1(n743), .A2(n623), .ZN(n562) );
  XOR2_X1 U647 ( .A(KEYINPUT85), .B(KEYINPUT46), .Z(n561) );
  XNOR2_X1 U648 ( .A(n562), .B(n561), .ZN(n588) );
  BUF_X1 U649 ( .A(n563), .Z(n567) );
  INV_X1 U650 ( .A(n598), .ZN(n564) );
  NAND2_X1 U651 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U652 ( .A1(n567), .A2(n566), .ZN(n569) );
  INV_X1 U653 ( .A(KEYINPUT106), .ZN(n568) );
  XNOR2_X1 U654 ( .A(n569), .B(n568), .ZN(n744) );
  INV_X1 U655 ( .A(n665), .ZN(n571) );
  NOR2_X1 U656 ( .A1(n572), .A2(n571), .ZN(n575) );
  INV_X1 U657 ( .A(n573), .ZN(n574) );
  NAND2_X1 U658 ( .A1(n575), .A2(n574), .ZN(n593) );
  NOR2_X1 U659 ( .A1(n593), .A2(n576), .ZN(n577) );
  XNOR2_X1 U660 ( .A(n577), .B(KEYINPUT36), .ZN(n578) );
  INV_X1 U661 ( .A(n672), .ZN(n579) );
  NAND2_X1 U662 ( .A1(n744), .A2(n579), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n581), .A2(n580), .ZN(n583) );
  INV_X1 U664 ( .A(KEYINPUT78), .ZN(n582) );
  XNOR2_X2 U665 ( .A(n583), .B(n582), .ZN(n659) );
  NAND2_X1 U666 ( .A1(n659), .A2(n680), .ZN(n584) );
  XNOR2_X1 U667 ( .A(n584), .B(KEYINPUT47), .ZN(n585) );
  NOR2_X1 U668 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U669 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U670 ( .A(KEYINPUT84), .B(KEYINPUT48), .ZN(n589) );
  XNOR2_X1 U671 ( .A(n590), .B(n589), .ZN(n600) );
  OR2_X1 U672 ( .A1(n592), .A2(n591), .ZN(n674) );
  NOR2_X1 U673 ( .A1(n690), .A2(n593), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT43), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n625) );
  NAND2_X1 U677 ( .A1(n674), .A2(n625), .ZN(n599) );
  NOR2_X2 U678 ( .A1(n600), .A2(n599), .ZN(n605) );
  INV_X1 U679 ( .A(n602), .ZN(n603) );
  XNOR2_X1 U680 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n608), .B(KEYINPUT55), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n612), .B(n611), .ZN(n614) );
  NOR2_X1 U684 ( .A1(n737), .A2(G952), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n613), .B(KEYINPUT89), .ZN(n640) );
  NAND2_X1 U686 ( .A1(n614), .A2(n640), .ZN(n616) );
  INV_X1 U687 ( .A(KEYINPUT56), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(G51) );
  XNOR2_X1 U689 ( .A(n617), .B(KEYINPUT59), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n620), .A2(n640), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(G60) );
  XOR2_X1 U693 ( .A(G137), .B(n623), .Z(G39) );
  XOR2_X1 U694 ( .A(G140), .B(KEYINPUT115), .Z(n624) );
  XNOR2_X1 U695 ( .A(n625), .B(n624), .ZN(G42) );
  XNOR2_X1 U696 ( .A(G119), .B(KEYINPUT127), .ZN(n627) );
  XOR2_X1 U697 ( .A(n627), .B(n626), .Z(G21) );
  XNOR2_X1 U698 ( .A(n628), .B(G110), .ZN(G12) );
  XOR2_X1 U699 ( .A(KEYINPUT88), .B(KEYINPUT109), .Z(n629) );
  XNOR2_X1 U700 ( .A(n629), .B(KEYINPUT62), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U702 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n634), .A2(n640), .ZN(n636) );
  XNOR2_X1 U704 ( .A(KEYINPUT110), .B(KEYINPUT63), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(G57) );
  NAND2_X1 U706 ( .A1(n645), .A2(G217), .ZN(n639) );
  XOR2_X1 U707 ( .A(KEYINPUT124), .B(n637), .Z(n638) );
  XNOR2_X1 U708 ( .A(n639), .B(n638), .ZN(n641) );
  INV_X1 U709 ( .A(n640), .ZN(n651) );
  NOR2_X1 U710 ( .A1(n641), .A2(n651), .ZN(G66) );
  XOR2_X1 U711 ( .A(n643), .B(n642), .Z(n644) );
  NOR2_X1 U712 ( .A1(n644), .A2(n651), .ZN(G63) );
  NAND2_X1 U713 ( .A1(n645), .A2(G469), .ZN(n650) );
  XNOR2_X1 U714 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n646), .B(KEYINPUT58), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U717 ( .A(n650), .B(n649), .ZN(n652) );
  NOR2_X1 U718 ( .A1(n652), .A2(n651), .ZN(G54) );
  XOR2_X1 U719 ( .A(G101), .B(n653), .Z(G3) );
  XOR2_X1 U720 ( .A(G104), .B(KEYINPUT111), .Z(n655) );
  NAND2_X1 U721 ( .A1(n349), .A2(n665), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n655), .B(n654), .ZN(G6) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n657) );
  NAND2_X1 U724 ( .A1(n349), .A2(n669), .ZN(n656) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U726 ( .A(G107), .B(n658), .ZN(G9) );
  XOR2_X1 U727 ( .A(G128), .B(KEYINPUT29), .Z(n661) );
  NAND2_X1 U728 ( .A1(n669), .A2(n662), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n661), .B(n660), .ZN(G30) );
  NAND2_X1 U730 ( .A1(n662), .A2(n665), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n663), .B(KEYINPUT112), .ZN(n664) );
  XNOR2_X1 U732 ( .A(G146), .B(n664), .ZN(G48) );
  XOR2_X1 U733 ( .A(G113), .B(KEYINPUT113), .Z(n667) );
  NAND2_X1 U734 ( .A1(n668), .A2(n665), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n667), .B(n666), .ZN(G15) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n670), .B(KEYINPUT114), .ZN(n671) );
  XNOR2_X1 U738 ( .A(G116), .B(n671), .ZN(G18) );
  XNOR2_X1 U739 ( .A(G125), .B(n672), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n673), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U741 ( .A(n674), .ZN(n675) );
  XOR2_X1 U742 ( .A(G134), .B(n675), .Z(G36) );
  XNOR2_X1 U743 ( .A(KEYINPUT80), .B(KEYINPUT2), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n345), .A2(n676), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n682), .A2(n681), .ZN(n679) );
  NAND2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n686) );
  NAND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n684) );
  NAND2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  AND2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n715), .A2(n687), .ZN(n708) );
  XNOR2_X1 U751 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n688) );
  XNOR2_X1 U752 ( .A(n688), .B(KEYINPUT119), .ZN(n704) );
  INV_X1 U753 ( .A(n689), .ZN(n702) );
  XNOR2_X1 U754 ( .A(KEYINPUT117), .B(KEYINPUT50), .ZN(n691) );
  XNOR2_X1 U755 ( .A(n692), .B(n691), .ZN(n698) );
  XOR2_X1 U756 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n696) );
  NAND2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U758 ( .A(n696), .B(n695), .ZN(n697) );
  NAND2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U761 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U762 ( .A(n704), .B(n703), .ZN(n706) );
  INV_X1 U763 ( .A(n705), .ZN(n714) );
  NOR2_X1 U764 ( .A1(n706), .A2(n714), .ZN(n707) );
  NOR2_X1 U765 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U766 ( .A(n709), .B(KEYINPUT120), .ZN(n710) );
  XNOR2_X1 U767 ( .A(KEYINPUT52), .B(n710), .ZN(n711) );
  NOR2_X1 U768 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U769 ( .A(KEYINPUT121), .B(n713), .Z(n717) );
  NOR2_X1 U770 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U772 ( .A(KEYINPUT122), .B(n718), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U774 ( .A1(n722), .A2(n721), .ZN(n730) );
  NOR2_X1 U775 ( .A1(n723), .A2(G953), .ZN(n728) );
  NAND2_X1 U776 ( .A1(G953), .A2(G224), .ZN(n724) );
  XOR2_X1 U777 ( .A(KEYINPUT61), .B(n724), .Z(n725) );
  NOR2_X1 U778 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U779 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U780 ( .A(n730), .B(n729), .ZN(G69) );
  XOR2_X1 U781 ( .A(n732), .B(n731), .Z(n735) );
  XOR2_X1 U782 ( .A(n735), .B(n733), .Z(n734) );
  NOR2_X1 U783 ( .A1(n734), .A2(G953), .ZN(n740) );
  XNOR2_X1 U784 ( .A(G227), .B(n735), .ZN(n736) );
  NAND2_X1 U785 ( .A1(n736), .A2(G900), .ZN(n738) );
  NOR2_X1 U786 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U787 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U788 ( .A(KEYINPUT126), .B(n741), .ZN(G72) );
  XNOR2_X1 U789 ( .A(G122), .B(n742), .ZN(G24) );
  XOR2_X1 U790 ( .A(n743), .B(G131), .Z(G33) );
  XNOR2_X1 U791 ( .A(n343), .B(n744), .ZN(G45) );
endmodule

