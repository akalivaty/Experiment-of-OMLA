//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n582, new_n583, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n640, new_n641, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  XNOR2_X1  g003(.A(KEYINPUT66), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT67), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n465), .A2(new_n469), .A3(G137), .A4(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n468), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G101), .A3(new_n470), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n463), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n472), .B1(new_n471), .B2(new_n474), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n465), .A2(new_n469), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(new_n470), .ZN(new_n487));
  MUX2_X1   g062(.A(G100), .B(G112), .S(G2105), .Z(new_n488));
  AOI22_X1  g063(.A1(new_n487), .A2(G124), .B1(G2104), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n486), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n489), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT72), .ZN(G162));
  NAND4_X1  g069(.A1(new_n477), .A2(new_n478), .A3(G138), .A4(new_n470), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n465), .A2(new_n469), .A3(G126), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n497), .B1(new_n500), .B2(G2105), .ZN(new_n501));
  NAND2_X1  g076(.A1(G102), .A2(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT4), .A2(G138), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n486), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n470), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(KEYINPUT73), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n508), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(new_n511), .B2(new_n513), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT74), .A3(G50), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT5), .B(G543), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(new_n510), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n512), .A2(KEYINPUT6), .A3(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT6), .B1(new_n512), .B2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n514), .A2(KEYINPUT75), .A3(new_n522), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n521), .B(new_n524), .C1(new_n525), .C2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n515), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n519), .A2(KEYINPUT77), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(KEYINPUT5), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  NAND2_X1  g115(.A1(KEYINPUT5), .A2(G543), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(KEYINPUT5), .A2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(KEYINPUT5), .A2(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT76), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  AND2_X1   g122(.A1(G63), .A2(G651), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n538), .A2(G51), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  XNOR2_X1  g126(.A(KEYINPUT78), .B(G89), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n532), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n553), .A2(KEYINPUT79), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(KEYINPUT79), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n549), .B1(new_n554), .B2(new_n555), .ZN(G286));
  INV_X1    g131(.A(G286), .ZN(G168));
  NAND2_X1  g132(.A1(G77), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G64), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n546), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n510), .B1(new_n560), .B2(KEYINPUT80), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n561), .B1(KEYINPUT80), .B2(new_n560), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n514), .A2(KEYINPUT75), .A3(new_n522), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT75), .B1(new_n514), .B2(new_n522), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(G90), .A2(new_n565), .B1(new_n538), .B2(G52), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G301));
  INV_X1    g142(.A(G301), .ZN(G171));
  AOI22_X1  g143(.A1(new_n547), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n510), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n538), .A2(G43), .ZN(new_n572));
  INV_X1    g147(.A(G81), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n573), .B2(new_n532), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n574), .A2(KEYINPUT81), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(KEYINPUT81), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n571), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G860), .ZN(G153));
  AND3_X1   g154(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G36), .ZN(G176));
  NAND2_X1  g156(.A1(G1), .A2(G3), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT8), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n580), .A2(new_n583), .ZN(G188));
  NAND2_X1  g159(.A1(new_n519), .A2(G53), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT9), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n522), .A2(G65), .ZN(new_n587));
  AND2_X1   g162(.A1(G78), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n565), .A2(G91), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n586), .A2(new_n589), .ZN(new_n594));
  INV_X1    g169(.A(new_n592), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT82), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G299));
  INV_X1    g173(.A(G74), .ZN(new_n599));
  NOR3_X1   g174(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT76), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G49), .B2(new_n519), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n530), .A2(G87), .A3(new_n531), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G288));
  NAND3_X1  g180(.A1(new_n530), .A2(G86), .A3(new_n531), .ZN(new_n606));
  OAI21_X1  g181(.A(G61), .B1(new_n543), .B2(new_n544), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n608));
  INV_X1    g183(.A(G73), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n518), .ZN(new_n610));
  NAND3_X1  g185(.A1(KEYINPUT83), .A2(G73), .A3(G543), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G48), .B2(new_n519), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n606), .A2(new_n613), .ZN(G305));
  AOI22_X1  g189(.A1(G85), .A2(new_n565), .B1(new_n538), .B2(G47), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT84), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n547), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n617), .A2(new_n510), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(G290));
  NOR2_X1   g194(.A1(new_n538), .A2(KEYINPUT85), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT85), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n536), .B2(new_n537), .ZN(new_n622));
  OAI21_X1  g197(.A(G54), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n530), .A2(G92), .A3(new_n531), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n522), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n510), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(new_n627), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n623), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(G171), .A2(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT87), .Z(G284));
  INV_X1    g210(.A(new_n634), .ZN(G321));
  NAND2_X1  g211(.A1(G286), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n597), .ZN(G297));
  OAI21_X1  g213(.A(new_n637), .B1(G868), .B2(new_n597), .ZN(G280));
  INV_X1    g214(.A(new_n631), .ZN(new_n640));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(G860), .ZN(G148));
  NOR2_X1   g217(.A1(new_n577), .A2(G868), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n631), .A2(G559), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(G868), .B2(new_n644), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g221(.A1(new_n466), .A2(new_n468), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n647), .A2(G2105), .A3(new_n479), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT12), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  MUX2_X1   g226(.A(G99), .B(G111), .S(G2105), .Z(new_n652));
  AOI22_X1  g227(.A1(new_n487), .A2(G123), .B1(G2104), .B2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G135), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n653), .B1(new_n654), .B2(new_n492), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT88), .B(G2096), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n651), .A2(new_n657), .ZN(G156));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT15), .B(G2435), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2427), .ZN(new_n662));
  INV_X1    g237(.A(G2430), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n659), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1341), .B(G1348), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n665), .A2(new_n671), .ZN(new_n673));
  AND3_X1   g248(.A1(new_n672), .A2(G14), .A3(new_n673), .ZN(G401));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT18), .ZN(new_n681));
  INV_X1    g256(.A(new_n677), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(KEYINPUT17), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n678), .B1(new_n684), .B2(new_n675), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(new_n676), .B2(new_n683), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n676), .A2(new_n679), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n682), .B1(new_n687), .B2(KEYINPUT17), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n681), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G2096), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G2100), .ZN(G227));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1961), .B(G1966), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT20), .Z(new_n700));
  NOR2_X1   g275(.A1(new_n693), .A2(new_n695), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n702), .A2(new_n698), .A3(new_n696), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n703), .C1(new_n698), .C2(new_n702), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1991), .B(G1996), .Z(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n706), .B(new_n709), .ZN(G229));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n711));
  INV_X1    g286(.A(G87), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n563), .A2(new_n564), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n519), .A2(G49), .ZN(new_n714));
  AOI21_X1  g289(.A(G74), .B1(new_n542), .B2(new_n545), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n510), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n711), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n603), .A2(KEYINPUT91), .A3(new_n604), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G23), .B(new_n719), .S(G16), .Z(new_n720));
  XOR2_X1   g295(.A(KEYINPUT33), .B(G1976), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G6), .B(G305), .S(G16), .Z(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT32), .B(G1981), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G16), .A2(G22), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G166), .B2(G16), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT92), .B(G1971), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR3_X1   g304(.A1(new_n722), .A2(new_n725), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT34), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT93), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n491), .A2(G131), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n487), .A2(G119), .ZN(new_n735));
  AND2_X1   g310(.A1(G107), .A2(G2105), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G95), .B2(new_n470), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n734), .B(new_n735), .C1(new_n461), .C2(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G25), .B(new_n738), .S(G29), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT90), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G16), .A2(G24), .ZN(new_n744));
  INV_X1    g319(.A(G290), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1986), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n743), .B(new_n747), .C1(new_n731), .C2(new_n730), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n733), .A2(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT36), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(KEYINPUT36), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G16), .A2(G19), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n578), .B2(G16), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT95), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1341), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT25), .Z(new_n758));
  INV_X1    g333(.A(G139), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n492), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(G115), .A2(G2104), .ZN(new_n761));
  INV_X1    g336(.A(G127), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n479), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(KEYINPUT96), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n470), .B1(new_n763), .B2(KEYINPUT96), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G29), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n768), .B2(G33), .ZN(new_n770));
  INV_X1    g345(.A(G2072), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT97), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n770), .A2(new_n771), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(KEYINPUT97), .ZN(new_n775));
  NAND2_X1  g350(.A1(G164), .A2(G29), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G27), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2078), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n773), .A2(new_n774), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT31), .B(G11), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT30), .B(G28), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(new_n768), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n655), .B2(new_n768), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT99), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n768), .A2(G26), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT28), .Z(new_n787));
  MUX2_X1   g362(.A(G104), .B(G116), .S(G2105), .Z(new_n788));
  AOI22_X1  g363(.A1(new_n487), .A2(G128), .B1(G2104), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G140), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n492), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n787), .B1(new_n791), .B2(G29), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2067), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n785), .B(new_n793), .C1(new_n778), .C2(new_n777), .ZN(new_n794));
  INV_X1    g369(.A(G16), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G5), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G171), .B2(new_n795), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1961), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n780), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(G21), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G168), .B2(new_n795), .ZN(new_n801));
  INV_X1    g376(.A(G1966), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(KEYINPUT24), .A2(G34), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(KEYINPUT24), .A2(G34), .ZN(new_n806));
  AOI21_X1  g381(.A(G29), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G160), .B2(G29), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(G2084), .ZN(new_n809));
  OR2_X1    g384(.A1(G29), .A2(G32), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n491), .A2(G141), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n487), .A2(G129), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n647), .A2(G2105), .ZN(new_n813));
  NAND3_X1  g388(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT26), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n813), .A2(G105), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n811), .A2(new_n812), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT98), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n810), .B1(new_n820), .B2(new_n768), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT27), .B(G1996), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n821), .A2(new_n822), .B1(G2084), .B2(new_n808), .ZN(new_n824));
  AND4_X1   g399(.A1(new_n803), .A2(new_n809), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(G4), .A2(G16), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT94), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n631), .B2(new_n795), .ZN(new_n828));
  INV_X1    g403(.A(G1348), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n768), .A2(G35), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G162), .B2(new_n768), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT29), .Z(new_n833));
  INV_X1    g408(.A(G2090), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n756), .A2(new_n799), .A3(new_n825), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n795), .A2(G20), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT23), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n597), .B2(new_n795), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT100), .ZN(new_n840));
  INV_X1    g415(.A(G1956), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n842), .B(new_n843), .C1(new_n834), .C2(new_n833), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n836), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n752), .A2(new_n848), .ZN(G150));
  INV_X1    g424(.A(G150), .ZN(G311));
  AOI22_X1  g425(.A1(new_n547), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(new_n510), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n565), .A2(G93), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n538), .A2(G55), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n577), .A2(new_n855), .ZN(new_n858));
  INV_X1    g433(.A(new_n855), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n859), .B(new_n571), .C1(new_n575), .C2(new_n576), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n640), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G860), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n864), .A2(new_n865), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n857), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT102), .Z(G145));
  XNOR2_X1  g446(.A(new_n649), .B(new_n738), .ZN(new_n872));
  MUX2_X1   g447(.A(G106), .B(G118), .S(G2105), .Z(new_n873));
  AOI22_X1  g448(.A1(new_n487), .A2(G130), .B1(G2104), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G142), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n874), .B1(new_n875), .B2(new_n492), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n872), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n767), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n820), .B(KEYINPUT103), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n791), .B(new_n506), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n820), .A2(KEYINPUT103), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n820), .A2(KEYINPUT103), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n882), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(KEYINPUT104), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n819), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n880), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n767), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT104), .B1(new_n881), .B2(new_n884), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n877), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT105), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n892), .B(new_n877), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  OR3_X1    g468(.A1(new_n888), .A2(new_n877), .A3(new_n889), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(G162), .B(G160), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n655), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n890), .A2(new_n897), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n900), .B2(new_n894), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g478(.A1(new_n855), .A2(G868), .ZN(new_n904));
  XNOR2_X1  g479(.A(G290), .B(new_n719), .ZN(new_n905));
  XOR2_X1   g480(.A(G303), .B(G305), .Z(new_n906));
  XOR2_X1   g481(.A(new_n905), .B(new_n906), .Z(new_n907));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n908));
  NAND3_X1  g483(.A1(G299), .A2(new_n908), .A3(new_n640), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT106), .B1(new_n597), .B2(new_n631), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n909), .A2(new_n910), .B1(new_n597), .B2(new_n631), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT41), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n861), .B(new_n644), .Z(new_n917));
  OR2_X1    g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n912), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n907), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n923), .ZN(new_n925));
  INV_X1    g500(.A(new_n907), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n926), .A3(new_n921), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n904), .B1(new_n928), .B2(G868), .ZN(G295));
  AOI21_X1  g504(.A(new_n904), .B1(new_n928), .B2(G868), .ZN(G331));
  NAND2_X1  g505(.A1(G168), .A2(G171), .ZN(new_n931));
  NAND2_X1  g506(.A1(G286), .A2(G301), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n861), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n858), .A2(new_n931), .A3(new_n860), .A4(new_n932), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n913), .A2(new_n915), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n912), .A2(new_n934), .A3(new_n935), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n907), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n907), .B1(new_n937), .B2(new_n938), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n937), .A2(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n926), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n940), .A4(new_n939), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(KEYINPUT107), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT44), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n943), .B(new_n947), .C1(KEYINPUT107), .C2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(G397));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n506), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(KEYINPUT108), .ZN(new_n957));
  AOI21_X1  g532(.A(G1384), .B1(new_n501), .B2(new_n505), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n954), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n484), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n962), .A2(G40), .A3(new_n475), .A4(new_n482), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n791), .B(G2067), .Z(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n967), .A2(KEYINPUT110), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(KEYINPUT110), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n819), .A2(G1996), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n820), .B2(G1996), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n968), .A2(new_n969), .B1(new_n964), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(G290), .A2(G1986), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT109), .ZN(new_n974));
  INV_X1    g549(.A(G1986), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n975), .B2(new_n745), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n964), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n742), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n738), .A2(new_n742), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n964), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n972), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT111), .Z(new_n982));
  INV_X1    g557(.A(G8), .ZN(new_n983));
  INV_X1    g558(.A(G40), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n483), .A2(new_n984), .A3(new_n484), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n985), .B2(new_n958), .ZN(new_n986));
  INV_X1    g561(.A(G86), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n563), .A2(new_n564), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n612), .A2(G651), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n519), .A2(G48), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(G1981), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1981), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n606), .A2(new_n993), .A3(new_n613), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT49), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(KEYINPUT49), .A3(new_n994), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n992), .A2(KEYINPUT116), .A3(KEYINPUT49), .A4(new_n994), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI211_X1 g575(.A(G1976), .B(G288), .C1(new_n1000), .C2(new_n986), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n606), .A2(new_n993), .A3(new_n613), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n986), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n985), .A2(new_n958), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n717), .A2(G1976), .A3(new_n718), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n1005), .A2(G8), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1976), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(G288), .B2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1000), .A2(new_n986), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n986), .A2(new_n1006), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT52), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1004), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n995), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n993), .B1(new_n606), .B2(new_n613), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1002), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT116), .B1(new_n1016), .B2(KEYINPUT49), .ZN(new_n1017));
  INV_X1    g592(.A(new_n999), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n986), .B(new_n1014), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n986), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1020));
  AND4_X1   g595(.A1(new_n1004), .A2(new_n1019), .A3(new_n1012), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT112), .B(G1971), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n985), .B1(new_n956), .B2(new_n954), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n958), .A2(KEYINPUT45), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n963), .B1(new_n958), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n956), .A2(new_n1029), .A3(KEYINPUT50), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT113), .B1(new_n958), .B2(new_n1027), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT114), .B(G2090), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1026), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n1035));
  NOR3_X1   g610(.A1(G166), .A2(new_n1035), .A3(new_n983), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1036), .A2(KEYINPUT115), .A3(new_n1037), .ZN(new_n1041));
  OAI211_X1 g616(.A(G8), .B(new_n1034), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1003), .B1(new_n1022), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1034), .A2(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n1038), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(KEYINPUT119), .B(new_n1045), .C1(new_n1013), .C2(new_n1021), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1042), .A2(KEYINPUT63), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n802), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1051));
  INV_X1    g626(.A(G2084), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1028), .A2(new_n1030), .A3(new_n1052), .A4(new_n1031), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(G8), .A3(G168), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1050), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1048), .A2(new_n1049), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT63), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n985), .B1(new_n958), .B2(new_n1027), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n985), .B(KEYINPUT118), .C1(new_n958), .C2(new_n1027), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n958), .A2(new_n1027), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1032), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1026), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G8), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n1038), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1042), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1058), .B1(new_n1070), .B2(new_n1055), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1043), .B1(new_n1057), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n590), .B2(new_n592), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n594), .A2(new_n595), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1059), .A2(new_n1060), .B1(new_n1027), .B2(new_n958), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1956), .B1(new_n1077), .B2(new_n1062), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n963), .B1(new_n958), .B2(KEYINPUT45), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n956), .A2(new_n954), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1076), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1064), .A2(new_n841), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1082), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1076), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1087), .A3(KEYINPUT61), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1005), .A2(G2067), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n829), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(new_n631), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1089), .B(new_n640), .C1(new_n1090), .C2(new_n829), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT60), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(new_n640), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1088), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT61), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n1005), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1996), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1079), .A2(new_n1080), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1005), .A2(KEYINPUT121), .A3(new_n1101), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT122), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1104), .A2(new_n1106), .A3(new_n1110), .A4(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1100), .B1(new_n1112), .B2(new_n578), .ZN(new_n1113));
  AOI211_X1 g688(.A(KEYINPUT59), .B(new_n577), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1086), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1087), .B1(new_n1116), .B2(new_n1092), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT120), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1119), .B(new_n1087), .C1(new_n1116), .C2(new_n1092), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1099), .A2(new_n1115), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(G2078), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n961), .A2(new_n1079), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1961), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1090), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1079), .A2(new_n1080), .A3(new_n778), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1122), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G171), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1079), .A2(new_n1080), .A3(KEYINPUT53), .A4(new_n778), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1126), .A2(new_n1128), .A3(G301), .A4(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1130), .A2(KEYINPUT54), .A3(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1070), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1126), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1129), .A2(G171), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1135), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(G286), .A2(G8), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1051), .A2(new_n1053), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1145), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT51), .ZN(new_n1150));
  OAI21_X1  g725(.A(G8), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1144), .B(KEYINPUT124), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g728(.A(KEYINPUT51), .B(new_n1145), .C1(new_n1054), .C2(G8), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1149), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1134), .A2(new_n1143), .A3(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1072), .B(KEYINPUT126), .C1(new_n1121), .C2(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1155), .A2(KEYINPUT62), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(KEYINPUT62), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1070), .B1(new_n1140), .B2(new_n1139), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1166), .A2(new_n1088), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1163), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1169), .A2(new_n1155), .A3(new_n1143), .A4(new_n1134), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT126), .B1(new_n1170), .B2(new_n1072), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n982), .B1(new_n1162), .B2(new_n1171), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n965), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT46), .B1(new_n965), .B2(G1996), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n966), .A2(new_n886), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1173), .A2(new_n1174), .B1(new_n964), .B2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT47), .Z(new_n1177));
  NOR2_X1   g752(.A1(new_n974), .A2(new_n965), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT48), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n972), .A2(new_n980), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n791), .A2(G2067), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n972), .B2(new_n978), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n1183), .A2(KEYINPUT127), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n965), .B1(new_n1183), .B2(KEYINPUT127), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1181), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1172), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g762(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1189));
  NAND3_X1  g763(.A1(new_n902), .A2(new_n948), .A3(new_n1189), .ZN(G225));
  INV_X1    g764(.A(G225), .ZN(G308));
endmodule


