//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT67), .Z(new_n463));
  OAI21_X1  g038(.A(G2105), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(KEYINPUT68), .A3(G101), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(G101), .A3(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n468), .A2(G137), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n464), .A2(new_n475), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n467), .A2(new_n469), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n479), .B(new_n482), .C1(G136), .C2(new_n468), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n469), .B2(G114), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n492), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT71), .B1(new_n494), .B2(new_n489), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n465), .B2(new_n466), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n497), .B(new_n500), .C1(new_n466), .C2(new_n465), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n493), .A2(new_n495), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(KEYINPUT73), .B2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT73), .B1(new_n508), .B2(KEYINPUT5), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n511), .B(G543), .C1(new_n512), .C2(KEYINPUT72), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n510), .A2(G62), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT74), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n505), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n510), .A2(G88), .A3(new_n513), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(G166));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n510), .A2(new_n513), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT75), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n521), .A2(G51), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n510), .A2(G89), .A3(new_n513), .A4(new_n518), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n527), .A2(new_n533), .ZN(G168));
  NAND3_X1  g109(.A1(new_n510), .A2(G64), .A3(new_n513), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n505), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n510), .A2(new_n513), .A3(new_n518), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n539), .A2(G90), .B1(G52), .B2(new_n521), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  NAND4_X1  g117(.A1(new_n510), .A2(G81), .A3(new_n513), .A4(new_n518), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(new_n520), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n510), .A2(G56), .A3(new_n513), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n505), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  OAI211_X1 g129(.A(G65), .B(new_n513), .C1(new_n507), .C2(new_n509), .ZN(new_n555));
  AND2_X1   g130(.A1(G78), .A2(G543), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n555), .A2(new_n557), .A3(KEYINPUT78), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(G651), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n560), .A2(KEYINPUT79), .A3(G651), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(KEYINPUT76), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n521), .A2(G53), .A3(new_n568), .ZN(new_n569));
  XOR2_X1   g144(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n520), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n539), .ZN(new_n574));
  INV_X1    g149(.A(G91), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n566), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G168), .ZN(G286));
  NAND2_X1  g154(.A1(new_n514), .A2(new_n516), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(new_n523), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT80), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n584), .B1(new_n517), .B2(new_n523), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(G303));
  AOI22_X1  g161(.A1(new_n539), .A2(G87), .B1(G49), .B2(new_n521), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n510), .A2(new_n513), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n589), .B2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT81), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(G288));
  OAI211_X1 g171(.A(G61), .B(new_n513), .C1(new_n507), .C2(new_n509), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n505), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n510), .A2(G86), .A3(new_n513), .A4(new_n518), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n602));
  INV_X1    g177(.A(G48), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n520), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n518), .A2(KEYINPUT82), .A3(G48), .A4(G543), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n600), .A2(new_n601), .A3(new_n606), .ZN(G305));
  AOI22_X1  g182(.A1(new_n589), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(new_n505), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n539), .A2(G85), .B1(G47), .B2(new_n521), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  AND3_X1   g187(.A1(new_n539), .A2(KEYINPUT10), .A3(G92), .ZN(new_n613));
  AOI21_X1  g188(.A(KEYINPUT10), .B1(new_n539), .B2(G92), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n588), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G651), .ZN(new_n619));
  INV_X1    g194(.A(G54), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n520), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n612), .B1(new_n622), .B2(G868), .ZN(G284));
  XOR2_X1   g198(.A(G284), .B(KEYINPUT83), .Z(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n576), .B1(new_n564), .B2(new_n565), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(G868), .B2(new_n626), .ZN(G297));
  OAI21_X1  g202(.A(new_n625), .B1(G868), .B2(new_n626), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n622), .B1(new_n629), .B2(G860), .ZN(G148));
  INV_X1    g205(.A(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n545), .B2(new_n548), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n619), .B1(new_n620), .B2(new_n520), .C1(new_n613), .C2(new_n614), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n633), .A2(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n632), .B1(new_n634), .B2(new_n631), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n460), .A2(new_n470), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(KEYINPUT12), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(KEYINPUT12), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n468), .A2(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n480), .A2(G123), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n469), .A2(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n641), .A2(new_n642), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n643), .A2(new_n649), .A3(new_n650), .ZN(G156));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(new_n665), .A3(G14), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT84), .ZN(G401));
  XNOR2_X1  g242(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT85), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n668), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2100), .ZN(new_n676));
  INV_X1    g251(.A(new_n672), .ZN(new_n677));
  NOR2_X1   g252(.A1(G2072), .A2(G2078), .ZN(new_n678));
  OAI22_X1  g253(.A1(new_n677), .A2(new_n668), .B1(new_n442), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2096), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n676), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n685), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(new_n689), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n702), .A2(new_n705), .A3(new_n703), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(G229));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n468), .A2(G131), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n480), .A2(G119), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n469), .A2(G107), .ZN(new_n715));
  OAI21_X1  g290(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n713), .B(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT88), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n712), .B1(new_n719), .B2(new_n711), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  XOR2_X1   g296(.A(new_n720), .B(new_n721), .Z(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(KEYINPUT89), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G24), .ZN(new_n725));
  INV_X1    g300(.A(G290), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1986), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n724), .A2(G23), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n592), .B2(new_n724), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT33), .B(G1976), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n724), .A2(G22), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G166), .B2(new_n724), .ZN(new_n735));
  INV_X1    g310(.A(G1971), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G6), .A2(G16), .ZN(new_n738));
  INV_X1    g313(.A(G305), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G16), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT32), .B(G1981), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n733), .A2(new_n737), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(KEYINPUT34), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(KEYINPUT34), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n722), .A2(KEYINPUT89), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n729), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT90), .B(KEYINPUT36), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G29), .A2(G35), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G162), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2090), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G164), .A2(new_n711), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G27), .B2(new_n711), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n724), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n724), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(G1966), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n756), .A2(new_n757), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n760), .A2(G1966), .ZN(new_n763));
  NOR4_X1   g338(.A1(new_n758), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G34), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n765), .A2(KEYINPUT24), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(KEYINPUT24), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n711), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G160), .B2(new_n711), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT92), .Z(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT93), .ZN(new_n773));
  NOR2_X1   g348(.A1(G5), .A2(G16), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT95), .Z(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G301), .B2(new_n724), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT96), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G1961), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n754), .A2(new_n764), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n770), .A2(new_n771), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n468), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n480), .A2(G129), .ZN(new_n782));
  NAND3_X1  g357(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT26), .Z(new_n784));
  NAND3_X1  g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(new_n711), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n711), .B2(G32), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT27), .B(G1996), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n780), .B1(new_n788), .B2(new_n789), .C1(new_n777), .C2(G1961), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT97), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n468), .A2(G140), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n480), .A2(G128), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n469), .A2(G116), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G29), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n711), .A2(G26), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT28), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2067), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n788), .A2(new_n789), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT31), .B(G11), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT94), .B(G28), .Z(new_n804));
  AOI21_X1  g379(.A(G29), .B1(new_n804), .B2(KEYINPUT30), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(KEYINPUT30), .B2(new_n804), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n803), .B(new_n806), .C1(new_n648), .C2(new_n711), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n711), .A2(G33), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(new_n469), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n811));
  NAND2_X1  g386(.A1(G103), .A2(G2104), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G2105), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n469), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n468), .A2(G139), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n808), .B1(new_n817), .B2(new_n711), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n807), .B1(new_n818), .B2(G2072), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n802), .B(new_n819), .C1(G2072), .C2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n622), .A2(G16), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G4), .B2(G16), .ZN(new_n822));
  INV_X1    g397(.A(G1348), .ZN(new_n823));
  AOI211_X1 g398(.A(new_n801), .B(new_n820), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(G16), .A2(G19), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n549), .B2(G16), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT91), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(G1341), .Z(new_n828));
  OAI211_X1 g403(.A(new_n824), .B(new_n828), .C1(new_n823), .C2(new_n822), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n724), .A2(G20), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT23), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n626), .B2(new_n724), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT100), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT99), .B(G1956), .Z(new_n834));
  AND2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR4_X1   g410(.A1(new_n779), .A2(new_n791), .A3(new_n829), .A4(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n833), .A2(new_n834), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n749), .A2(new_n836), .A3(new_n837), .ZN(G150));
  INV_X1    g413(.A(G150), .ZN(G311));
  AOI22_X1  g414(.A1(new_n539), .A2(G93), .B1(G55), .B2(new_n521), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n510), .A2(G67), .A3(new_n513), .ZN(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G651), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n622), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  INV_X1    g424(.A(new_n545), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n546), .A2(new_n547), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G651), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n850), .A2(new_n840), .A3(new_n852), .A4(new_n844), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n510), .A2(G93), .A3(new_n513), .A4(new_n518), .ZN(new_n854));
  INV_X1    g429(.A(G55), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n520), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n505), .B1(new_n841), .B2(new_n842), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n548), .A2(new_n545), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n849), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT101), .ZN(new_n863));
  INV_X1    g438(.A(G860), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n847), .B1(new_n863), .B2(new_n865), .ZN(G145));
  INV_X1    g441(.A(new_n501), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n500), .B1(new_n460), .B2(new_n497), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT102), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n499), .A2(new_n870), .A3(new_n501), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n490), .A2(new_n492), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(new_n796), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n796), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n719), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n718), .A3(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n468), .A2(G142), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n480), .A2(G130), .ZN(new_n883));
  OR2_X1    g458(.A1(G106), .A2(G2105), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n884), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n640), .A2(new_n882), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(new_n639), .A3(new_n638), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n817), .A2(new_n786), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n816), .A2(new_n785), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n889), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n881), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(G160), .B(new_n648), .ZN(new_n896));
  XNOR2_X1  g471(.A(G162), .B(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n881), .B1(new_n892), .B2(new_n893), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n879), .A3(new_n880), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n897), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT103), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n904));
  AOI211_X1 g479(.A(new_n904), .B(new_n897), .C1(new_n899), .C2(new_n900), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n898), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n859), .B(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n634), .ZN(new_n910));
  NAND2_X1  g485(.A1(G299), .A2(new_n633), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n622), .A2(new_n626), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n910), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n915), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n917), .B1(new_n918), .B2(new_n910), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT42), .ZN(new_n920));
  XNOR2_X1  g495(.A(G290), .B(new_n739), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n591), .B(G166), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n920), .A2(new_n923), .ZN(new_n925));
  OAI21_X1  g500(.A(G868), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n845), .A2(new_n631), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(G295));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n927), .ZN(G331));
  NAND2_X1  g504(.A1(new_n916), .A2(new_n914), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n510), .A2(G90), .A3(new_n513), .A4(new_n518), .ZN(new_n931));
  INV_X1    g506(.A(G52), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n931), .B1(new_n932), .B2(new_n520), .ZN(new_n933));
  OAI22_X1  g508(.A1(new_n527), .A2(new_n533), .B1(new_n537), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT75), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n526), .B(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n531), .A2(new_n532), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n936), .A2(new_n538), .A3(new_n937), .A4(new_n540), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  OR3_X1    g514(.A1(new_n939), .A2(new_n859), .A3(KEYINPUT107), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n934), .A2(new_n938), .A3(new_n853), .A4(new_n858), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT107), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n939), .A2(new_n859), .A3(KEYINPUT106), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT106), .B1(new_n939), .B2(new_n859), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n940), .B(new_n942), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n859), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(KEYINPUT108), .A3(new_n941), .ZN(new_n947));
  OR3_X1    g522(.A1(new_n939), .A2(new_n859), .A3(KEYINPUT108), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n930), .A2(new_n945), .B1(new_n949), .B2(new_n918), .ZN(new_n950));
  AOI21_X1  g525(.A(G37), .B1(new_n950), .B2(new_n923), .ZN(new_n951));
  XNOR2_X1  g526(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n918), .A2(KEYINPUT109), .A3(new_n913), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n914), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n916), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n949), .ZN(new_n957));
  INV_X1    g532(.A(new_n945), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n956), .A2(new_n957), .B1(new_n958), .B2(new_n918), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n951), .B(new_n952), .C1(new_n959), .C2(new_n923), .ZN(new_n960));
  INV_X1    g535(.A(new_n952), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n930), .A2(new_n945), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n949), .A2(new_n918), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n923), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G37), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n950), .A2(new_n923), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n961), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n960), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n966), .A2(new_n967), .A3(new_n961), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n951), .B1(new_n959), .B2(new_n923), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n970), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n972));
  MUX2_X1   g547(.A(new_n969), .B(new_n972), .S(KEYINPUT44), .Z(G397));
  INV_X1    g548(.A(G1966), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n464), .A2(new_n475), .A3(G40), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n872), .B2(new_n874), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n975), .B(new_n976), .C1(new_n977), .C2(KEYINPUT45), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n873), .B1(new_n869), .B2(new_n871), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(G1384), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n975), .B1(new_n984), .B2(new_n976), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n974), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT118), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n977), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n503), .A2(new_n979), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n976), .A3(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n992), .A2(G2084), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n994), .B(new_n974), .C1(new_n981), .C2(new_n985), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n987), .A2(G168), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n996), .A2(G8), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n996), .B2(G8), .ZN(new_n1000));
  NAND2_X1  g575(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n987), .A2(new_n993), .A3(new_n995), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(G8), .A3(G286), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT62), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1000), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n996), .A2(G8), .A3(new_n998), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n1001), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT62), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n1005), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n583), .A2(G8), .A3(new_n585), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n583), .A2(new_n585), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n990), .A2(new_n982), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n976), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n736), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n875), .A2(new_n979), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT50), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT112), .B(G2090), .Z(new_n1025));
  NAND3_X1  g600(.A1(new_n503), .A2(new_n988), .A3(new_n979), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1024), .A2(new_n976), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1018), .B1(new_n1028), .B2(KEYINPUT116), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1022), .A2(new_n1030), .A3(new_n1027), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1017), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n1033));
  OAI21_X1  g608(.A(G1981), .B1(new_n599), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G305), .B(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT115), .B1(new_n1035), .B2(KEYINPUT49), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1034), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(G305), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n464), .A2(new_n475), .A3(G40), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n983), .A2(new_n1044), .A3(G1384), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1045), .B2(new_n1018), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n875), .A2(new_n976), .A3(new_n979), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(KEYINPUT113), .A3(G8), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1046), .A2(new_n1048), .B1(new_n1035), .B2(KEYINPUT49), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1042), .A2(new_n1049), .ZN(new_n1050));
  AND4_X1   g625(.A1(new_n976), .A2(new_n989), .A3(new_n991), .A4(new_n1025), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1044), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1971), .B1(new_n1052), .B2(new_n1020), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1017), .B(G8), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n592), .A2(G1976), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1045), .A2(new_n1043), .A3(new_n1018), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT113), .B1(new_n1047), .B2(G8), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT52), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1060));
  INV_X1    g635(.A(G1976), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n593), .A2(new_n1061), .A3(new_n595), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .A4(new_n1055), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1050), .A2(new_n1054), .A3(new_n1059), .A4(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1032), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1052), .A2(new_n757), .A3(new_n1020), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  INV_X1    g643(.A(G1961), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1067), .A2(new_n1068), .B1(new_n992), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n984), .A2(new_n976), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT117), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1068), .A2(G2078), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1072), .A2(new_n978), .A3(new_n980), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G301), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1066), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1007), .A2(new_n1012), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT63), .ZN(new_n1079));
  OAI21_X1  g654(.A(G8), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1017), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1042), .A2(new_n1049), .B1(new_n1058), .B2(KEYINPUT52), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n1054), .A4(new_n1064), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G286), .A2(new_n1018), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n995), .A2(new_n993), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1072), .A2(new_n978), .A3(new_n980), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n994), .B1(new_n1087), .B2(new_n974), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT119), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n1085), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1084), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1092), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1004), .B2(new_n1085), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1066), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(new_n1096), .B2(new_n1079), .ZN(new_n1097));
  NOR2_X1   g672(.A1(G305), .A2(G1981), .ZN(new_n1098));
  NOR2_X1   g673(.A1(G288), .A2(G1976), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1050), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1048), .B2(new_n1046), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1083), .A2(new_n1064), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(new_n1054), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1078), .B1(new_n1097), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT63), .B1(new_n1107), .B2(new_n1066), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT120), .B(new_n1104), .C1(new_n1108), .C2(new_n1093), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1019), .A2(new_n984), .A3(new_n976), .A4(new_n1073), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1070), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(G171), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1070), .A2(G301), .A3(new_n1074), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(KEYINPUT54), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1111), .A2(G171), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1075), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1066), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1956), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n977), .A2(new_n988), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1026), .A2(new_n976), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT56), .B(G2072), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT57), .B1(new_n573), .B2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1126), .B(new_n576), .C1(new_n564), .C2(new_n565), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1126), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n626), .A2(new_n1128), .ZN(new_n1129));
  OAI221_X1 g704(.A(new_n1122), .B1(new_n1021), .B2(new_n1124), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1122), .B1(new_n1021), .B2(new_n1124), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1130), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT58), .B(G1341), .ZN(new_n1138));
  OAI22_X1  g713(.A1(new_n1021), .A2(G1996), .B1(new_n1045), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n549), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT59), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n992), .A2(new_n823), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1047), .A2(G2067), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1145), .A2(KEYINPUT123), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT123), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n622), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT123), .B(new_n633), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1137), .B(new_n1141), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1130), .A2(new_n622), .A3(new_n1145), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1154), .A2(new_n1133), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1118), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1010), .A2(new_n1005), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1077), .A2(new_n1106), .A3(new_n1109), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1023), .A2(new_n982), .A3(new_n976), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT110), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1161), .A2(G1996), .A3(new_n785), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT111), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n796), .B(G2067), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1160), .A2(G1996), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1161), .A2(new_n1164), .B1(new_n786), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n718), .B(new_n721), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1161), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1163), .B(new_n1166), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  OR2_X1    g744(.A1(G290), .A2(G1986), .ZN(new_n1170));
  NAND2_X1  g745(.A1(G290), .A2(G1986), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1160), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1159), .A2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1165), .B(KEYINPUT46), .Z(new_n1175));
  OAI21_X1  g750(.A(new_n1161), .B1(new_n785), .B2(new_n1164), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1178));
  XNOR2_X1  g753(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1170), .A2(new_n1160), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT48), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1179), .B1(new_n1169), .B2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1163), .A2(new_n721), .A3(new_n719), .A4(new_n1166), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n796), .A2(G2067), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1168), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1174), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g762(.A1(new_n681), .A2(G319), .A3(new_n666), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n1189), .B1(new_n707), .B2(new_n708), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n1190), .A2(new_n906), .ZN(new_n1191));
  INV_X1    g765(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n969), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1193), .A2(KEYINPUT126), .ZN(new_n1194));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n969), .A2(new_n1195), .A3(new_n1192), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n1194), .A2(KEYINPUT127), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n1198));
  AOI211_X1 g772(.A(KEYINPUT126), .B(new_n1191), .C1(new_n968), .C2(new_n960), .ZN(new_n1199));
  AOI21_X1  g773(.A(new_n1195), .B1(new_n969), .B2(new_n1192), .ZN(new_n1200));
  OAI21_X1  g774(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1197), .A2(new_n1201), .ZN(G308));
  NAND2_X1  g776(.A1(new_n1194), .A2(new_n1196), .ZN(G225));
endmodule


