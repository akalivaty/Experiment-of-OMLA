

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766;

  OR2_X1 U377 ( .A1(n690), .A2(G902), .ZN(n427) );
  AND2_X1 U378 ( .A1(n425), .A2(n632), .ZN(n355) );
  XOR2_X1 U379 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n356) );
  XNOR2_X2 U380 ( .A(n422), .B(KEYINPUT0), .ZN(n644) );
  XNOR2_X2 U381 ( .A(n427), .B(G472), .ZN(n565) );
  NOR2_X1 U382 ( .A1(n581), .A2(n582), .ZN(n618) );
  INV_X1 U383 ( .A(n686), .ZN(n687) );
  XNOR2_X1 U384 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n487) );
  AND2_X1 U385 ( .A1(n381), .A2(n611), .ZN(n753) );
  NAND2_X1 U386 ( .A1(n398), .A2(n396), .ZN(n673) );
  AND2_X1 U387 ( .A1(n401), .A2(n399), .ZN(n398) );
  OR2_X1 U388 ( .A1(n765), .A2(n766), .ZN(n430) );
  NOR2_X1 U389 ( .A1(n553), .A2(n446), .ZN(n445) );
  XNOR2_X1 U390 ( .A(n565), .B(KEYINPUT6), .ZN(n634) );
  XNOR2_X1 U391 ( .A(n616), .B(KEYINPUT91), .ZN(n617) );
  XNOR2_X1 U392 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U393 ( .A(n443), .B(n365), .ZN(n734) );
  XNOR2_X1 U394 ( .A(n428), .B(G146), .ZN(n443) );
  XNOR2_X1 U395 ( .A(n522), .B(n521), .ZN(n428) );
  XNOR2_X1 U396 ( .A(n487), .B(n489), .ZN(n410) );
  XNOR2_X1 U397 ( .A(n534), .B(n484), .ZN(n380) );
  XNOR2_X1 U398 ( .A(n460), .B(G146), .ZN(n486) );
  XNOR2_X1 U399 ( .A(KEYINPUT4), .B(G137), .ZN(n519) );
  AND2_X1 U400 ( .A1(n599), .A2(n431), .ZN(n357) );
  XNOR2_X1 U401 ( .A(n600), .B(KEYINPUT39), .ZN(n609) );
  XNOR2_X1 U402 ( .A(n658), .B(KEYINPUT45), .ZN(n358) );
  BUF_X1 U403 ( .A(n730), .Z(n359) );
  NAND2_X1 U404 ( .A1(n526), .A2(n380), .ZN(n362) );
  NAND2_X1 U405 ( .A1(n360), .A2(n361), .ZN(n363) );
  NAND2_X1 U406 ( .A1(n362), .A2(n363), .ZN(n702) );
  INV_X1 U407 ( .A(n526), .ZN(n360) );
  INV_X1 U408 ( .A(n380), .ZN(n361) );
  XNOR2_X1 U409 ( .A(n658), .B(KEYINPUT45), .ZN(n678) );
  XNOR2_X1 U410 ( .A(n570), .B(n569), .ZN(n578) );
  NAND2_X1 U411 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U412 ( .A(n430), .B(n429), .ZN(n383) );
  XNOR2_X1 U413 ( .A(n417), .B(n372), .ZN(n446) );
  OR2_X1 U414 ( .A1(n734), .A2(G902), .ZN(n535) );
  XNOR2_X1 U415 ( .A(n511), .B(KEYINPUT25), .ZN(n512) );
  XNOR2_X1 U416 ( .A(n423), .B(n473), .ZN(n522) );
  INV_X1 U417 ( .A(G134), .ZN(n473) );
  XNOR2_X1 U418 ( .A(n441), .B(n440), .ZN(n738) );
  XNOR2_X1 U419 ( .A(n464), .B(n370), .ZN(n440) );
  XNOR2_X1 U420 ( .A(n470), .B(n751), .ZN(n441) );
  XNOR2_X1 U421 ( .A(n379), .B(n395), .ZN(n378) );
  XNOR2_X1 U422 ( .A(n488), .B(n486), .ZN(n395) );
  XNOR2_X1 U423 ( .A(n410), .B(n423), .ZN(n379) );
  XOR2_X1 U424 ( .A(G104), .B(G122), .Z(n467) );
  INV_X1 U425 ( .A(KEYINPUT67), .ZN(n465) );
  AND2_X1 U426 ( .A1(n444), .A2(KEYINPUT34), .ZN(n424) );
  OR2_X1 U427 ( .A1(n446), .A2(n630), .ZN(n426) );
  XNOR2_X1 U428 ( .A(n382), .B(n416), .ZN(n381) );
  XNOR2_X1 U429 ( .A(G116), .B(G113), .ZN(n421) );
  XNOR2_X1 U430 ( .A(G119), .B(G137), .ZN(n505) );
  XNOR2_X1 U431 ( .A(n461), .B(KEYINPUT10), .ZN(n751) );
  XOR2_X1 U432 ( .A(KEYINPUT8), .B(n474), .Z(n504) );
  NAND2_X1 U433 ( .A1(G234), .A2(n754), .ZN(n474) );
  AND2_X1 U434 ( .A1(n719), .A2(n438), .ZN(n606) );
  INV_X1 U435 ( .A(n577), .ZN(n439) );
  INV_X1 U436 ( .A(n642), .ZN(n431) );
  OR2_X1 U437 ( .A1(n613), .A2(n388), .ZN(n387) );
  INV_X1 U438 ( .A(n615), .ZN(n390) );
  NOR2_X1 U439 ( .A1(n403), .A2(n624), .ZN(n402) );
  NOR2_X1 U440 ( .A1(n400), .A2(n367), .ZN(n399) );
  NOR2_X1 U441 ( .A1(n625), .A2(KEYINPUT105), .ZN(n400) );
  XNOR2_X1 U442 ( .A(n483), .B(n434), .ZN(n543) );
  XNOR2_X1 U443 ( .A(n435), .B(G478), .ZN(n434) );
  INV_X1 U444 ( .A(KEYINPUT103), .ZN(n435) );
  XNOR2_X1 U445 ( .A(n472), .B(n471), .ZN(n581) );
  NAND2_X1 U446 ( .A1(n374), .A2(G210), .ZN(n454) );
  INV_X1 U447 ( .A(KEYINPUT46), .ZN(n429) );
  INV_X1 U448 ( .A(KEYINPUT48), .ZN(n416) );
  XNOR2_X1 U449 ( .A(G902), .B(KEYINPUT15), .ZN(n684) );
  XNOR2_X1 U450 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U451 ( .A(G113), .B(G143), .ZN(n466) );
  XOR2_X1 U452 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n463) );
  INV_X1 U453 ( .A(G125), .ZN(n460) );
  XNOR2_X1 U454 ( .A(n561), .B(KEYINPUT90), .ZN(n613) );
  NAND2_X1 U455 ( .A1(G953), .A2(n389), .ZN(n388) );
  INV_X1 U456 ( .A(G900), .ZN(n389) );
  INV_X1 U457 ( .A(n543), .ZN(n582) );
  AND2_X1 U458 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U459 ( .A(n443), .B(n527), .ZN(n690) );
  INV_X1 U460 ( .A(KEYINPUT102), .ZN(n476) );
  NAND2_X1 U461 ( .A1(n426), .A2(n368), .ZN(n392) );
  NAND2_X1 U462 ( .A1(n355), .A2(n424), .ZN(n393) );
  XNOR2_X1 U463 ( .A(n566), .B(n386), .ZN(n385) );
  INV_X1 U464 ( .A(KEYINPUT28), .ZN(n386) );
  INV_X1 U465 ( .A(n630), .ZN(n444) );
  XNOR2_X1 U466 ( .A(KEYINPUT16), .B(G122), .ZN(n484) );
  XNOR2_X1 U467 ( .A(n507), .B(n456), .ZN(n508) );
  XNOR2_X1 U468 ( .A(n738), .B(n457), .ZN(n739) );
  XNOR2_X1 U469 ( .A(KEYINPUT92), .B(G140), .ZN(n532) );
  NOR2_X1 U470 ( .A1(n686), .A2(n664), .ZN(n665) );
  AND2_X1 U471 ( .A1(n608), .A2(n449), .ZN(n725) );
  INV_X1 U472 ( .A(KEYINPUT40), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n437), .B(n436), .ZN(n580) );
  INV_X1 U474 ( .A(KEYINPUT36), .ZN(n436) );
  NAND2_X1 U475 ( .A1(n606), .A2(n579), .ZN(n437) );
  NOR2_X1 U476 ( .A1(n597), .A2(n449), .ZN(n584) );
  BUF_X1 U477 ( .A(G110), .Z(n411) );
  NAND2_X1 U478 ( .A1(n397), .A2(n624), .ZN(n396) );
  XNOR2_X1 U479 ( .A(n744), .B(n412), .ZN(n746) );
  XNOR2_X1 U480 ( .A(n745), .B(n743), .ZN(n412) );
  INV_X1 U481 ( .A(KEYINPUT56), .ZN(n450) );
  INV_X1 U482 ( .A(n750), .ZN(n452) );
  INV_X2 U483 ( .A(G953), .ZN(n754) );
  XOR2_X1 U484 ( .A(n494), .B(n493), .Z(n364) );
  XOR2_X1 U485 ( .A(n534), .B(n533), .Z(n365) );
  AND2_X1 U486 ( .A1(n390), .A2(n387), .ZN(n366) );
  OR2_X1 U487 ( .A1(n636), .A2(n641), .ZN(n367) );
  AND2_X1 U488 ( .A1(n632), .A2(n631), .ZN(n368) );
  OR2_X1 U489 ( .A1(n592), .A2(n591), .ZN(n369) );
  AND2_X1 U490 ( .A1(G214), .A2(n523), .ZN(n370) );
  AND2_X1 U491 ( .A1(n634), .A2(n625), .ZN(n371) );
  XOR2_X1 U492 ( .A(KEYINPUT106), .B(KEYINPUT33), .Z(n372) );
  XNOR2_X1 U493 ( .A(n702), .B(n378), .ZN(n730) );
  XNOR2_X1 U494 ( .A(n731), .B(n359), .ZN(n373) );
  NOR2_X1 U495 ( .A1(n587), .A2(n603), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n409), .B(n408), .ZN(n765) );
  AND2_X2 U497 ( .A1(n406), .A2(n687), .ZN(n374) );
  AND2_X2 U498 ( .A1(n406), .A2(n687), .ZN(n375) );
  XNOR2_X1 U499 ( .A(n578), .B(n571), .ZN(n405) );
  XNOR2_X1 U500 ( .A(n391), .B(KEYINPUT35), .ZN(n652) );
  NAND2_X1 U501 ( .A1(n393), .A2(n392), .ZN(n391) );
  NOR2_X2 U502 ( .A1(n668), .A2(G953), .ZN(n670) );
  BUF_X1 U503 ( .A(n405), .Z(n376) );
  BUF_X1 U504 ( .A(n578), .Z(n377) );
  NAND2_X2 U505 ( .A1(n407), .A2(n685), .ZN(n406) );
  NAND2_X1 U506 ( .A1(n730), .A2(n684), .ZN(n495) );
  XNOR2_X2 U507 ( .A(n413), .B(n421), .ZN(n526) );
  NOR2_X1 U508 ( .A1(n602), .A2(n369), .ZN(n384) );
  NOR2_X1 U509 ( .A1(n593), .A2(n376), .ZN(n717) );
  NAND2_X1 U510 ( .A1(n385), .A2(n585), .ZN(n593) );
  AND2_X2 U511 ( .A1(n673), .A2(n394), .ZN(n655) );
  XNOR2_X1 U512 ( .A(n394), .B(n676), .ZN(G21) );
  XNOR2_X2 U513 ( .A(n404), .B(n629), .ZN(n394) );
  INV_X1 U514 ( .A(n627), .ZN(n397) );
  NAND2_X1 U515 ( .A1(n627), .A2(n402), .ZN(n401) );
  INV_X1 U516 ( .A(n625), .ZN(n403) );
  NAND2_X1 U517 ( .A1(n627), .A2(n455), .ZN(n404) );
  NOR2_X2 U518 ( .A1(n405), .A2(n617), .ZN(n422) );
  NAND2_X1 U519 ( .A1(n406), .A2(n687), .ZN(n727) );
  NAND2_X1 U520 ( .A1(n447), .A2(n682), .ZN(n407) );
  NAND2_X1 U521 ( .A1(n609), .A2(n601), .ZN(n409) );
  XNOR2_X2 U522 ( .A(n485), .B(n420), .ZN(n413) );
  XNOR2_X1 U523 ( .A(n414), .B(n742), .ZN(G60) );
  NOR2_X2 U524 ( .A1(n741), .A2(n750), .ZN(n414) );
  XNOR2_X1 U525 ( .A(n415), .B(KEYINPUT120), .ZN(G54) );
  NOR2_X2 U526 ( .A1(n737), .A2(n750), .ZN(n415) );
  INV_X1 U527 ( .A(n565), .ZN(n587) );
  NAND2_X1 U528 ( .A1(n418), .A2(n604), .ZN(n417) );
  XNOR2_X2 U529 ( .A(n585), .B(KEYINPUT1), .ZN(n604) );
  NOR2_X1 U530 ( .A1(n634), .A2(n586), .ZN(n418) );
  XNOR2_X2 U531 ( .A(n419), .B(G107), .ZN(n534) );
  XNOR2_X2 U532 ( .A(G104), .B(G110), .ZN(n419) );
  XNOR2_X2 U533 ( .A(G101), .B(KEYINPUT68), .ZN(n420) );
  XNOR2_X2 U534 ( .A(n442), .B(G143), .ZN(n423) );
  INV_X1 U535 ( .A(n446), .ZN(n425) );
  XNOR2_X1 U536 ( .A(n428), .B(n751), .ZN(n757) );
  NAND2_X1 U537 ( .A1(n432), .A2(n431), .ZN(n596) );
  NAND2_X1 U538 ( .A1(n585), .A2(n552), .ZN(n642) );
  XNOR2_X1 U539 ( .A(n433), .B(KEYINPUT30), .ZN(n432) );
  NOR2_X1 U540 ( .A1(n634), .A2(n439), .ZN(n438) );
  XNOR2_X2 U541 ( .A(G128), .B(KEYINPUT73), .ZN(n442) );
  NOR2_X1 U542 ( .A1(n594), .A2(n446), .ZN(n557) );
  NAND2_X1 U543 ( .A1(n627), .A2(n371), .ZN(n635) );
  XNOR2_X1 U544 ( .A(n679), .B(n448), .ZN(n447) );
  INV_X1 U545 ( .A(KEYINPUT78), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n568), .B(KEYINPUT38), .ZN(n598) );
  INV_X1 U547 ( .A(n568), .ZN(n449) );
  XNOR2_X2 U548 ( .A(n495), .B(n364), .ZN(n568) );
  XNOR2_X1 U549 ( .A(n451), .B(n450), .ZN(G51) );
  NAND2_X1 U550 ( .A1(n453), .A2(n452), .ZN(n451) );
  XNOR2_X1 U551 ( .A(n454), .B(n373), .ZN(n453) );
  AND2_X1 U552 ( .A1(n626), .A2(n634), .ZN(n455) );
  XOR2_X1 U553 ( .A(n506), .B(n505), .Z(n456) );
  XNOR2_X1 U554 ( .A(KEYINPUT85), .B(KEYINPUT59), .ZN(n457) );
  INV_X1 U555 ( .A(n724), .ZN(n610) );
  NOR2_X1 U556 ( .A1(n725), .A2(n610), .ZN(n611) );
  XNOR2_X1 U557 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U558 ( .A(n502), .B(n501), .ZN(n503) );
  BUF_X1 U559 ( .A(n565), .Z(n641) );
  XNOR2_X1 U560 ( .A(n509), .B(n508), .ZN(n748) );
  BUF_X1 U561 ( .A(n529), .Z(n636) );
  AND2_X1 U562 ( .A1(n693), .A2(G953), .ZN(n750) );
  INV_X1 U563 ( .A(n671), .ZN(n672) );
  XNOR2_X1 U564 ( .A(n670), .B(n669), .ZN(G75) );
  XOR2_X1 U565 ( .A(KEYINPUT69), .B(KEYINPUT14), .Z(n459) );
  NAND2_X1 U566 ( .A1(G234), .A2(G237), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n459), .B(n458), .ZN(n560) );
  NAND2_X1 U568 ( .A1(G952), .A2(n560), .ZN(n562) );
  XNOR2_X1 U569 ( .A(n486), .B(G140), .ZN(n461) );
  XNOR2_X1 U570 ( .A(KEYINPUT98), .B(KEYINPUT11), .ZN(n462) );
  XNOR2_X1 U571 ( .A(n463), .B(n462), .ZN(n464) );
  NOR2_X1 U572 ( .A1(G953), .A2(G237), .ZN(n523) );
  XNOR2_X1 U573 ( .A(n465), .B(G131), .ZN(n520) );
  XNOR2_X1 U574 ( .A(n520), .B(KEYINPUT99), .ZN(n469) );
  XNOR2_X1 U575 ( .A(n467), .B(n466), .ZN(n468) );
  NOR2_X1 U576 ( .A1(G902), .A2(n738), .ZN(n472) );
  XNOR2_X1 U577 ( .A(KEYINPUT13), .B(G475), .ZN(n471) );
  NAND2_X1 U578 ( .A1(G217), .A2(n504), .ZN(n481) );
  XNOR2_X1 U579 ( .A(G107), .B(KEYINPUT101), .ZN(n475) );
  XNOR2_X1 U580 ( .A(n356), .B(n475), .ZN(n479) );
  XNOR2_X1 U581 ( .A(G116), .B(G122), .ZN(n477) );
  XNOR2_X1 U582 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U583 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U584 ( .A(n522), .B(n482), .Z(n745) );
  NOR2_X1 U585 ( .A1(G902), .A2(n745), .ZN(n483) );
  XNOR2_X2 U586 ( .A(KEYINPUT3), .B(G119), .ZN(n485) );
  XOR2_X1 U587 ( .A(KEYINPUT18), .B(KEYINPUT86), .Z(n488) );
  NAND2_X1 U588 ( .A1(n754), .A2(G224), .ZN(n489) );
  INV_X1 U589 ( .A(G902), .ZN(n491) );
  INV_X1 U590 ( .A(G237), .ZN(n490) );
  NAND2_X1 U591 ( .A1(n491), .A2(n490), .ZN(n496) );
  NAND2_X1 U592 ( .A1(n496), .A2(G210), .ZN(n494) );
  INV_X1 U593 ( .A(KEYINPUT87), .ZN(n492) );
  XNOR2_X1 U594 ( .A(n492), .B(KEYINPUT88), .ZN(n493) );
  AND2_X1 U595 ( .A1(n496), .A2(G214), .ZN(n603) );
  OR2_X1 U596 ( .A1(n598), .A2(n603), .ZN(n497) );
  XOR2_X1 U597 ( .A(KEYINPUT110), .B(n497), .Z(n546) );
  NAND2_X1 U598 ( .A1(n618), .A2(n546), .ZN(n498) );
  XOR2_X1 U599 ( .A(KEYINPUT41), .B(n498), .Z(n594) );
  XOR2_X1 U600 ( .A(KEYINPUT95), .B(KEYINPUT24), .Z(n500) );
  XNOR2_X1 U601 ( .A(KEYINPUT94), .B(KEYINPUT23), .ZN(n499) );
  XNOR2_X1 U602 ( .A(n500), .B(n499), .ZN(n502) );
  XOR2_X1 U603 ( .A(KEYINPUT93), .B(KEYINPUT71), .Z(n501) );
  XNOR2_X1 U604 ( .A(n751), .B(n503), .ZN(n509) );
  NAND2_X1 U605 ( .A1(G221), .A2(n504), .ZN(n507) );
  XOR2_X1 U606 ( .A(n411), .B(G128), .Z(n506) );
  NOR2_X1 U607 ( .A1(G902), .A2(n748), .ZN(n513) );
  NAND2_X1 U608 ( .A1(n684), .A2(G234), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n510), .B(KEYINPUT20), .ZN(n514) );
  NAND2_X1 U610 ( .A1(n514), .A2(G217), .ZN(n511) );
  XNOR2_X1 U611 ( .A(n513), .B(n512), .ZN(n529) );
  NAND2_X1 U612 ( .A1(n514), .A2(G221), .ZN(n516) );
  XOR2_X1 U613 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n515) );
  XNOR2_X1 U614 ( .A(n516), .B(n515), .ZN(n619) );
  NOR2_X1 U615 ( .A1(n636), .A2(n619), .ZN(n517) );
  XNOR2_X1 U616 ( .A(n517), .B(KEYINPUT114), .ZN(n518) );
  XNOR2_X1 U617 ( .A(n518), .B(KEYINPUT49), .ZN(n528) );
  XNOR2_X1 U618 ( .A(n520), .B(n519), .ZN(n521) );
  NAND2_X1 U619 ( .A1(G210), .A2(n523), .ZN(n524) );
  XNOR2_X1 U620 ( .A(n524), .B(KEYINPUT5), .ZN(n525) );
  XNOR2_X1 U621 ( .A(n526), .B(n525), .ZN(n527) );
  INV_X1 U622 ( .A(G472), .ZN(n688) );
  NAND2_X1 U623 ( .A1(n528), .A2(n587), .ZN(n538) );
  NAND2_X1 U624 ( .A1(n529), .A2(n619), .ZN(n586) );
  NAND2_X1 U625 ( .A1(G227), .A2(n754), .ZN(n530) );
  XNOR2_X1 U626 ( .A(G101), .B(n530), .ZN(n531) );
  XNOR2_X1 U627 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X2 U628 ( .A(n535), .B(G469), .ZN(n585) );
  INV_X1 U629 ( .A(n604), .ZN(n625) );
  NAND2_X1 U630 ( .A1(n586), .A2(n625), .ZN(n536) );
  XOR2_X1 U631 ( .A(KEYINPUT50), .B(n536), .Z(n537) );
  NOR2_X1 U632 ( .A1(n538), .A2(n537), .ZN(n540) );
  NOR2_X1 U633 ( .A1(n586), .A2(n587), .ZN(n539) );
  AND2_X1 U634 ( .A1(n539), .A2(n604), .ZN(n638) );
  OR2_X1 U635 ( .A1(n540), .A2(n638), .ZN(n541) );
  XNOR2_X1 U636 ( .A(KEYINPUT51), .B(n541), .ZN(n542) );
  NOR2_X1 U637 ( .A1(n594), .A2(n542), .ZN(n554) );
  AND2_X1 U638 ( .A1(n581), .A2(n543), .ZN(n601) );
  INV_X1 U639 ( .A(n601), .ZN(n545) );
  NOR2_X1 U640 ( .A1(n543), .A2(n581), .ZN(n721) );
  INV_X1 U641 ( .A(n721), .ZN(n544) );
  NAND2_X1 U642 ( .A1(n545), .A2(n544), .ZN(n645) );
  NAND2_X1 U643 ( .A1(n546), .A2(n645), .ZN(n547) );
  XNOR2_X1 U644 ( .A(KEYINPUT115), .B(n547), .ZN(n551) );
  INV_X1 U645 ( .A(n618), .ZN(n549) );
  AND2_X1 U646 ( .A1(n598), .A2(n603), .ZN(n548) );
  NOR2_X1 U647 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U648 ( .A1(n551), .A2(n550), .ZN(n553) );
  INV_X1 U649 ( .A(n586), .ZN(n552) );
  NOR2_X1 U650 ( .A1(n554), .A2(n445), .ZN(n555) );
  XNOR2_X1 U651 ( .A(n555), .B(KEYINPUT52), .ZN(n556) );
  NOR2_X1 U652 ( .A1(n562), .A2(n556), .ZN(n558) );
  NOR2_X1 U653 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U654 ( .A(KEYINPUT116), .B(n559), .Z(n666) );
  NAND2_X1 U655 ( .A1(n560), .A2(G902), .ZN(n561) );
  NOR2_X1 U656 ( .A1(G953), .A2(n562), .ZN(n615) );
  XNOR2_X1 U657 ( .A(KEYINPUT74), .B(n366), .ZN(n597) );
  INV_X1 U658 ( .A(n619), .ZN(n563) );
  OR2_X1 U659 ( .A1(n597), .A2(n563), .ZN(n564) );
  NOR2_X1 U660 ( .A1(n636), .A2(n564), .ZN(n577) );
  NAND2_X1 U661 ( .A1(n577), .A2(n641), .ZN(n566) );
  INV_X1 U662 ( .A(n603), .ZN(n567) );
  NAND2_X1 U663 ( .A1(n568), .A2(n567), .ZN(n570) );
  INV_X1 U664 ( .A(KEYINPUT81), .ZN(n569) );
  XNOR2_X1 U665 ( .A(KEYINPUT65), .B(KEYINPUT19), .ZN(n571) );
  NAND2_X1 U666 ( .A1(n717), .A2(n645), .ZN(n572) );
  XNOR2_X1 U667 ( .A(n572), .B(KEYINPUT47), .ZN(n573) );
  NAND2_X1 U668 ( .A1(n573), .A2(KEYINPUT76), .ZN(n576) );
  NAND2_X1 U669 ( .A1(n645), .A2(KEYINPUT47), .ZN(n574) );
  INV_X1 U670 ( .A(KEYINPUT76), .ZN(n590) );
  NAND2_X1 U671 ( .A1(n574), .A2(n590), .ZN(n575) );
  NAND2_X1 U672 ( .A1(n576), .A2(n575), .ZN(n602) );
  XNOR2_X1 U673 ( .A(KEYINPUT108), .B(n601), .ZN(n719) );
  INV_X1 U674 ( .A(n377), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n580), .A2(n604), .ZN(n675) );
  NAND2_X1 U676 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U677 ( .A(n583), .B(KEYINPUT107), .ZN(n632) );
  NAND2_X1 U678 ( .A1(n632), .A2(n584), .ZN(n588) );
  NOR2_X1 U679 ( .A1(n588), .A2(n596), .ZN(n589) );
  XNOR2_X1 U680 ( .A(n589), .B(KEYINPUT109), .ZN(n764) );
  NAND2_X1 U681 ( .A1(n675), .A2(n764), .ZN(n592) );
  AND2_X1 U682 ( .A1(n717), .A2(n590), .ZN(n591) );
  NOR2_X1 U683 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U684 ( .A(n595), .B(KEYINPUT42), .ZN(n766) );
  NOR2_X1 U685 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U686 ( .A1(n357), .A2(n432), .ZN(n600) );
  NOR2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U689 ( .A(n607), .B(KEYINPUT43), .ZN(n608) );
  NAND2_X1 U690 ( .A1(n609), .A2(n721), .ZN(n724) );
  AND2_X1 U691 ( .A1(n753), .A2(KEYINPUT2), .ZN(n660) );
  NOR2_X1 U692 ( .A1(G898), .A2(n754), .ZN(n612) );
  XNOR2_X1 U693 ( .A(KEYINPUT89), .B(n612), .ZN(n703) );
  NOR2_X1 U694 ( .A1(n613), .A2(n703), .ZN(n614) );
  OR2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U696 ( .A(n620), .B(KEYINPUT104), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n644), .A2(n621), .ZN(n623) );
  INV_X1 U698 ( .A(KEYINPUT22), .ZN(n622) );
  XNOR2_X2 U699 ( .A(n623), .B(n622), .ZN(n627) );
  INV_X1 U700 ( .A(KEYINPUT105), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n636), .A2(n625), .ZN(n626) );
  XNOR2_X1 U702 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT64), .ZN(n629) );
  INV_X1 U704 ( .A(n644), .ZN(n630) );
  INV_X1 U705 ( .A(KEYINPUT34), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n655), .A2(n652), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n633), .A2(KEYINPUT44), .ZN(n649) );
  XNOR2_X1 U708 ( .A(n635), .B(KEYINPUT79), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n707) );
  NAND2_X1 U710 ( .A1(n444), .A2(n638), .ZN(n640) );
  XOR2_X1 U711 ( .A(KEYINPUT31), .B(KEYINPUT97), .Z(n639) );
  XNOR2_X1 U712 ( .A(n640), .B(n639), .ZN(n722) );
  NOR2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U714 ( .A1(n444), .A2(n643), .ZN(n710) );
  OR2_X1 U715 ( .A1(n722), .A2(n710), .ZN(n646) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n647) );
  AND2_X1 U717 ( .A1(n707), .A2(n647), .ZN(n648) );
  NAND2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n651) );
  INV_X1 U719 ( .A(KEYINPUT80), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(n657) );
  BUF_X1 U721 ( .A(n652), .Z(n671) );
  INV_X1 U722 ( .A(KEYINPUT44), .ZN(n653) );
  AND2_X1 U723 ( .A1(n671), .A2(n653), .ZN(n654) );
  NAND2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  INV_X1 U726 ( .A(n358), .ZN(n659) );
  INV_X1 U727 ( .A(n659), .ZN(n697) );
  AND2_X1 U728 ( .A1(n660), .A2(n697), .ZN(n686) );
  NOR2_X1 U729 ( .A1(n358), .A2(KEYINPUT2), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(KEYINPUT77), .ZN(n663) );
  OR2_X1 U731 ( .A1(KEYINPUT2), .A2(n753), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n667), .B(KEYINPUT117), .ZN(n668) );
  XNOR2_X1 U735 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n669) );
  XOR2_X1 U736 ( .A(G122), .B(n672), .Z(G24) );
  XNOR2_X1 U737 ( .A(n673), .B(n411), .ZN(G12) );
  XOR2_X1 U738 ( .A(G125), .B(KEYINPUT37), .Z(n674) );
  XNOR2_X1 U739 ( .A(n675), .B(n674), .ZN(G27) );
  XOR2_X1 U740 ( .A(G119), .B(KEYINPUT127), .Z(n676) );
  INV_X1 U741 ( .A(n684), .ZN(n677) );
  NAND2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  INV_X1 U743 ( .A(KEYINPUT70), .ZN(n680) );
  XNOR2_X1 U744 ( .A(n753), .B(n680), .ZN(n681) );
  INV_X1 U745 ( .A(n681), .ZN(n682) );
  INV_X1 U746 ( .A(KEYINPUT2), .ZN(n683) );
  OR2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U748 ( .A1(n727), .A2(n688), .ZN(n692) );
  XOR2_X1 U749 ( .A(KEYINPUT84), .B(KEYINPUT62), .Z(n689) );
  XNOR2_X1 U750 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U751 ( .A(n692), .B(n691), .ZN(n694) );
  INV_X1 U752 ( .A(G952), .ZN(n693) );
  NOR2_X1 U753 ( .A1(n694), .A2(n750), .ZN(n696) );
  XOR2_X1 U754 ( .A(KEYINPUT82), .B(KEYINPUT63), .Z(n695) );
  XNOR2_X1 U755 ( .A(n696), .B(n695), .ZN(G57) );
  NAND2_X1 U756 ( .A1(n697), .A2(n754), .ZN(n701) );
  NAND2_X1 U757 ( .A1(G953), .A2(G224), .ZN(n698) );
  XNOR2_X1 U758 ( .A(KEYINPUT61), .B(n698), .ZN(n699) );
  NAND2_X1 U759 ( .A1(n699), .A2(G898), .ZN(n700) );
  NAND2_X1 U760 ( .A1(n701), .A2(n700), .ZN(n706) );
  INV_X1 U761 ( .A(n703), .ZN(n704) );
  NOR2_X1 U762 ( .A1(n702), .A2(n704), .ZN(n705) );
  XNOR2_X1 U763 ( .A(n706), .B(n705), .ZN(G69) );
  XNOR2_X1 U764 ( .A(G101), .B(n707), .ZN(G3) );
  XOR2_X1 U765 ( .A(G104), .B(KEYINPUT111), .Z(n709) );
  NAND2_X1 U766 ( .A1(n710), .A2(n719), .ZN(n708) );
  XNOR2_X1 U767 ( .A(n709), .B(n708), .ZN(G6) );
  XOR2_X1 U768 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n712) );
  NAND2_X1 U769 ( .A1(n710), .A2(n721), .ZN(n711) );
  XNOR2_X1 U770 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U771 ( .A(G107), .B(n713), .ZN(G9) );
  XOR2_X1 U772 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n715) );
  NAND2_X1 U773 ( .A1(n717), .A2(n721), .ZN(n714) );
  XNOR2_X1 U774 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U775 ( .A(G128), .B(n716), .ZN(G30) );
  NAND2_X1 U776 ( .A1(n717), .A2(n719), .ZN(n718) );
  XNOR2_X1 U777 ( .A(n718), .B(G146), .ZN(G48) );
  NAND2_X1 U778 ( .A1(n719), .A2(n722), .ZN(n720) );
  XNOR2_X1 U779 ( .A(n720), .B(G113), .ZN(G15) );
  NAND2_X1 U780 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U781 ( .A(n723), .B(G116), .ZN(G18) );
  XNOR2_X1 U782 ( .A(G134), .B(n724), .ZN(G36) );
  XNOR2_X1 U783 ( .A(n725), .B(G140), .ZN(n726) );
  XNOR2_X1 U784 ( .A(n726), .B(KEYINPUT113), .ZN(G42) );
  XOR2_X1 U785 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n729) );
  XNOR2_X1 U786 ( .A(KEYINPUT83), .B(KEYINPUT75), .ZN(n728) );
  XNOR2_X1 U787 ( .A(n729), .B(n728), .ZN(n731) );
  NAND2_X1 U788 ( .A1(n375), .A2(G469), .ZN(n736) );
  XNOR2_X1 U789 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n732) );
  XNOR2_X1 U790 ( .A(n732), .B(KEYINPUT57), .ZN(n733) );
  XNOR2_X1 U791 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U792 ( .A1(n375), .A2(G475), .ZN(n740) );
  XNOR2_X1 U793 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U794 ( .A(KEYINPUT60), .B(KEYINPUT66), .ZN(n742) );
  NAND2_X1 U795 ( .A1(n374), .A2(G478), .ZN(n744) );
  XOR2_X1 U796 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n743) );
  NOR2_X1 U797 ( .A1(n750), .A2(n746), .ZN(G63) );
  NAND2_X1 U798 ( .A1(n374), .A2(G217), .ZN(n747) );
  XNOR2_X1 U799 ( .A(n748), .B(n747), .ZN(n749) );
  NOR2_X1 U800 ( .A1(n750), .A2(n749), .ZN(G66) );
  XNOR2_X1 U801 ( .A(n757), .B(KEYINPUT123), .ZN(n752) );
  XNOR2_X1 U802 ( .A(n753), .B(n752), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U804 ( .A(KEYINPUT124), .B(n756), .ZN(n763) );
  XNOR2_X1 U805 ( .A(n757), .B(G227), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(G900), .ZN(n759) );
  XOR2_X1 U807 ( .A(KEYINPUT125), .B(n759), .Z(n760) );
  NAND2_X1 U808 ( .A1(G953), .A2(n760), .ZN(n761) );
  XNOR2_X1 U809 ( .A(KEYINPUT126), .B(n761), .ZN(n762) );
  NAND2_X1 U810 ( .A1(n763), .A2(n762), .ZN(G72) );
  XNOR2_X1 U811 ( .A(G143), .B(n764), .ZN(G45) );
  XOR2_X1 U812 ( .A(n765), .B(G131), .Z(G33) );
  XOR2_X1 U813 ( .A(G137), .B(n766), .Z(G39) );
endmodule

