//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957;
  OR2_X1    g000(.A1(G15gat), .A2(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G15gat), .A2(G22gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT89), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT16), .B1(new_n202), .B2(new_n203), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n206), .A2(G1gat), .A3(G8gat), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n209));
  INV_X1    g008(.A(new_n203), .ZN(new_n210));
  NOR2_X1   g009(.A1(G15gat), .A2(G22gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G1gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n208), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n205), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(G8gat), .B1(new_n206), .B2(G1gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n213), .A3(new_n208), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT89), .A4(new_n204), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT17), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT87), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(G29gat), .A3(G36gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G29gat), .A2(G36gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT87), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NOR3_X1   g025(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n222), .B(new_n224), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G50gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G43gat), .ZN(new_n230));
  INV_X1    g029(.A(G43gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G50gat), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT15), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT88), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(KEYINPUT88), .A3(new_n233), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G43gat), .B(G50gat), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n239), .A2(KEYINPUT15), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n226), .A2(new_n227), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(KEYINPUT15), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n224), .A2(new_n222), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n240), .A2(new_n241), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n220), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n228), .A2(KEYINPUT88), .A3(new_n233), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT88), .B1(new_n228), .B2(new_n233), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n220), .B(new_n244), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n219), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n219), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n244), .B1(new_n246), .B2(new_n247), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G229gat), .A2(G233gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT18), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n228), .A2(new_n233), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n236), .A2(new_n237), .B1(new_n240), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n219), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n254), .B(KEYINPUT13), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n259), .A2(new_n219), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n252), .A2(KEYINPUT17), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n248), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n267), .B2(new_n219), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(KEYINPUT18), .A3(new_n254), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n257), .A2(new_n264), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT11), .B(G169gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(G197gat), .ZN(new_n272));
  XOR2_X1   g071(.A(G113gat), .B(G141gat), .Z(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT12), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n257), .A2(new_n269), .A3(new_n275), .A4(new_n264), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT86), .ZN(new_n281));
  XOR2_X1   g080(.A(G1gat), .B(G29gat), .Z(new_n282));
  XNOR2_X1  g081(.A(G57gat), .B(G85gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g085(.A(G148gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(G141gat), .ZN(new_n288));
  INV_X1    g087(.A(G141gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(G148gat), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT74), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT2), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n292), .B1(G155gat), .B2(G162gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(G148gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n287), .A2(G141gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT75), .B1(new_n300), .B2(new_n292), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n291), .A2(new_n295), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G155gat), .B(G162gat), .Z(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n293), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT76), .B(G148gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n296), .B1(new_n306), .B2(new_n289), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT3), .ZN(new_n310));
  INV_X1    g109(.A(G120gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G113gat), .ZN(new_n312));
  INV_X1    g111(.A(G113gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G120gat), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT1), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G127gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G113gat), .B(G120gat), .ZN(new_n318));
  OAI21_X1  g117(.A(G127gat), .B1(new_n318), .B2(KEYINPUT1), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G134gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n319), .A3(G134gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n302), .A2(new_n303), .B1(new_n307), .B2(new_n305), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n323), .A3(new_n322), .ZN(new_n329));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT77), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n317), .A2(new_n319), .A3(G134gat), .ZN(new_n335));
  AOI21_X1  g134(.A(G134gat), .B1(new_n317), .B2(new_n319), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n337), .B2(new_n325), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n328), .B(new_n332), .C1(new_n333), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT5), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n309), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n329), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n342), .B2(new_n331), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n331), .A2(KEYINPUT5), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n328), .B(new_n345), .C1(new_n333), .C2(new_n338), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n286), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n346), .ZN(new_n350));
  INV_X1    g149(.A(new_n286), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n344), .A2(new_n286), .A3(new_n346), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n349), .B1(new_n354), .B2(new_n348), .ZN(new_n355));
  INV_X1    g154(.A(G218gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G197gat), .B(G204gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT71), .B(G218gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(new_n358), .B2(KEYINPUT22), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G211gat), .ZN(new_n360));
  INV_X1    g159(.A(G211gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(KEYINPUT22), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n356), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n360), .A2(new_n356), .A3(new_n362), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G226gat), .ZN(new_n367));
  INV_X1    g166(.A(G233gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n372), .A2(new_n373), .B1(G169gat), .B2(G176gat), .ZN(new_n374));
  INV_X1    g173(.A(G183gat), .ZN(new_n375));
  INV_X1    g174(.A(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI211_X1 g176(.A(KEYINPUT65), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT65), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT66), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(KEYINPUT25), .B(new_n374), .C1(new_n382), .C2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n387));
  INV_X1    g186(.A(new_n374), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n377), .A2(new_n383), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(new_n379), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n387), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n370), .A2(KEYINPUT26), .ZN(new_n393));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n370), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT67), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT27), .B(G183gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT28), .B1(new_n401), .B2(G190gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT28), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n403), .A3(new_n376), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT67), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n399), .A2(new_n402), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n392), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n369), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n369), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n392), .B2(new_n406), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n366), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT72), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n407), .A2(new_n369), .ZN(new_n414));
  INV_X1    g213(.A(new_n366), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n392), .B2(new_n406), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n414), .B(new_n415), .C1(new_n369), .C2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n409), .A2(new_n411), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(KEYINPUT72), .A3(new_n415), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  INV_X1    g222(.A(G64gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(G92gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(new_n422), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n427), .B(KEYINPUT73), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n418), .A2(new_n420), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT30), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n427), .B1(new_n418), .B2(new_n420), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n355), .A2(new_n434), .A3(KEYINPUT85), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT85), .B1(new_n355), .B2(new_n434), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n337), .B1(new_n392), .B2(new_n406), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G227gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(new_n368), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n392), .A2(new_n337), .A3(new_n406), .ZN(new_n443));
  NAND2_X1  g242(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n439), .A2(new_n442), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n443), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n447), .A2(new_n438), .A3(new_n441), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n441), .B1(new_n447), .B2(new_n438), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT32), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G15gat), .B(G43gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(G71gat), .B(G99gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n455), .B(new_n456), .Z(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n457), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n451), .B(KEYINPUT32), .C1(new_n453), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n450), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n460), .A3(new_n450), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT70), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT70), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n458), .A2(new_n464), .A3(new_n460), .A4(new_n450), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT31), .B(G50gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT80), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(G78gat), .ZN(new_n469));
  INV_X1    g268(.A(G106gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G22gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n327), .A2(new_n408), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT81), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT81), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n327), .A2(new_n476), .A3(new_n408), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n366), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n364), .A2(new_n408), .A3(new_n365), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n326), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n309), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n478), .A2(G228gat), .A3(new_n481), .A4(G233gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n474), .A2(new_n366), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n325), .B1(new_n479), .B2(new_n326), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n473), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n472), .B1(new_n487), .B2(KEYINPUT83), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n482), .A2(new_n473), .A3(new_n486), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n488), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT82), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n489), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n482), .A2(KEYINPUT82), .A3(new_n473), .A4(new_n486), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n472), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT35), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n466), .A2(new_n492), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n281), .B1(new_n437), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n355), .A2(new_n434), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n355), .A2(new_n434), .A3(KEYINPUT85), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n498), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT86), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n461), .B(KEYINPUT69), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n463), .A2(new_n465), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n492), .A4(new_n496), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT35), .B1(new_n509), .B2(new_n500), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n499), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n434), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n328), .B1(new_n333), .B2(new_n338), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n513), .A2(new_n331), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT39), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n342), .A2(new_n331), .ZN(new_n516));
  OR3_X1    g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(KEYINPUT84), .A2(KEYINPUT40), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n514), .A2(new_n515), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n517), .A2(new_n286), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n286), .A3(new_n520), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n518), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n512), .A2(new_n352), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n492), .A2(new_n496), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT37), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT38), .B1(new_n421), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT37), .B1(new_n418), .B2(new_n420), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n528), .A2(new_n428), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n433), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n527), .B1(new_n412), .B2(new_n417), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT38), .B1(new_n533), .B2(new_n430), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n530), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n524), .B(new_n526), .C1(new_n535), .C2(new_n355), .ZN(new_n536));
  AOI211_X1 g335(.A(KEYINPUT36), .B(new_n461), .C1(new_n463), .C2(new_n465), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n507), .A2(new_n508), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(KEYINPUT36), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n525), .A2(new_n500), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n280), .B1(new_n511), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G57gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G64gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n424), .A2(G57gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT9), .ZN(new_n546));
  NAND2_X1  g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n547), .ZN(new_n549));
  NOR2_X1   g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G71gat), .ZN(new_n553));
  INV_X1    g352(.A(G78gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT91), .B1(new_n555), .B2(new_n547), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n548), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT92), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g358(.A(KEYINPUT92), .B(new_n548), .C1(new_n552), .C2(new_n556), .ZN(new_n560));
  INV_X1    g359(.A(new_n548), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT90), .B1(new_n549), .B2(new_n550), .ZN(new_n562));
  OR3_X1    g361(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT90), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT21), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n219), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G183gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(new_n361), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n574), .B1(new_n570), .B2(new_n571), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n565), .A2(new_n566), .ZN(new_n577));
  XOR2_X1   g376(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OR3_X1    g379(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n575), .B2(new_n576), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n426), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n585), .B2(new_n426), .ZN(new_n588));
  NAND3_X1  g387(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G99gat), .B(G106gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n586), .A2(new_n591), .A3(new_n588), .A4(new_n589), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(KEYINPUT94), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(new_n596), .A3(new_n592), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n267), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G190gat), .B(G218gat), .Z(new_n600));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT93), .Z(new_n602));
  INV_X1    g401(.A(KEYINPUT41), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n595), .A2(new_n597), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n604), .B1(new_n252), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n599), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n603), .ZN(new_n608));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT95), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n600), .B1(new_n599), .B2(new_n606), .ZN(new_n613));
  MUX2_X1   g412(.A(new_n611), .B(new_n610), .S(new_n613), .Z(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n614), .B2(new_n607), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n605), .A2(new_n565), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n593), .A2(new_n594), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n618), .A2(new_n559), .A3(new_n560), .A4(new_n564), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT10), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n598), .A2(new_n621), .A3(new_n565), .ZN(new_n622));
  INV_X1    g421(.A(G230gat), .ZN(new_n623));
  OAI22_X1  g422(.A1(new_n620), .A2(new_n622), .B1(new_n623), .B2(new_n368), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n617), .A2(new_n619), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n623), .A2(new_n368), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  INV_X1    g428(.A(G176gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n628), .B(new_n633), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n583), .A2(new_n616), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n542), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT96), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n542), .A2(new_n638), .A3(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n355), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT97), .B(G1gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(G1324gat));
  NAND2_X1  g443(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n640), .A2(new_n512), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n208), .B1(new_n640), .B2(new_n512), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n648), .B1(new_n652), .B2(new_n650), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n649), .B1(new_n648), .B2(new_n650), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(G1325gat));
  AOI21_X1  g454(.A(G15gat), .B1(new_n640), .B2(new_n466), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n539), .B1(new_n637), .B2(new_n639), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(G15gat), .B2(new_n657), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n640), .A2(new_n525), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT43), .B(G22gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  INV_X1    g460(.A(new_n583), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n634), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n615), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n542), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n666), .A2(G29gat), .A3(new_n355), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT45), .Z(new_n668));
  AOI21_X1  g467(.A(new_n615), .B1(new_n511), .B2(new_n541), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT18), .B1(new_n268), .B2(new_n254), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n251), .B1(new_n266), .B2(new_n248), .ZN(new_n673));
  INV_X1    g472(.A(new_n254), .ZN(new_n674));
  NOR4_X1   g473(.A1(new_n673), .A2(new_n256), .A3(new_n265), .A4(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n275), .B1(new_n676), .B2(new_n264), .ZN(new_n677));
  INV_X1    g476(.A(new_n278), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT99), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n277), .A2(new_n680), .A3(new_n278), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n664), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n671), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(G29gat), .B1(new_n685), .B2(new_n355), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n686), .ZN(G1328gat));
  OR3_X1    g486(.A1(new_n666), .A2(G36gat), .A3(new_n434), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n688), .A2(KEYINPUT100), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(KEYINPUT100), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT46), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G36gat), .B1(new_n685), .B2(new_n434), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n689), .B2(new_n690), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(G1329gat));
  NAND2_X1  g494(.A1(new_n511), .A2(new_n541), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n616), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n670), .ZN(new_n698));
  INV_X1    g497(.A(new_n539), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n669), .A2(KEYINPUT44), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .A4(new_n684), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G43gat), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n542), .A2(new_n231), .A3(new_n466), .A4(new_n665), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(KEYINPUT47), .A3(new_n703), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n701), .A2(KEYINPUT102), .A3(G43gat), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT102), .B1(new_n701), .B2(G43gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n703), .B(KEYINPUT103), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT101), .B(KEYINPUT47), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n704), .B1(new_n708), .B2(new_n709), .ZN(G1330gat));
  NAND3_X1  g509(.A1(new_n671), .A2(new_n525), .A3(new_n684), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G50gat), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT48), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n542), .A2(new_n229), .A3(new_n525), .A4(new_n665), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n712), .B(new_n715), .C1(new_n713), .C2(KEYINPUT48), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1331gat));
  AOI211_X1 g518(.A(new_n583), .B(new_n616), .C1(new_n511), .C2(new_n541), .ZN(new_n720));
  INV_X1    g519(.A(new_n634), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n682), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n355), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT105), .B(G57gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1332gat));
  NOR2_X1   g525(.A1(new_n723), .A2(new_n434), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(G1333gat));
  NAND4_X1  g530(.A1(new_n720), .A2(G71gat), .A3(new_n699), .A4(new_n722), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT106), .Z(new_n733));
  INV_X1    g532(.A(new_n466), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n553), .B1(new_n723), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT50), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n733), .A2(new_n738), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1334gat));
  NOR2_X1   g539(.A1(new_n723), .A2(new_n526), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(new_n554), .ZN(G1335gat));
  NAND2_X1  g541(.A1(new_n583), .A2(new_n683), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT107), .Z(new_n744));
  NAND4_X1  g543(.A1(new_n698), .A2(new_n634), .A3(new_n700), .A4(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n745), .A2(new_n585), .A3(new_n355), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n696), .A2(new_n616), .A3(new_n744), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT51), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n669), .A2(new_n749), .A3(new_n744), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(new_n641), .A3(new_n634), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n746), .B1(new_n585), .B2(new_n752), .ZN(G1336gat));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  OAI21_X1  g553(.A(G92gat), .B1(new_n745), .B2(new_n434), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(KEYINPUT108), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n751), .A2(new_n426), .A3(new_n512), .A4(new_n634), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n755), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n757), .B(new_n755), .C1(KEYINPUT108), .C2(new_n754), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1337gat));
  OAI21_X1  g560(.A(G99gat), .B1(new_n745), .B2(new_n539), .ZN(new_n762));
  INV_X1    g561(.A(G99gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n751), .A2(new_n763), .A3(new_n634), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n764), .B2(new_n734), .ZN(G1338gat));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n748), .A2(new_n525), .A3(new_n634), .A4(new_n750), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n470), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n671), .A2(new_n525), .A3(new_n634), .A4(new_n744), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n470), .B1(new_n770), .B2(KEYINPUT109), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n766), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT109), .B1(new_n745), .B2(new_n526), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G106gat), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n770), .A2(new_n769), .ZN(new_n776));
  OAI211_X1 g575(.A(KEYINPUT53), .B(new_n775), .C1(new_n776), .C2(new_n768), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n773), .A2(new_n777), .ZN(G1339gat));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  INV_X1    g578(.A(new_n565), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n626), .B(new_n781), .C1(new_n625), .C2(KEYINPUT10), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n624), .A3(KEYINPUT54), .ZN(new_n783));
  XOR2_X1   g582(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n784));
  OAI221_X1 g583(.A(new_n784), .B1(new_n623), .B2(new_n368), .C1(new_n620), .C2(new_n622), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n783), .A2(KEYINPUT55), .A3(new_n633), .A4(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n628), .A2(new_n633), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n785), .A2(new_n633), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT55), .B1(new_n789), .B2(new_n783), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n277), .A2(new_n680), .A3(new_n278), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n680), .B1(new_n277), .B2(new_n278), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n268), .B2(new_n254), .ZN(new_n796));
  OAI211_X1 g595(.A(KEYINPUT111), .B(new_n674), .C1(new_n673), .C2(new_n265), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n253), .A2(new_n260), .A3(new_n262), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT112), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n274), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n634), .A2(new_n801), .A3(new_n278), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n616), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n791), .A2(new_n278), .A3(new_n801), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n615), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n779), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n616), .A2(new_n278), .A3(new_n801), .A4(new_n791), .ZN(new_n807));
  INV_X1    g606(.A(new_n802), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n682), .B2(new_n791), .ZN(new_n809));
  OAI211_X1 g608(.A(KEYINPUT113), .B(new_n807), .C1(new_n809), .C2(new_n616), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n810), .A3(new_n583), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n635), .A2(new_n683), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n526), .A2(new_n466), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n512), .A2(new_n355), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G113gat), .B1(new_n820), .B2(new_n280), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n525), .B(new_n538), .C1(new_n811), .C2(new_n812), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n817), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n313), .A3(new_n682), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(G1340gat));
  OAI21_X1  g624(.A(G120gat), .B1(new_n820), .B2(new_n721), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n311), .A3(new_n634), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1341gat));
  NOR3_X1   g627(.A1(new_n820), .A2(new_n316), .A3(new_n583), .ZN(new_n829));
  AOI21_X1  g628(.A(G127gat), .B1(new_n823), .B2(new_n662), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(G1342gat));
  NAND3_X1  g630(.A1(new_n822), .A2(new_n321), .A3(new_n817), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n832), .A2(KEYINPUT56), .A3(new_n615), .ZN(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n820), .B2(new_n615), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT56), .B1(new_n832), .B2(new_n615), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT114), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n789), .A2(new_n783), .ZN(new_n838));
  XOR2_X1   g637(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n840), .A2(new_n279), .A3(new_n787), .A4(new_n786), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n842), .A3(new_n802), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n841), .B2(new_n802), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n615), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n848), .B(new_n615), .C1(new_n844), .C2(new_n845), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n807), .A3(new_n849), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n850), .A2(new_n583), .B1(new_n635), .B2(new_n683), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT57), .B1(new_n851), .B2(new_n526), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n526), .B1(new_n811), .B2(new_n812), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n699), .A2(new_n818), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G141gat), .B1(new_n857), .B2(new_n280), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n853), .A2(new_n856), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n289), .A3(new_n279), .ZN(new_n860));
  XOR2_X1   g659(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n860), .ZN(new_n863));
  INV_X1    g662(.A(new_n857), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n682), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(G141gat), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(G1344gat));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n855), .A3(new_n634), .A4(new_n856), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n870), .A3(new_n306), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT120), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n841), .A2(new_n802), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT116), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n616), .B1(new_n874), .B2(new_n843), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n583), .B1(new_n875), .B2(new_n805), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n635), .A2(new_n280), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n876), .A2(KEYINPUT121), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT121), .B1(new_n876), .B2(new_n877), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n854), .B(new_n525), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n853), .A2(new_n854), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n880), .A2(new_n634), .A3(new_n856), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G148gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT59), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n885), .A3(new_n870), .A4(new_n306), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n872), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n306), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n859), .A2(new_n888), .A3(new_n634), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT119), .Z(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n890), .ZN(G1345gat));
  AOI21_X1  g690(.A(G155gat), .B1(new_n859), .B2(new_n662), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n662), .A2(G155gat), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT122), .Z(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n864), .B2(new_n894), .ZN(G1346gat));
  AOI21_X1  g694(.A(G162gat), .B1(new_n859), .B2(new_n616), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n857), .A2(new_n615), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n641), .A2(new_n434), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT123), .B1(new_n816), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n814), .B1(new_n811), .B2(new_n812), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n903), .A3(new_n899), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n280), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n822), .A2(new_n899), .ZN(new_n907));
  INV_X1    g706(.A(G169gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n908), .A3(new_n682), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(new_n909), .ZN(G1348gat));
  NOR3_X1   g709(.A1(new_n905), .A2(new_n630), .A3(new_n721), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n913));
  AOI21_X1  g712(.A(G176gat), .B1(new_n907), .B2(new_n634), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G1349gat));
  NAND3_X1  g714(.A1(new_n907), .A2(new_n400), .A3(new_n662), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n905), .A2(new_n583), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n375), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n902), .A2(new_n903), .A3(new_n899), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n903), .B1(new_n902), .B2(new_n899), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n921), .A2(new_n922), .A3(new_n615), .ZN(new_n923));
  OAI211_X1 g722(.A(KEYINPUT125), .B(new_n920), .C1(new_n923), .C2(new_n376), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n376), .A3(new_n616), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n901), .A2(new_n616), .A3(new_n904), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n926), .A2(G190gat), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n924), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n924), .A2(KEYINPUT126), .A3(new_n925), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1351gat));
  NOR2_X1   g733(.A1(new_n699), .A2(new_n900), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n853), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(G197gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n937), .A3(new_n682), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n880), .A2(new_n881), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n939), .A2(new_n935), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n940), .A2(new_n279), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n941), .B2(new_n937), .ZN(G1352gat));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n634), .A3(new_n935), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT127), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n939), .A2(new_n945), .A3(new_n634), .A4(new_n935), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(G204gat), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n936), .A2(new_n632), .A3(new_n634), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1353gat));
  NAND3_X1  g749(.A1(new_n936), .A2(new_n361), .A3(new_n662), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n939), .A2(new_n662), .A3(new_n935), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(G1354gat));
  AOI21_X1  g754(.A(G218gat), .B1(new_n936), .B2(new_n616), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n616), .A2(new_n358), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n940), .B2(new_n957), .ZN(G1355gat));
endmodule


