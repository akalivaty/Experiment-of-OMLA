//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT66), .B(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT67), .B(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT68), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT69), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT71), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT70), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n458), .B1(new_n464), .B2(G101), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  AOI211_X1 g041(.A(KEYINPUT71), .B(new_n466), .C1(new_n461), .C2(new_n463), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n476), .B2(new_n462), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n468), .A2(new_n477), .ZN(G160));
  AOI21_X1  g053(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(G136), .B2(new_n471), .ZN(G162));
  OR2_X1    g059(.A1(new_n462), .A2(G114), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n479), .A2(G126), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n489), .B1(new_n494), .B2(KEYINPUT73), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n489), .A2(KEYINPUT72), .A3(KEYINPUT73), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n475), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(KEYINPUT72), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n488), .A2(new_n495), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(KEYINPUT75), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n506), .A2(new_n509), .A3(G62), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n501), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT74), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(KEYINPUT74), .A2(KEYINPUT6), .A3(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n503), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n515), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(new_n506), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n511), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n525), .B(new_n527), .C1(new_n528), .C2(new_n520), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n516), .B(KEYINPUT77), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n529), .B1(G51), .B2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n530), .A2(G52), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n501), .ZN(new_n534));
  AND2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n514), .B2(new_n515), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G90), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n532), .A2(new_n534), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(new_n530), .A2(G43), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n538), .A2(G81), .B1(new_n545), .B2(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT78), .Z(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g126(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n552));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n516), .A2(G53), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n516), .A2(new_n558), .A3(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n538), .A2(G91), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT81), .B(G65), .Z(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(new_n537), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT80), .Z(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n560), .A2(new_n561), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(new_n529), .ZN(new_n568));
  INV_X1    g143(.A(G51), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n516), .B(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n568), .B1(new_n569), .B2(new_n571), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  NAND3_X1  g148(.A1(new_n519), .A2(G87), .A3(new_n506), .ZN(new_n574));
  INV_X1    g149(.A(new_n515), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT6), .B1(KEYINPUT74), .B2(G651), .ZN(new_n576));
  OAI211_X1 g151(.A(G49), .B(G543), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n504), .A2(new_n578), .A3(new_n505), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n574), .A2(new_n577), .A3(new_n580), .ZN(G288));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  INV_X1    g157(.A(G73), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n537), .A2(new_n582), .B1(new_n583), .B2(new_n503), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(G48), .B2(new_n516), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n519), .A2(G86), .A3(new_n506), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n538), .A2(G85), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI221_X1 g165(.A(new_n588), .B1(new_n501), .B2(new_n589), .C1(new_n571), .C2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n538), .A2(KEYINPUT10), .A3(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n520), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n537), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n593), .A2(new_n596), .B1(G651), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n530), .A2(G54), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n592), .B1(new_n602), .B2(G868), .ZN(G284));
  XNOR2_X1  g178(.A(G284), .B(KEYINPUT82), .ZN(G321));
  XNOR2_X1  g179(.A(G299), .B(KEYINPUT83), .ZN(new_n605));
  MUX2_X1   g180(.A(new_n605), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g181(.A(new_n605), .B(G286), .S(G868), .Z(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n602), .B1(new_n608), .B2(G860), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT84), .ZN(G148));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n608), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  INV_X1    g190(.A(G111), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G2105), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n471), .A2(G135), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT85), .Z(new_n619));
  AOI211_X1 g194(.A(new_n617), .B(new_n619), .C1(G123), .C2(new_n479), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2096), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n464), .A2(new_n475), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT13), .Z(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n621), .A2(new_n626), .A3(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n629), .B(new_n630), .Z(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT87), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n634), .A2(new_n635), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n641), .B1(new_n638), .B2(new_n639), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n632), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n646), .A2(new_n631), .A3(new_n642), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G14), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n648), .B1(new_n645), .B2(new_n647), .ZN(new_n651));
  OAI21_X1  g226(.A(KEYINPUT88), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n651), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n654));
  NAND4_X1  g229(.A1(new_n653), .A2(new_n654), .A3(G14), .A4(new_n649), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT17), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT90), .ZN(new_n666));
  INV_X1    g241(.A(new_n664), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n658), .A2(new_n660), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n667), .B(new_n668), .C1(new_n659), .C2(new_n661), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n658), .A3(new_n660), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G2100), .ZN(new_n674));
  NAND4_X1  g249(.A1(new_n666), .A2(new_n625), .A3(new_n669), .A4(new_n672), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT91), .B(G2096), .ZN(new_n676));
  AND3_X1   g251(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n676), .B1(new_n674), .B2(new_n675), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT93), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  OR3_X1    g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n688), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n685), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n685), .A2(new_n689), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n690), .A2(new_n693), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G1981), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n697), .B(G1981), .ZN(new_n701));
  INV_X1    g276(.A(G1986), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n682), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n700), .A2(new_n703), .A3(new_n682), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n706), .ZN(new_n709));
  INV_X1    g284(.A(new_n707), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n704), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n708), .A2(new_n711), .ZN(G229));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G21), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G168), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G1966), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT102), .ZN(new_n717));
  NOR2_X1   g292(.A1(G171), .A2(new_n713), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G5), .B2(new_n713), .ZN(new_n719));
  INV_X1    g294(.A(G1961), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n715), .A2(G1966), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT31), .B(G11), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT30), .B(G28), .Z(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G29), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n620), .B2(G29), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n721), .A2(new_n722), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT103), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n717), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n713), .A2(G20), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT23), .ZN(new_n731));
  INV_X1    g306(.A(G299), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n713), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1956), .ZN(new_n734));
  NOR2_X1   g309(.A1(G29), .A2(G35), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G162), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT104), .B(KEYINPUT29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2090), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n740));
  NAND2_X1  g315(.A1(G103), .A2(G2104), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G2105), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n471), .A2(G139), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n462), .B2(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G33), .B(new_n746), .S(G29), .Z(new_n747));
  AOI21_X1  g322(.A(new_n739), .B1(G2072), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT100), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT26), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  AOI22_X1  g327(.A1(G129), .A2(new_n479), .B1(new_n471), .B2(G141), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n464), .A2(G105), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n757), .B2(G32), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n747), .A2(G2072), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT99), .ZN(new_n763));
  INV_X1    g338(.A(G34), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n764), .A2(KEYINPUT24), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(KEYINPUT24), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n757), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G160), .B2(new_n757), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G2084), .Z(new_n769));
  NAND4_X1  g344(.A1(new_n748), .A2(new_n761), .A3(new_n763), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n759), .A2(new_n760), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(KEYINPUT101), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(KEYINPUT101), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n734), .B(new_n770), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n757), .A2(G26), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT28), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n479), .A2(G128), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n780));
  INV_X1    g355(.A(G116), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(G2105), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G140), .B2(new_n471), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT98), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n776), .B1(new_n786), .B2(new_n757), .ZN(new_n787));
  INV_X1    g362(.A(G2067), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n713), .A2(G4), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n602), .B2(new_n713), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1348), .Z(new_n792));
  INV_X1    g367(.A(G1341), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n547), .A2(G16), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n713), .A2(G19), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n719), .A2(new_n720), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n757), .A2(G27), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n757), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2078), .ZN(new_n800));
  INV_X1    g375(.A(new_n796), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(G1341), .ZN(new_n802));
  AND4_X1   g377(.A1(new_n789), .A2(new_n792), .A3(new_n797), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n728), .B1(new_n717), .B2(new_n727), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n729), .A2(new_n774), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n713), .A2(G6), .ZN(new_n806));
  INV_X1    g381(.A(G305), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n713), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT96), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT32), .B(G1981), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n713), .A2(G22), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G166), .B2(new_n713), .ZN(new_n813));
  INV_X1    g388(.A(G1971), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  MUX2_X1   g390(.A(G23), .B(G288), .S(G16), .Z(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT33), .B(G1976), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  OR3_X1    g394(.A1(new_n811), .A2(KEYINPUT34), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT34), .B1(new_n811), .B2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n479), .A2(G119), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n825));
  INV_X1    g400(.A(G107), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(G2105), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G131), .B2(new_n471), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  MUX2_X1   g404(.A(G25), .B(new_n829), .S(G29), .Z(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT35), .B(G1991), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT95), .Z(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n830), .B(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n713), .A2(G24), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G290), .B2(G16), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n834), .B1(new_n702), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n702), .B2(new_n836), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n820), .A2(new_n821), .A3(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n805), .B1(new_n840), .B2(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  INV_X1    g418(.A(new_n805), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(G150));
  NAND2_X1  g420(.A1(new_n602), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n537), .B2(new_n849), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n538), .A2(G93), .B1(new_n850), .B2(G651), .ZN(new_n851));
  INV_X1    g426(.A(G55), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n571), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n547), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n530), .A2(G55), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n542), .A2(new_n855), .A3(new_n546), .A4(new_n851), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n847), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT105), .Z(new_n861));
  AOI21_X1  g436(.A(G860), .B1(new_n858), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n853), .A2(G860), .ZN(new_n864));
  XOR2_X1   g439(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(G145));
  XOR2_X1   g442(.A(G160), .B(G162), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT107), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(new_n620), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n620), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n784), .B(KEYINPUT98), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n499), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n786), .A2(G164), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT108), .ZN(new_n877));
  INV_X1    g452(.A(G118), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n876), .A2(new_n877), .B1(new_n878), .B2(G2105), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n877), .B2(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n471), .A2(G142), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n479), .A2(G130), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n874), .A2(new_n875), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n829), .B(new_n623), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n756), .B(new_n746), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n883), .B1(new_n874), .B2(new_n875), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n885), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n874), .A2(new_n875), .ZN(new_n893));
  INV_X1    g468(.A(new_n883), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n895), .A2(new_n884), .B1(new_n889), .B2(new_n888), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n872), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n890), .B1(new_n885), .B2(new_n891), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n895), .A2(new_n884), .A3(new_n889), .A4(new_n888), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n871), .A4(new_n870), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g478(.A(G290), .B(G305), .ZN(new_n904));
  XNOR2_X1  g479(.A(G166), .B(G288), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(KEYINPUT42), .Z(new_n907));
  XNOR2_X1  g482(.A(new_n857), .B(new_n611), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n600), .A2(new_n601), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(G299), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n566), .A2(new_n561), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n912), .A2(new_n560), .B1(new_n600), .B2(new_n601), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n911), .B2(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n910), .A2(G299), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n912), .A2(new_n600), .A3(new_n560), .A4(new_n601), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(KEYINPUT41), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n909), .B1(new_n908), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n914), .ZN(new_n923));
  INV_X1    g498(.A(new_n908), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n907), .A2(new_n915), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n907), .B1(new_n925), .B2(new_n915), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n853), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(G868), .B2(new_n929), .ZN(G295));
  OAI21_X1  g505(.A(new_n928), .B1(G868), .B2(new_n929), .ZN(G331));
  INV_X1    g506(.A(new_n906), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n854), .A2(G301), .A3(new_n856), .ZN(new_n933));
  AOI21_X1  g508(.A(G301), .B1(new_n854), .B2(new_n856), .ZN(new_n934));
  OAI21_X1  g509(.A(G286), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n547), .A2(new_n853), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n542), .A2(new_n546), .B1(new_n855), .B2(new_n851), .ZN(new_n937));
  OAI21_X1  g512(.A(G171), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n854), .A2(G301), .A3(new_n856), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(G168), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n935), .A2(new_n921), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n914), .B1(new_n935), .B2(new_n940), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n932), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n933), .A2(new_n934), .A3(G286), .ZN(new_n946));
  AOI21_X1  g521(.A(G168), .B1(new_n938), .B2(new_n939), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n923), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n948), .A2(new_n942), .A3(new_n906), .A4(new_n941), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n901), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT111), .B1(new_n950), .B2(KEYINPUT43), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n948), .A2(new_n942), .A3(new_n941), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n955), .B2(new_n932), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n956), .B2(new_n949), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n951), .A2(new_n952), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n954), .A3(new_n949), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT111), .A4(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(G397));
  NAND2_X1  g537(.A1(new_n786), .A2(new_n788), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n873), .A2(G2067), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n756), .B(G1996), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n829), .B(new_n833), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  OAI211_X1 g544(.A(G126), .B(G2105), .C1(new_n492), .C2(new_n493), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n485), .A2(new_n487), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n498), .A2(new_n497), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n462), .A2(G138), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n469), .B2(new_n470), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT73), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT4), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n969), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT112), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT45), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n492), .A2(new_n493), .ZN(new_n983));
  INV_X1    g558(.A(G125), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n473), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n985), .A2(G2105), .B1(G137), .B2(new_n471), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n986), .B(G40), .C1(new_n465), .C2(new_n467), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n968), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(G290), .A2(G1986), .ZN(new_n990));
  AND2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT113), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT114), .B(G8), .ZN(new_n995));
  INV_X1    g570(.A(G40), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n468), .A2(new_n477), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n995), .B1(new_n978), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n999));
  INV_X1    g574(.A(G1976), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G288), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI211_X1 g578(.A(KEYINPUT115), .B(KEYINPUT52), .C1(G288), .C2(new_n1000), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(G288), .A2(new_n1000), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n998), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT49), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT117), .B(G86), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n519), .A2(new_n506), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n698), .B1(new_n585), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n582), .B1(new_n504), .B2(new_n505), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n583), .A2(new_n503), .ZN(new_n1013));
  OAI21_X1  g588(.A(G651), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n516), .A2(G48), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT116), .B(G1981), .Z(new_n1016));
  AND4_X1   g591(.A1(new_n586), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1008), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(G160), .A2(G40), .A3(new_n969), .A4(new_n499), .ZN(new_n1019));
  INV_X1    g594(.A(new_n995), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n585), .A2(new_n586), .A3(new_n1016), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1014), .A2(new_n1015), .A3(new_n1010), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G1981), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1023), .A3(KEYINPUT49), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1020), .B(new_n1006), .C1(new_n987), .C2(new_n977), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1007), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(G166), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT55), .B(G8), .C1(new_n511), .C2(new_n521), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n499), .B2(new_n969), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(new_n987), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1971), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G2090), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n977), .A2(KEYINPUT50), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n499), .A2(new_n1040), .A3(new_n969), .ZN(new_n1041));
  AND4_X1   g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n997), .A4(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(G8), .B(new_n1033), .C1(new_n1037), .C2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1028), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n977), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(new_n997), .A3(new_n1036), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n814), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1039), .A2(new_n997), .A3(new_n1041), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(G2090), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1033), .B1(new_n1050), .B2(new_n1020), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT125), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1033), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1037), .A2(new_n1042), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n995), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT125), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n1043), .A4(new_n1028), .ZN(new_n1057));
  INV_X1    g632(.A(G2078), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1035), .A2(new_n1058), .A3(new_n1036), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT123), .B(G1961), .Z(new_n1061));
  AOI22_X1  g636(.A1(new_n1059), .A2(new_n1060), .B1(new_n1049), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1036), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1046), .A2(new_n997), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1046), .A2(KEYINPUT120), .A3(new_n997), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1060), .A2(G2078), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1062), .A2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(G301), .B(KEYINPUT54), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT124), .B(G2078), .Z(new_n1072));
  NOR4_X1   g647(.A1(new_n1063), .A2(new_n1060), .A3(new_n987), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1071), .B1(new_n982), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1070), .A2(new_n1071), .B1(new_n1074), .B2(new_n1062), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1052), .A2(new_n1057), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G286), .A2(new_n1020), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1049), .A2(G2084), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1065), .B1(new_n1034), .B2(new_n987), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1067), .A2(new_n1080), .A3(new_n1036), .ZN(new_n1081));
  INV_X1    g656(.A(G1966), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1077), .B(new_n1078), .C1(new_n1083), .C2(new_n995), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1966), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1086));
  OAI21_X1  g661(.A(G8), .B1(new_n1086), .B2(new_n1079), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1077), .B1(new_n1087), .B2(new_n1078), .ZN(new_n1088));
  OAI211_X1 g663(.A(G286), .B(new_n1020), .C1(new_n1086), .C2(new_n1079), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n912), .B(new_n560), .C1(KEYINPUT121), .C2(KEYINPUT57), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n566), .A2(KEYINPUT121), .A3(new_n561), .ZN(new_n1093));
  NAND3_X1  g668(.A1(G299), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n987), .B1(KEYINPUT50), .B2(new_n977), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1956), .B1(new_n1097), .B2(new_n1041), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(G2072), .ZN(new_n1100));
  AND4_X1   g675(.A1(new_n997), .A2(new_n1046), .A3(new_n1036), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1096), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1348), .B1(new_n1097), .B2(new_n1041), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1019), .A2(G2067), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1102), .B1(new_n1105), .B2(new_n910), .ZN(new_n1106));
  INV_X1    g681(.A(G1956), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1049), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1035), .A2(new_n1036), .A3(new_n1100), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n1095), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1108), .A2(new_n1109), .A3(new_n1095), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1095), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1039), .A2(new_n997), .A3(new_n1041), .ZN(new_n1116));
  OAI221_X1 g691(.A(KEYINPUT60), .B1(G2067), .B2(new_n1019), .C1(new_n1116), .C2(G1348), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1119), .A3(new_n602), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1102), .A2(KEYINPUT61), .A3(new_n1110), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1115), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n987), .A2(new_n977), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT58), .B(G1341), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n1047), .A2(G1996), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n548), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(KEYINPUT59), .A3(new_n548), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1128), .B(new_n1129), .C1(new_n602), .C2(new_n1117), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1111), .B1(new_n1122), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1076), .A2(new_n1090), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(G288), .A2(G1976), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1017), .B1(new_n1025), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n998), .B(KEYINPUT118), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1028), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1136), .A2(new_n1138), .B1(new_n1139), .B2(new_n1043), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1083), .A2(new_n995), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(G168), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1055), .A2(new_n1043), .A3(new_n1028), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1044), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1050), .A2(G8), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1141), .B1(new_n1147), .B2(new_n1053), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1146), .A2(new_n1148), .A3(G168), .A4(new_n1142), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1140), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1132), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1078), .B1(new_n1083), .B2(new_n1030), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n1089), .A3(KEYINPUT51), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1153), .A2(new_n1084), .A3(KEYINPUT62), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT62), .B1(new_n1153), .B2(new_n1084), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1052), .A2(new_n1057), .A3(G171), .A4(new_n1070), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n994), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n988), .A2(new_n990), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT48), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1159), .A2(KEYINPUT48), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n989), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n988), .ZN(new_n1163));
  OR3_X1    g738(.A1(new_n1163), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT46), .B1(new_n1163), .B2(G1996), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n963), .A2(new_n964), .A3(new_n756), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1164), .A2(new_n1165), .B1(new_n988), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT47), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1162), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n829), .A2(new_n832), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n966), .B2(new_n1163), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1173), .A2(new_n1174), .A3(new_n963), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1173), .B2(new_n963), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1175), .A2(new_n1176), .A3(new_n1163), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1158), .A2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g754(.A(G319), .B1(new_n677), .B2(new_n678), .ZN(new_n1181));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g757(.A(KEYINPUT127), .B(G319), .C1(new_n677), .C2(new_n678), .ZN(new_n1184));
  AOI22_X1  g758(.A1(new_n708), .A2(new_n711), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g759(.A1(new_n656), .A2(new_n1185), .A3(new_n902), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n1186), .B1(new_n959), .B2(new_n960), .ZN(G308));
  NAND2_X1  g761(.A1(new_n959), .A2(new_n960), .ZN(new_n1188));
  NAND4_X1  g762(.A1(new_n1188), .A2(new_n656), .A3(new_n902), .A4(new_n1185), .ZN(G225));
endmodule


