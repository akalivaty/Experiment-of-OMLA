//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT80), .ZN(new_n193));
  INV_X1    g007(.A(G227), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G953), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n193), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G137), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n199), .A2(new_n201), .A3(new_n205), .A4(new_n202), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT81), .A3(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n212), .A2(new_n208), .A3(KEYINPUT81), .A4(G104), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G107), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n210), .A2(new_n211), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n215), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n214), .A2(G107), .ZN(new_n218));
  OAI21_X1  g032(.A(G101), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n223), .A3(G143), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n224), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT1), .B1(new_n225), .B2(G146), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n224), .A2(new_n226), .B1(G128), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n216), .B(new_n219), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT10), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n225), .A2(G146), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT64), .B(G146), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(G143), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n237), .B2(G143), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n240), .B2(new_n227), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n224), .A2(new_n226), .A3(new_n228), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n233), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n216), .A2(new_n219), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT84), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n227), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n221), .A2(new_n223), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n235), .B1(new_n247), .B2(new_n225), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n242), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(new_n244), .A3(KEYINPUT84), .A4(KEYINPUT10), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n234), .B1(new_n245), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n210), .A2(new_n213), .A3(new_n215), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT82), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT82), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n210), .A2(new_n256), .A3(new_n213), .A4(new_n215), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n254), .A2(new_n255), .A3(G101), .A4(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n224), .A2(new_n259), .A3(new_n226), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n260), .B1(new_n248), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n254), .A2(G101), .A3(new_n257), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n216), .A2(KEYINPUT4), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT83), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n267), .A2(KEYINPUT83), .A3(new_n268), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n266), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n207), .B1(new_n252), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT87), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n249), .A2(new_n244), .A3(KEYINPUT10), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT84), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n278), .A2(new_n250), .B1(new_n233), .B2(new_n232), .ZN(new_n279));
  INV_X1    g093(.A(new_n266), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n267), .A2(KEYINPUT83), .A3(new_n268), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT83), .B1(new_n267), .B2(new_n268), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT87), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n207), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n275), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n207), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n279), .A2(new_n288), .A3(new_n283), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n196), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n216), .A2(new_n219), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n241), .A2(new_n242), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT85), .A3(new_n232), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n241), .A2(new_n291), .A3(new_n294), .A4(new_n242), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n293), .A2(KEYINPUT12), .A3(new_n207), .A4(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT12), .ZN(new_n299));
  INV_X1    g113(.A(new_n293), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n207), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n301), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n303), .A2(KEYINPUT86), .A3(KEYINPUT12), .A4(new_n293), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n298), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n305), .A2(new_n289), .A3(new_n196), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n190), .B(new_n191), .C1(new_n290), .C2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n190), .A2(new_n191), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n196), .B1(new_n305), .B2(new_n289), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n289), .A2(new_n196), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n287), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n308), .B1(new_n311), .B2(G469), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n189), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(G110), .B(G122), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G116), .B(G119), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT2), .B(G113), .Z(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(KEYINPUT65), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT2), .B(G113), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT65), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n317), .A2(KEYINPUT66), .A3(new_n316), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT66), .B1(new_n317), .B2(new_n316), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n258), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(new_n271), .B2(new_n272), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n316), .A2(KEYINPUT5), .ZN(new_n329));
  INV_X1    g143(.A(G116), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n330), .A2(KEYINPUT5), .A3(G119), .ZN(new_n331));
  INV_X1    g145(.A(G113), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n324), .B2(new_n325), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(new_n291), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n315), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n336), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n281), .A2(new_n282), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n314), .B(new_n338), .C1(new_n339), .C2(new_n327), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n340), .A3(KEYINPUT6), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n264), .A2(G125), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(KEYINPUT88), .C1(G125), .C2(new_n249), .ZN(new_n343));
  OR3_X1    g157(.A1(new_n249), .A2(KEYINPUT88), .A3(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G224), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G953), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n345), .B(new_n347), .Z(new_n348));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n315), .C1(new_n328), .C2(new_n336), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n341), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n314), .B(KEYINPUT8), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n317), .A2(new_n316), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT66), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n355), .A2(new_n323), .B1(new_n329), .B2(new_n333), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT89), .A3(new_n244), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n335), .A2(new_n291), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT89), .B1(new_n356), .B2(new_n244), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n352), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT7), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n347), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n345), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n343), .B(new_n344), .C1(new_n362), .C2(new_n347), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n366), .B2(new_n340), .ZN(new_n367));
  OAI21_X1  g181(.A(G210), .B1(G237), .B2(G902), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n351), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n368), .B(KEYINPUT90), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n351), .B2(new_n367), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G214), .B1(G237), .B2(G902), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT92), .ZN(new_n377));
  NOR2_X1   g191(.A1(G475), .A2(G902), .ZN(new_n378));
  INV_X1    g192(.A(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G125), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(KEYINPUT16), .ZN(new_n381));
  INV_X1    g195(.A(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G140), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n383), .A3(KEYINPUT16), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT74), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n381), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n380), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n220), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n387), .ZN(new_n389));
  XNOR2_X1  g203(.A(G125), .B(G140), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT74), .B1(new_n390), .B2(KEYINPUT16), .ZN(new_n391));
  OAI211_X1 g205(.A(G146), .B(new_n389), .C1(new_n391), .C2(new_n381), .ZN(new_n392));
  NOR2_X1   g206(.A1(G237), .A2(G953), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n393), .A2(G143), .A3(G214), .ZN(new_n394));
  AOI21_X1  g208(.A(G143), .B1(new_n393), .B2(G214), .ZN(new_n395));
  OAI21_X1  g209(.A(G131), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT17), .ZN(new_n397));
  INV_X1    g211(.A(G237), .ZN(new_n398));
  INV_X1    g212(.A(G953), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(G214), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n225), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n393), .A2(G143), .A3(G214), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n205), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n396), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(KEYINPUT17), .B(G131), .C1(new_n394), .C2(new_n395), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n388), .A2(new_n392), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(G113), .B(G122), .Z(new_n407));
  XOR2_X1   g221(.A(KEYINPUT91), .B(G104), .Z(new_n408));
  XOR2_X1   g222(.A(new_n407), .B(new_n408), .Z(new_n409));
  AND3_X1   g223(.A1(new_n237), .A2(new_n390), .A3(KEYINPUT77), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT77), .B1(new_n237), .B2(new_n390), .ZN(new_n411));
  OAI22_X1  g225(.A1(new_n410), .A2(new_n411), .B1(new_n220), .B2(new_n390), .ZN(new_n412));
  NAND2_X1  g226(.A1(KEYINPUT18), .A2(G131), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n401), .A2(new_n402), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT18), .B(G131), .C1(new_n394), .C2(new_n395), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n406), .A2(new_n409), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n396), .A2(new_n403), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n380), .A2(new_n383), .A3(KEYINPUT19), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT19), .B1(new_n380), .B2(new_n383), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n237), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n392), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n409), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n378), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT20), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n418), .A2(new_n421), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n386), .A2(new_n220), .A3(new_n387), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n390), .A2(new_n220), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n237), .A2(new_n390), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT77), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n237), .A2(new_n390), .A3(KEYINPUT77), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n415), .A2(new_n414), .ZN(new_n434));
  OAI22_X1  g248(.A1(new_n426), .A2(new_n427), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n409), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n406), .A2(new_n416), .A3(new_n409), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n378), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n425), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n409), .B1(new_n406), .B2(new_n416), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n191), .B1(new_n417), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G475), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n377), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n440), .B1(new_n439), .B2(new_n378), .ZN(new_n447));
  INV_X1    g261(.A(new_n378), .ZN(new_n448));
  AOI211_X1 g262(.A(KEYINPUT20), .B(new_n448), .C1(new_n437), .C2(new_n438), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n445), .B(new_n377), .C1(new_n447), .C2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G478), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(KEYINPUT15), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n225), .A2(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n227), .A2(G143), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G134), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n456), .A3(new_n198), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G122), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G116), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n330), .A2(G122), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n463), .A3(new_n208), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n330), .A2(KEYINPUT14), .A3(G122), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n463), .ZN(new_n466));
  OAI211_X1 g280(.A(G107), .B(new_n465), .C1(new_n466), .C2(KEYINPUT14), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(G107), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n469), .A2(new_n464), .A3(KEYINPUT93), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT93), .B1(new_n469), .B2(new_n464), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT13), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n456), .B1(new_n455), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n455), .A2(new_n473), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n455), .A2(KEYINPUT94), .A3(new_n473), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n459), .B1(new_n479), .B2(new_n198), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n468), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G217), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n187), .A2(new_n482), .A3(G953), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n468), .B(new_n483), .C1(new_n472), .C2(new_n480), .ZN(new_n486));
  AOI21_X1  g300(.A(G902), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT95), .B1(new_n487), .B2(KEYINPUT96), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT95), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n489), .B(G902), .C1(new_n485), .C2(new_n486), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n454), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n485), .A2(new_n486), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT96), .A3(new_n191), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n489), .ZN(new_n494));
  INV_X1    g308(.A(new_n454), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT21), .B(G898), .ZN(new_n498));
  NAND2_X1  g312(.A1(G234), .A2(G237), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n498), .A2(G902), .A3(G953), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n399), .A2(G952), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(G234), .B2(G237), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n504), .B(KEYINPUT97), .Z(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n452), .A2(new_n497), .A3(new_n506), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n313), .A2(new_n376), .A3(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n509));
  NAND2_X1  g323(.A1(new_n393), .A2(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G101), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n355), .A2(new_n323), .B1(new_n318), .B2(new_n321), .ZN(new_n515));
  INV_X1    g329(.A(new_n202), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n198), .A2(G137), .ZN(new_n517));
  OAI21_X1  g331(.A(G131), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n518), .A2(new_n206), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n249), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n238), .A2(new_n262), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n207), .A2(new_n521), .A3(new_n260), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT30), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n515), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n520), .A2(new_n522), .A3(new_n515), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n514), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n515), .B1(new_n520), .B2(new_n522), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT28), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n534), .A3(new_n513), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n530), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT69), .ZN(new_n538));
  INV_X1    g352(.A(new_n531), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n528), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT70), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT28), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n532), .A2(KEYINPUT70), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n534), .B(KEYINPUT71), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n514), .A2(new_n536), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n530), .A2(new_n535), .A3(new_n548), .A4(new_n536), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n538), .A2(new_n191), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G472), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n532), .A2(new_n534), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n514), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n527), .A2(new_n529), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT31), .B1(new_n554), .B2(new_n513), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  NOR4_X1   g370(.A1(new_n527), .A2(new_n556), .A3(new_n529), .A4(new_n514), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(G472), .A2(G902), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT68), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n558), .A2(KEYINPUT32), .A3(new_n561), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n551), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n482), .B1(G234), .B2(new_n191), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n388), .A2(new_n392), .ZN(new_n568));
  INV_X1    g382(.A(G119), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G128), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n227), .A2(KEYINPUT23), .A3(G119), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n569), .A2(G128), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(KEYINPUT23), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G110), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n227), .A2(G119), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n570), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT72), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n570), .A3(KEYINPUT72), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT24), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G110), .ZN(new_n582));
  INV_X1    g396(.A(G110), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT24), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT73), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(KEYINPUT24), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n581), .A2(G110), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT73), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n568), .B(new_n574), .C1(new_n580), .C2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT78), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT76), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n573), .A2(G110), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT72), .B1(new_n575), .B2(new_n570), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n575), .A2(new_n570), .A3(KEYINPUT72), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n588), .B1(new_n586), .B2(new_n587), .ZN(new_n599));
  OAI22_X1  g413(.A1(new_n596), .A2(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT75), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT75), .B1(new_n580), .B2(new_n590), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n593), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n601), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n580), .A2(new_n590), .A3(KEYINPUT75), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n605), .A2(KEYINPUT76), .A3(new_n595), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n431), .A2(new_n432), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n392), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n592), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  AOI211_X1 g426(.A(KEYINPUT78), .B(new_n610), .C1(new_n604), .C2(new_n607), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n591), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n399), .A2(G221), .A3(G234), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT79), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT22), .B(G137), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n591), .B(new_n618), .C1(new_n612), .C2(new_n613), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT25), .B1(new_n622), .B2(new_n191), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT25), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n624), .B(G902), .C1(new_n620), .C2(new_n621), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n567), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n567), .A2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n566), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n508), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G101), .ZN(G3));
  NAND2_X1  g445(.A1(new_n558), .A2(new_n191), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n632), .A2(G472), .B1(new_n561), .B2(new_n558), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n626), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n368), .B1(new_n351), .B2(new_n367), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n374), .B(new_n505), .C1(new_n369), .C2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n453), .A2(G902), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n492), .A2(new_n638), .A3(KEYINPUT33), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT33), .B1(new_n492), .B2(new_n638), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n641), .B1(G478), .B2(new_n487), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n452), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n634), .A2(new_n313), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT99), .Z(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND2_X1  g462(.A1(new_n442), .A2(new_n445), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n497), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n636), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n634), .A2(new_n313), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT100), .Z(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT35), .B(G107), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  INV_X1    g470(.A(new_n633), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n618), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n614), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n627), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n657), .B1(new_n626), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n508), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  NAND2_X1  g478(.A1(new_n626), .A2(new_n660), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n374), .B1(new_n369), .B2(new_n635), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n499), .A2(new_n667), .A3(G902), .A4(G953), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n503), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n497), .A2(new_n650), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  AND4_X1   g485(.A1(new_n566), .A2(new_n665), .A3(new_n671), .A4(new_n313), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n227), .ZN(G30));
  INV_X1    g487(.A(new_n665), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n540), .A2(new_n514), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n554), .A2(new_n513), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n191), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G472), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n564), .A2(new_n565), .A3(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n446), .A2(new_n451), .ZN(new_n682));
  INV_X1    g496(.A(new_n497), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n374), .A2(new_n674), .A3(new_n681), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n669), .B(KEYINPUT39), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n313), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n373), .B(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n685), .A2(new_n688), .A3(new_n689), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT103), .B(G143), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G45));
  AOI22_X1  g508(.A1(G472), .A2(new_n550), .B1(new_n562), .B2(new_n563), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n565), .A2(new_n695), .B1(new_n626), .B2(new_n660), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n452), .A2(new_n642), .A3(new_n669), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n697), .B1(new_n666), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n666), .ZN(new_n700));
  INV_X1    g514(.A(new_n698), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(KEYINPUT104), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n696), .A2(new_n313), .A3(new_n699), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  INV_X1    g518(.A(new_n628), .ZN(new_n705));
  INV_X1    g519(.A(new_n607), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n578), .A2(new_n579), .B1(new_n585), .B2(new_n589), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n594), .B1(new_n707), .B2(KEYINPUT75), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT76), .B1(new_n708), .B2(new_n605), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n611), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT78), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n608), .A2(new_n592), .A3(new_n611), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n618), .B1(new_n713), .B2(new_n591), .ZN(new_n714));
  INV_X1    g528(.A(new_n621), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n191), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n624), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n622), .A2(KEYINPUT25), .A3(new_n191), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n705), .B1(new_n719), .B2(new_n567), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n285), .B1(new_n284), .B2(new_n207), .ZN(new_n721));
  AOI211_X1 g535(.A(KEYINPUT87), .B(new_n288), .C1(new_n279), .C2(new_n283), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n289), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n196), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n306), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(G469), .B1(new_n725), .B2(G902), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n726), .A2(new_n188), .A3(new_n307), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n720), .A2(new_n727), .A3(new_n644), .A4(new_n566), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  NAND4_X1  g544(.A1(new_n720), .A2(new_n727), .A3(new_n652), .A4(new_n566), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  NAND3_X1  g546(.A1(new_n665), .A2(new_n566), .A3(new_n683), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n682), .A2(new_n505), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n727), .A2(new_n736), .A3(new_n700), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n726), .A2(new_n307), .A3(new_n188), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT105), .B1(new_n738), .B2(new_n666), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  INV_X1    g556(.A(KEYINPUT71), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n534), .B(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n543), .B2(new_n542), .ZN(new_n745));
  OAI22_X1  g559(.A1(new_n745), .A2(new_n513), .B1(new_n555), .B2(new_n557), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n632), .A2(G472), .B1(new_n746), .B2(new_n561), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n626), .A2(new_n628), .A3(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n666), .A2(new_n683), .A3(new_n682), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n505), .A3(new_n727), .A4(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n626), .A2(new_n747), .A3(new_n628), .A4(new_n505), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n738), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(KEYINPUT106), .A3(new_n749), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G122), .ZN(G24));
  AND3_X1   g571(.A1(new_n665), .A2(new_n701), .A3(new_n747), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n736), .B1(new_n727), .B2(new_n700), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n738), .A2(KEYINPUT105), .A3(new_n666), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  NOR3_X1   g576(.A1(new_n369), .A2(new_n372), .A3(new_n375), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n313), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n698), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n565), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n558), .A2(KEYINPUT107), .A3(KEYINPUT32), .A4(new_n561), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n551), .A3(new_n564), .A4(new_n769), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n720), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n766), .B1(new_n720), .B2(new_n770), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n765), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT42), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n720), .A2(new_n566), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n698), .A2(KEYINPUT42), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n775), .A2(new_n764), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n205), .ZN(G33));
  NOR3_X1   g595(.A1(new_n775), .A2(new_n764), .A3(new_n670), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n198), .ZN(G36));
  OR2_X1    g597(.A1(new_n311), .A2(KEYINPUT45), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n311), .A2(KEYINPUT45), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(G469), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n190), .B2(new_n191), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n307), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n189), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n642), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n452), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT43), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n657), .A3(new_n665), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT44), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n373), .A2(new_n374), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n796), .B2(new_n797), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n792), .A2(new_n686), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  XNOR2_X1  g616(.A(new_n792), .B(KEYINPUT47), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n720), .A2(new_n566), .A3(new_n799), .A4(new_n698), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  NAND3_X1  g622(.A1(new_n720), .A2(new_n188), .A3(new_n374), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT110), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n691), .A2(new_n452), .A3(new_n793), .A4(new_n681), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n726), .A2(new_n307), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT49), .Z(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n502), .A2(new_n795), .A3(new_n727), .A4(new_n763), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n665), .A3(new_n747), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT113), .Z(new_n817));
  NAND2_X1  g631(.A1(new_n720), .A2(new_n502), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n818), .A2(new_n681), .A3(new_n738), .A4(new_n799), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n682), .A3(new_n793), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n812), .A2(new_n188), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n803), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n795), .A2(new_n502), .A3(new_n748), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n799), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n824), .A2(new_n374), .A3(new_n691), .A4(new_n738), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT50), .Z(new_n828));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n826), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n771), .A2(new_n772), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n815), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT48), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n824), .B1(new_n737), .B2(new_n739), .ZN(new_n838));
  INV_X1    g652(.A(new_n643), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n501), .B(new_n838), .C1(new_n839), .C2(new_n819), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n828), .A2(new_n833), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n826), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  INV_X1    g658(.A(new_n672), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n626), .A2(new_n660), .A3(new_n669), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n313), .A3(new_n681), .A4(new_n749), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n761), .A2(new_n845), .A3(new_n703), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n672), .B1(new_n740), .B2(new_n758), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(KEYINPUT52), .A3(new_n703), .A4(new_n847), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT106), .B1(new_n754), .B2(new_n749), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n700), .A2(new_n684), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n753), .A2(new_n855), .A3(new_n738), .A4(new_n751), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n741), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n508), .B1(new_n629), .B2(new_n661), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n374), .B(new_n505), .C1(new_n369), .C2(new_n372), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n497), .B1(new_n446), .B2(new_n451), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT111), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n860), .A2(new_n861), .B1(new_n452), .B2(new_n642), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n682), .A2(KEYINPUT111), .A3(new_n497), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n634), .A2(new_n864), .A3(new_n313), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n858), .A2(new_n728), .A3(new_n731), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n857), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n782), .ZN(new_n868));
  INV_X1    g682(.A(new_n764), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n650), .A2(new_n669), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n733), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n871), .B2(new_n758), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n774), .A2(new_n779), .A3(new_n868), .A4(new_n872), .ZN(new_n873));
  AND4_X1   g687(.A1(KEYINPUT53), .A2(new_n853), .A3(new_n867), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n774), .A2(new_n779), .A3(new_n868), .A4(new_n872), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n865), .A2(new_n728), .A3(new_n731), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n756), .A2(new_n741), .A3(new_n858), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT53), .B1(new_n878), .B2(new_n853), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n844), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n778), .B(new_n782), .C1(new_n773), .C2(KEYINPUT42), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n867), .A2(new_n882), .A3(new_n872), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n850), .A2(new_n852), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n878), .A2(KEYINPUT53), .A3(new_n853), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(KEYINPUT54), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n834), .A2(new_n843), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(G952), .A2(G953), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n814), .B1(new_n889), .B2(new_n890), .ZN(G75));
  NOR2_X1   g705(.A1(new_n399), .A2(G952), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT114), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n341), .A2(new_n350), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n348), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n191), .B1(new_n885), .B2(new_n886), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(G210), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n898), .A2(new_n370), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n897), .A2(new_n900), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n894), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(G51));
  XNOR2_X1  g718(.A(new_n725), .B(KEYINPUT116), .ZN(new_n905));
  XOR2_X1   g719(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n308), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n888), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n786), .B(KEYINPUT117), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n898), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n892), .B1(new_n908), .B2(new_n910), .ZN(G54));
  NAND2_X1  g725(.A1(KEYINPUT58), .A2(G475), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT118), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n898), .A2(new_n439), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n439), .B1(new_n898), .B2(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n892), .ZN(G60));
  OR2_X1    g730(.A1(new_n639), .A2(new_n640), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n453), .A2(new_n191), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n919), .B(new_n920), .Z(new_n921));
  NOR2_X1   g735(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n880), .A2(new_n887), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT120), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n880), .A2(new_n887), .A3(new_n925), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n921), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n880), .A2(new_n887), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n894), .B1(new_n929), .B2(new_n918), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n927), .A2(KEYINPUT121), .A3(new_n930), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(G63));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n936));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT60), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n885), .B2(new_n886), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n894), .B1(new_n939), .B2(new_n659), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n940), .B2(KEYINPUT122), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n622), .B2(new_n939), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n941), .B(new_n942), .Z(G66));
  NAND2_X1  g757(.A1(new_n877), .A2(new_n399), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT123), .Z(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n498), .B2(new_n346), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n895), .B1(G898), .B2(new_n399), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G69));
  OAI21_X1  g763(.A(G953), .B1(new_n194), .B2(new_n667), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT125), .Z(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n524), .A2(new_n526), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n419), .A2(new_n420), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(G900), .B2(G953), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n851), .A2(new_n703), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n792), .A2(new_n686), .A3(new_n749), .A4(new_n835), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n882), .A2(new_n801), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n807), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n956), .B1(new_n960), .B2(G953), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n955), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n957), .A2(new_n692), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT62), .Z(new_n965));
  AOI21_X1  g779(.A(new_n799), .B1(new_n863), .B2(new_n862), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n629), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n801), .B1(new_n687), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT124), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n807), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n963), .B1(new_n970), .B2(new_n399), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n952), .B1(new_n962), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n970), .A2(new_n399), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n961), .B(new_n951), .C1(new_n973), .C2(new_n963), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(G72));
  XOR2_X1   g789(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n976));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n970), .B2(new_n877), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n979), .B(new_n513), .C1(new_n529), .C2(new_n527), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n677), .A2(new_n530), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n978), .B(new_n981), .C1(new_n874), .C2(new_n879), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n978), .B1(new_n960), .B2(new_n877), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n554), .A2(new_n514), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT127), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n892), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n980), .A2(new_n982), .A3(new_n986), .ZN(G57));
endmodule


