//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(new_n456), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(G101), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT70), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n473), .A2(new_n470), .A3(G101), .A4(G2104), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n469), .A2(G137), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n476), .B1(new_n467), .B2(new_n468), .ZN(new_n477));
  AND2_X1   g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n469), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n470), .B2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n467), .A2(new_n468), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT71), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n485), .B1(new_n488), .B2(G124), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(KEYINPUT73), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n491), .B(G138), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(G102), .A2(G2104), .ZN(new_n495));
  AOI21_X1  g070(.A(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n469), .B2(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(G126), .B1(new_n493), .B2(new_n492), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G114), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n500), .A2(new_n502), .A3(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n470), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n496), .A2(new_n497), .A3(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT5), .B1(new_n506), .B2(KEYINPUT74), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(G543), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n511), .A2(G62), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n517), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(new_n516), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT75), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT75), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n523), .B(new_n527), .C1(new_n524), .C2(new_n516), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n511), .A2(new_n512), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n526), .A2(new_n528), .A3(new_n530), .A4(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n513), .A2(new_n535), .B1(new_n536), .B2(new_n516), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n518), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  XOR2_X1   g118(.A(KEYINPUT77), .B(G81), .Z(new_n544));
  NAND2_X1  g119(.A1(new_n531), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n546), .B2(new_n516), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n511), .A2(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n518), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT78), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT79), .Z(G188));
  INV_X1    g133(.A(new_n516), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n559), .B(G53), .C1(KEYINPUT80), .C2(new_n560), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT80), .B(KEYINPUT9), .Z(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n516), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n507), .A2(new_n510), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n561), .A2(new_n564), .B1(G651), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n511), .A2(G91), .A3(new_n512), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT81), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G299));
  OR2_X1    g148(.A1(new_n517), .A2(new_n521), .ZN(G303));
  NAND4_X1  g149(.A1(new_n512), .A2(G87), .A3(new_n507), .A4(new_n510), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n512), .A2(G49), .A3(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(G74), .B1(new_n507), .B2(new_n510), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n518), .C2(new_n577), .ZN(G288));
  NAND4_X1  g153(.A1(new_n512), .A2(G86), .A3(new_n507), .A4(new_n510), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n507), .A2(new_n510), .A3(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n518), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n566), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n518), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n591), .B2(new_n590), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n531), .A2(G85), .B1(G47), .B2(new_n559), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G290));
  NAND3_X1  g170(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n513), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n596), .A2(new_n599), .B1(G54), .B2(new_n559), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n566), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT83), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n518), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(new_n603), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G171), .B2(new_n608), .ZN(G284));
  OAI21_X1  g185(.A(new_n609), .B1(G171), .B2(new_n608), .ZN(G321));
  NAND2_X1  g186(.A1(G299), .A2(new_n608), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G168), .B2(new_n608), .ZN(G280));
  XOR2_X1   g188(.A(G280), .B(KEYINPUT84), .Z(G297));
  INV_X1    g189(.A(new_n607), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g196(.A(G2096), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n469), .A2(G135), .ZN(new_n623));
  NOR2_X1   g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(new_n470), .B2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(new_n488), .B2(G123), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n622), .A2(new_n627), .B1(new_n631), .B2(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(G2100), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n632), .B(new_n633), .C1(new_n622), .C2(new_n627), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT86), .Z(G401));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT17), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(new_n652), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT87), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n657), .A2(new_n654), .A3(new_n652), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n658), .A2(new_n654), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n663), .B1(new_n653), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n622), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(G227));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT88), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n670), .B2(new_n673), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT90), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n675), .B(new_n677), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n670), .A2(new_n673), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n679), .A2(new_n672), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT91), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  MUX2_X1   g268(.A(G6), .B(G305), .S(G16), .Z(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT93), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT32), .B(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G23), .ZN(new_n700));
  INV_X1    g275(.A(G288), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n699), .A2(G22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT94), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n699), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT95), .Z(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n704), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n708), .A2(new_n709), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n698), .A2(new_n710), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n710), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT34), .B1(new_n714), .B2(new_n697), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G25), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(new_n470), .B2(G107), .ZN(new_n718));
  INV_X1    g293(.A(G95), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n470), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT92), .Z(new_n721));
  INV_X1    g296(.A(G131), .ZN(new_n722));
  INV_X1    g297(.A(new_n469), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n488), .A2(G119), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n717), .B1(new_n726), .B2(new_n716), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n727), .B(new_n729), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n699), .A2(G24), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G290), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1986), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n730), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n713), .A2(new_n715), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(KEYINPUT96), .A2(KEYINPUT36), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n713), .A2(new_n738), .A3(new_n715), .A4(new_n736), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n615), .A2(new_n699), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G4), .B2(new_n699), .ZN(new_n744));
  INV_X1    g319(.A(G1348), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n716), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n716), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT29), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n746), .B(new_n747), .C1(G2090), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(G2090), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT101), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n699), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n551), .B2(new_n699), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1341), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n699), .A2(G20), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT102), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT23), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G299), .B2(G16), .ZN(new_n760));
  INV_X1    g335(.A(G1956), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n716), .A2(G26), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n469), .A2(G140), .ZN(new_n765));
  NOR2_X1   g340(.A1(G104), .A2(G2105), .ZN(new_n766));
  OAI21_X1  g341(.A(G2104), .B1(new_n470), .B2(G116), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n488), .B2(G128), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n764), .B1(new_n769), .B2(new_n716), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n756), .A2(new_n762), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n751), .A2(new_n753), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n699), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n699), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1961), .ZN(new_n776));
  INV_X1    g351(.A(G32), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n488), .A2(G129), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n469), .A2(G141), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT97), .B(KEYINPUT26), .Z(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n470), .A2(G105), .A3(G2104), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n779), .A2(new_n780), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(G29), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT98), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT27), .B(G1996), .Z(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n791), .B1(new_n788), .B2(new_n789), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n776), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n716), .A2(G27), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G164), .B2(new_n716), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT99), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2078), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n699), .A2(G21), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G168), .B2(new_n699), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1966), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n716), .A2(G33), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT25), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n470), .ZN(new_n807));
  AOI211_X1 g382(.A(new_n805), .B(new_n807), .C1(G139), .C2(new_n469), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n803), .B1(new_n808), .B2(new_n716), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(G2072), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(G2072), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT30), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n812), .A2(G28), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n716), .B1(new_n812), .B2(G28), .ZN(new_n814));
  AND2_X1   g389(.A1(KEYINPUT31), .A2(G11), .ZN(new_n815));
  NOR2_X1   g390(.A1(KEYINPUT31), .A2(G11), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n813), .A2(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n627), .B2(G29), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n810), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n716), .B1(KEYINPUT24), .B2(G34), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(KEYINPUT24), .B2(G34), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n480), .B2(G29), .ZN(new_n822));
  INV_X1    g397(.A(G2084), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n802), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n795), .A2(new_n799), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT100), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n795), .A2(KEYINPUT100), .A3(new_n799), .A4(new_n825), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n773), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n742), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(G311));
  NAND3_X1  g407(.A1(new_n742), .A2(new_n830), .A3(KEYINPUT103), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT103), .B1(new_n742), .B2(new_n830), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(G150));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  INV_X1    g412(.A(G55), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n513), .A2(new_n837), .B1(new_n838), .B2(new_n516), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n511), .A2(G67), .ZN(new_n840));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n518), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n551), .A2(KEYINPUT104), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(KEYINPUT104), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n548), .A2(new_n549), .ZN(new_n846));
  OAI221_X1 g421(.A(new_n545), .B1(new_n546), .B2(new_n516), .C1(new_n846), .C2(new_n518), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT104), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n839), .B2(new_n842), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT38), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n615), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  INV_X1    g430(.A(G860), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n843), .A2(new_n856), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT105), .B(KEYINPUT37), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(G145));
  INV_X1    g437(.A(KEYINPUT73), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n863), .A2(KEYINPUT4), .A3(G138), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n467), .B2(new_n468), .ZN(new_n865));
  INV_X1    g440(.A(new_n495), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n470), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(new_n499), .B2(G114), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G126), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(new_n467), .B2(new_n468), .ZN(new_n872));
  OAI21_X1  g447(.A(G2105), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI211_X1 g448(.A(G138), .B(new_n470), .C1(new_n493), .C2(new_n492), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(KEYINPUT73), .B2(new_n490), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n867), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n769), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n808), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n726), .B(new_n629), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n469), .A2(G142), .ZN(new_n881));
  NOR2_X1   g456(.A1(G106), .A2(G2105), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(new_n470), .B2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n488), .B2(G130), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n785), .B(new_n885), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n880), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G162), .B(new_n480), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n627), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n887), .A2(new_n890), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g470(.A(new_n851), .B(new_n618), .Z(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n615), .A2(G299), .ZN(new_n898));
  INV_X1    g473(.A(G299), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n607), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(KEYINPUT106), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n615), .A2(new_n902), .A3(G299), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n897), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n898), .A2(KEYINPUT107), .A3(new_n900), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n615), .A2(KEYINPUT107), .A3(G299), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n905), .A2(new_n906), .A3(new_n897), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n896), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(new_n903), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n908), .B1(new_n896), .B2(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(G305), .ZN(new_n912));
  XNOR2_X1  g487(.A(G290), .B(new_n701), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(KEYINPUT108), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(KEYINPUT108), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n911), .B2(new_n917), .ZN(new_n919));
  OAI21_X1  g494(.A(G868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(G868), .B2(new_n843), .ZN(G295));
  OAI21_X1  g496(.A(new_n920), .B1(G868), .B2(new_n843), .ZN(G331));
  NAND2_X1  g497(.A1(new_n851), .A2(G171), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n844), .A2(new_n850), .A3(G301), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(G286), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(G168), .A3(new_n924), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n926), .B(new_n927), .C1(new_n907), .C2(new_n904), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n923), .A2(G168), .A3(new_n924), .ZN(new_n929));
  AOI21_X1  g504(.A(G168), .B1(new_n923), .B2(new_n924), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n903), .B(new_n901), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n931), .A3(new_n916), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n892), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n916), .B1(new_n928), .B2(new_n931), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(KEYINPUT109), .B(KEYINPUT43), .C1(new_n933), .C2(new_n934), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n929), .A2(new_n930), .A3(new_n897), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n905), .A2(new_n906), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n916), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n901), .A2(new_n903), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n941), .B1(new_n942), .B2(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n892), .A4(new_n932), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n938), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND4_X1   g523(.A1(KEYINPUT43), .A2(new_n943), .A3(new_n892), .A4(new_n932), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n933), .A2(new_n934), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT44), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(G397));
  XOR2_X1   g528(.A(KEYINPUT114), .B(G8), .Z(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(KEYINPUT112), .B(G1971), .Z(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n475), .A2(new_n479), .A3(G40), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n876), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n961));
  AOI21_X1  g536(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n958), .ZN(new_n965));
  NOR2_X1   g540(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n965), .B1(G164), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n876), .B2(new_n959), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n968), .A2(new_n970), .A3(G2090), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n955), .B1(new_n964), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G8), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n974));
  OR3_X1    g549(.A1(G166), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(G166), .B2(new_n973), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n972), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n977), .B(G8), .C1(new_n971), .C2(new_n964), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n965), .A2(new_n959), .A3(new_n876), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n955), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n983));
  INV_X1    g558(.A(G1976), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(G288), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n575), .A2(new_n576), .ZN(new_n986));
  OAI21_X1  g561(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(KEYINPUT115), .A3(G1976), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1981), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n582), .A2(new_n586), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(G1981), .B1(new_n581), .B2(new_n585), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(KEYINPUT49), .A3(new_n993), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n955), .A3(new_n981), .A4(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n985), .A2(new_n988), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(G288), .B2(new_n984), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(new_n955), .A3(new_n981), .A4(new_n1000), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n990), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n979), .A2(new_n980), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G2078), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n962), .A2(new_n1004), .A3(new_n963), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n958), .B1(new_n876), .B2(new_n966), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1961), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(G164), .B2(G1384), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n961), .A2(G1384), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n958), .B1(new_n876), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1006), .A2(G2078), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(G171), .B1(new_n1008), .B2(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1003), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1966), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n876), .A2(new_n1016), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n965), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT45), .B1(new_n876), .B2(new_n959), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1009), .A2(new_n823), .A3(new_n1010), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G286), .A2(new_n955), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1029), .A2(G8), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(new_n1030), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n954), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(KEYINPUT122), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n968), .A2(new_n970), .A3(G2084), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1966), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n955), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1036), .B1(new_n1045), .B2(KEYINPUT123), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT123), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1039), .A2(new_n1047), .A3(new_n1044), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1033), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1022), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT122), .B(new_n955), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1037), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1038), .A2(KEYINPUT122), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT123), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1036), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1048), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1032), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT126), .B1(new_n1059), .B2(KEYINPUT62), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT126), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1061), .B(new_n1050), .C1(new_n1058), .C2(new_n1032), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1051), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT127), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT127), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1051), .B(new_n1065), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n954), .B(G286), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n979), .A2(new_n980), .A3(new_n1002), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT63), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(KEYINPUT117), .A3(new_n1069), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n990), .A2(new_n998), .A3(new_n1001), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT116), .ZN(new_n1075));
  OAI21_X1  g650(.A(G8), .B1(new_n964), .B2(new_n971), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n978), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1042), .A2(new_n1069), .A3(G286), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1075), .A2(new_n980), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1072), .A2(new_n1073), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n998), .A2(new_n984), .A3(new_n701), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n982), .B1(new_n1081), .B2(new_n992), .ZN(new_n1082));
  INV_X1    g657(.A(new_n980), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1075), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1003), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1021), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n960), .A2(new_n961), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1089), .A2(new_n965), .A3(new_n963), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1018), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT124), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n1093));
  AOI211_X1 g668(.A(new_n1093), .B(G1961), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1091), .B(new_n1007), .C1(new_n1092), .C2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT125), .B1(new_n1095), .B2(G171), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1091), .A2(new_n1007), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT125), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .A4(G301), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1088), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1098), .A3(G171), .ZN(new_n1102));
  OAI21_X1  g677(.A(G301), .B1(new_n1008), .B2(new_n1020), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1102), .A2(KEYINPUT54), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1086), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(new_n1049), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n561), .A2(new_n564), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT57), .B1(new_n1107), .B2(KEYINPUT118), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G299), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n561), .B2(new_n564), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n569), .B(new_n572), .C1(new_n1111), .C2(KEYINPUT57), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1011), .A2(new_n761), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT119), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n962), .A2(new_n963), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1011), .A2(new_n745), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(G2067), .B2(new_n981), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1120), .A2(new_n615), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1113), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT61), .B1(new_n1122), .B2(KEYINPUT120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n1118), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1124), .A2(new_n1128), .A3(KEYINPUT121), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT121), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G1996), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1090), .A2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n981), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT59), .B1(new_n1136), .B2(new_n551), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1120), .A2(KEYINPUT60), .A3(new_n607), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1120), .A2(new_n615), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT60), .B1(new_n1121), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1126), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1136), .A2(KEYINPUT59), .A3(new_n551), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1123), .B1(new_n1131), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1085), .B1(new_n1106), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1064), .A2(new_n1066), .A3(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1089), .A2(new_n958), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n726), .A2(new_n728), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n724), .A2(new_n725), .A3(new_n729), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1152), .A2(KEYINPUT111), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n785), .B(G1996), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n769), .B(G2067), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1152), .A2(KEYINPUT111), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1153), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(G290), .A2(G1986), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n593), .A2(new_n733), .A3(new_n594), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1148), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1147), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1148), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1157), .A2(new_n1150), .ZN(new_n1166));
  INV_X1    g741(.A(G2067), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n769), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1165), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1148), .B1(new_n1156), .B2(new_n785), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1148), .A2(KEYINPUT46), .A3(new_n1132), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT46), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1165), .B2(G1996), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT47), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n1159), .A2(new_n1148), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1165), .A2(new_n1161), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1177), .B(KEYINPUT48), .Z(new_n1178));
  AOI211_X1 g753(.A(new_n1169), .B(new_n1175), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1164), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g755(.A1(G227), .A2(G401), .A3(new_n463), .ZN(new_n1182));
  AND2_X1   g756(.A1(new_n692), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g757(.A1(new_n946), .A2(new_n1183), .A3(new_n894), .ZN(G225));
  INV_X1    g758(.A(G225), .ZN(G308));
endmodule


