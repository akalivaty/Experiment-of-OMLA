

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769;

  OR2_X1 U370 ( .A1(n502), .A2(KEYINPUT83), .ZN(n494) );
  XNOR2_X1 U371 ( .A(n635), .B(KEYINPUT111), .ZN(n764) );
  NAND2_X1 U372 ( .A1(n608), .A2(n607), .ZN(n606) );
  XNOR2_X1 U373 ( .A(n556), .B(n450), .ZN(n449) );
  INV_X1 U374 ( .A(n515), .ZN(n559) );
  XNOR2_X1 U375 ( .A(n523), .B(n522), .ZN(n557) );
  XNOR2_X2 U376 ( .A(G101), .B(G104), .ZN(n531) );
  XNOR2_X1 U377 ( .A(n449), .B(n557), .ZN(n749) );
  XNOR2_X2 U378 ( .A(n503), .B(KEYINPUT77), .ZN(n673) );
  INV_X1 U379 ( .A(n675), .ZN(n632) );
  XNOR2_X1 U380 ( .A(n552), .B(n553), .ZN(n622) );
  INV_X1 U381 ( .A(G146), .ZN(n443) );
  INV_X1 U382 ( .A(G953), .ZN(n748) );
  BUF_X1 U383 ( .A(n603), .Z(n459) );
  XNOR2_X1 U384 ( .A(n443), .B(G125), .ZN(n558) );
  NOR2_X2 U385 ( .A1(n426), .A2(KEYINPUT69), .ZN(n597) );
  NOR2_X1 U386 ( .A1(n701), .A2(n622), .ZN(n624) );
  XNOR2_X1 U387 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U388 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n515) );
  INV_X1 U389 ( .A(G122), .ZN(n451) );
  BUF_X1 U390 ( .A(n652), .Z(n756) );
  NAND2_X1 U391 ( .A1(n494), .A2(n495), .ZN(n652) );
  AND2_X1 U392 ( .A1(n500), .A2(n496), .ZN(n495) );
  AND2_X1 U393 ( .A1(n374), .A2(n373), .ZN(n382) );
  NOR2_X1 U394 ( .A1(n768), .A2(n668), .ZN(n465) );
  NAND2_X1 U395 ( .A1(n436), .A2(n349), .ZN(n635) );
  AND2_X1 U396 ( .A1(n397), .A2(n398), .ZN(n389) );
  XNOR2_X1 U397 ( .A(n629), .B(n419), .ZN(n767) );
  XNOR2_X1 U398 ( .A(n431), .B(n430), .ZN(n699) );
  XNOR2_X1 U399 ( .A(n433), .B(n362), .ZN(n482) );
  XNOR2_X1 U400 ( .A(n383), .B(n456), .ZN(n631) );
  NAND2_X1 U401 ( .A1(n636), .A2(n691), .ZN(n634) );
  OR2_X2 U402 ( .A1(n416), .A2(n417), .ZN(n636) );
  XNOR2_X1 U403 ( .A(n445), .B(n749), .ZN(n655) );
  XNOR2_X1 U404 ( .A(n571), .B(n572), .ZN(n755) );
  XNOR2_X1 U405 ( .A(n557), .B(n525), .ZN(n529) );
  AND2_X1 U406 ( .A1(n509), .A2(n508), .ZN(n507) );
  XNOR2_X1 U407 ( .A(n558), .B(n442), .ZN(n570) );
  XNOR2_X1 U408 ( .A(n451), .B(KEYINPUT16), .ZN(n450) );
  XNOR2_X1 U409 ( .A(n399), .B(G902), .ZN(n651) );
  XNOR2_X1 U410 ( .A(KEYINPUT3), .B(KEYINPUT71), .ZN(n521) );
  NOR2_X1 U411 ( .A1(n673), .A2(n696), .ZN(n422) );
  XNOR2_X2 U412 ( .A(n483), .B(n363), .ZN(n741) );
  NOR2_X1 U413 ( .A1(n643), .A2(n671), .ZN(n374) );
  OR2_X1 U414 ( .A1(n727), .A2(G902), .ZN(n427) );
  XNOR2_X1 U415 ( .A(n764), .B(KEYINPUT85), .ZN(n373) );
  NAND2_X1 U416 ( .A1(n376), .A2(n375), .ZN(n381) );
  AND2_X1 U417 ( .A1(n378), .A2(n377), .ZN(n376) );
  NOR2_X1 U418 ( .A1(n767), .A2(n379), .ZN(n371) );
  NAND2_X1 U419 ( .A1(n655), .A2(n348), .ZN(n415) );
  INV_X1 U420 ( .A(KEYINPUT38), .ZN(n458) );
  INV_X1 U421 ( .A(n608), .ZN(n605) );
  INV_X1 U422 ( .A(KEYINPUT28), .ZN(n504) );
  NAND2_X1 U423 ( .A1(n769), .A2(n379), .ZN(n378) );
  NAND2_X1 U424 ( .A1(n767), .A2(n379), .ZN(n377) );
  INV_X1 U425 ( .A(KEYINPUT48), .ZN(n470) );
  NAND2_X1 U426 ( .A1(n382), .A2(n381), .ZN(n380) );
  NAND2_X1 U427 ( .A1(n499), .A2(n498), .ZN(n497) );
  INV_X1 U428 ( .A(KEYINPUT83), .ZN(n498) );
  INV_X1 U429 ( .A(n682), .ZN(n499) );
  NAND2_X1 U430 ( .A1(n348), .A2(n651), .ZN(n418) );
  INV_X1 U431 ( .A(KEYINPUT0), .ZN(n485) );
  NAND2_X1 U432 ( .A1(n488), .A2(KEYINPUT0), .ZN(n487) );
  INV_X1 U433 ( .A(n518), .ZN(n488) );
  NAND2_X1 U434 ( .A1(n409), .A2(n356), .ZN(n408) );
  XNOR2_X1 U435 ( .A(n541), .B(n540), .ZN(n583) );
  XNOR2_X1 U436 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n540) );
  XOR2_X1 U437 ( .A(KEYINPUT92), .B(G110), .Z(n543) );
  XNOR2_X1 U438 ( .A(G119), .B(G137), .ZN(n542) );
  XNOR2_X1 U439 ( .A(n539), .B(n355), .ZN(n469) );
  XNOR2_X1 U440 ( .A(G128), .B(G140), .ZN(n538) );
  XNOR2_X1 U441 ( .A(KEYINPUT70), .B(KEYINPUT10), .ZN(n442) );
  INV_X1 U442 ( .A(G134), .ZN(n519) );
  XNOR2_X1 U443 ( .A(G116), .B(G122), .ZN(n581) );
  XOR2_X1 U444 ( .A(KEYINPUT9), .B(G107), .Z(n582) );
  XNOR2_X1 U445 ( .A(n755), .B(n580), .ZN(n731) );
  XNOR2_X1 U446 ( .A(n576), .B(n463), .ZN(n578) );
  XNOR2_X1 U447 ( .A(n447), .B(n446), .ZN(n445) );
  XNOR2_X1 U448 ( .A(n448), .B(n491), .ZN(n447) );
  XNOR2_X1 U449 ( .A(n452), .B(KEYINPUT39), .ZN(n650) );
  NAND2_X1 U450 ( .A1(n479), .A2(n482), .ZN(n452) );
  NOR2_X1 U451 ( .A1(n618), .A2(n480), .ZN(n479) );
  AND2_X1 U452 ( .A1(n396), .A2(n395), .ZN(n392) );
  INV_X1 U453 ( .A(n358), .ZN(n395) );
  INV_X1 U454 ( .A(KEYINPUT33), .ZN(n430) );
  NAND2_X1 U455 ( .A1(n705), .A2(n428), .ZN(n431) );
  NOR2_X1 U456 ( .A1(n631), .A2(n429), .ZN(n428) );
  XNOR2_X1 U457 ( .A(G478), .B(n588), .ZN(n607) );
  NAND2_X1 U458 ( .A1(n473), .A2(n476), .ZN(n472) );
  NAND2_X1 U459 ( .A1(n555), .A2(n475), .ZN(n474) );
  NAND2_X1 U460 ( .A1(n684), .A2(n651), .ZN(n405) );
  INV_X1 U461 ( .A(KEYINPUT46), .ZN(n379) );
  XNOR2_X1 U462 ( .A(n422), .B(n421), .ZN(n643) );
  INV_X1 U463 ( .A(KEYINPUT47), .ZN(n421) );
  NAND2_X1 U464 ( .A1(n514), .A2(n513), .ZN(n512) );
  NAND2_X1 U465 ( .A1(n515), .A2(G137), .ZN(n514) );
  NAND2_X1 U466 ( .A1(n559), .A2(n516), .ZN(n513) );
  XOR2_X1 U467 ( .A(G131), .B(G140), .Z(n572) );
  INV_X1 U468 ( .A(n622), .ZN(n702) );
  XOR2_X1 U469 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n527) );
  XNOR2_X1 U470 ( .A(G131), .B(G101), .ZN(n526) );
  AND2_X1 U471 ( .A1(n412), .A2(n411), .ZN(n410) );
  NOR2_X1 U472 ( .A1(n617), .A2(n406), .ZN(n411) );
  AND2_X1 U473 ( .A1(n497), .A2(n681), .ZN(n496) );
  XNOR2_X1 U474 ( .A(n577), .B(n464), .ZN(n463) );
  INV_X1 U475 ( .A(KEYINPUT98), .ZN(n464) );
  NOR2_X1 U476 ( .A1(G237), .A2(G953), .ZN(n524) );
  XNOR2_X1 U477 ( .A(n558), .B(n490), .ZN(n448) );
  XNOR2_X1 U478 ( .A(KEYINPUT76), .B(KEYINPUT18), .ZN(n490) );
  XNOR2_X1 U479 ( .A(n492), .B(KEYINPUT17), .ZN(n491) );
  NAND2_X1 U480 ( .A1(n748), .A2(G224), .ZN(n492) );
  OR2_X1 U481 ( .A1(G237), .A2(G902), .ZN(n561) );
  INV_X1 U482 ( .A(n459), .ZN(n397) );
  NAND2_X1 U483 ( .A1(n622), .A2(n400), .ZN(n429) );
  NAND2_X1 U484 ( .A1(n415), .A2(n418), .ZN(n417) );
  INV_X1 U485 ( .A(G902), .ZN(n475) );
  NAND2_X1 U486 ( .A1(n477), .A2(G902), .ZN(n476) );
  INV_X1 U487 ( .A(n429), .ZN(n706) );
  AND2_X1 U488 ( .A1(n489), .A2(n487), .ZN(n486) );
  XNOR2_X1 U489 ( .A(n457), .B(KEYINPUT104), .ZN(n456) );
  INV_X1 U490 ( .A(KEYINPUT6), .ZN(n457) );
  XOR2_X1 U491 ( .A(G116), .B(G113), .Z(n522) );
  XNOR2_X1 U492 ( .A(n521), .B(n520), .ZN(n523) );
  INV_X1 U493 ( .A(G119), .ZN(n520) );
  INV_X1 U494 ( .A(n423), .ZN(n532) );
  XNOR2_X1 U495 ( .A(G110), .B(G107), .ZN(n423) );
  NAND2_X1 U496 ( .A1(n387), .A2(n386), .ZN(n684) );
  XNOR2_X1 U497 ( .A(n434), .B(n350), .ZN(n608) );
  OR2_X1 U498 ( .A1(n731), .A2(G902), .ZN(n434) );
  NAND2_X1 U499 ( .A1(G953), .A2(G900), .ZN(n760) );
  XNOR2_X1 U500 ( .A(n570), .B(n469), .ZN(n547) );
  XNOR2_X1 U501 ( .A(n420), .B(n586), .ZN(n734) );
  XNOR2_X1 U502 ( .A(n587), .B(n351), .ZN(n420) );
  XOR2_X1 U503 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n585) );
  XNOR2_X1 U504 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U505 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n419) );
  INV_X1 U506 ( .A(KEYINPUT40), .ZN(n432) );
  AND2_X1 U507 ( .A1(n438), .A2(n437), .ZN(n436) );
  AND2_X1 U508 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U509 ( .A(n592), .B(KEYINPUT32), .ZN(n768) );
  AND2_X1 U510 ( .A1(n611), .A2(n353), .ZN(n592) );
  AND2_X1 U511 ( .A1(n595), .A2(n354), .ZN(n668) );
  XNOR2_X1 U512 ( .A(n606), .B(KEYINPUT102), .ZN(n675) );
  INV_X1 U513 ( .A(KEYINPUT122), .ZN(n461) );
  OR2_X1 U514 ( .A1(n694), .A2(n701), .ZN(n347) );
  XNOR2_X1 U515 ( .A(n636), .B(n458), .ZN(n692) );
  XOR2_X1 U516 ( .A(n560), .B(KEYINPUT90), .Z(n348) );
  AND2_X1 U517 ( .A1(n435), .A2(n705), .ZN(n349) );
  XOR2_X1 U518 ( .A(n569), .B(n568), .Z(n350) );
  XOR2_X1 U519 ( .A(n582), .B(n581), .Z(n351) );
  XOR2_X1 U520 ( .A(n556), .B(n535), .Z(n352) );
  INV_X1 U521 ( .A(n701), .ZN(n400) );
  INV_X1 U522 ( .A(G137), .ZN(n516) );
  NOR2_X1 U523 ( .A1(n612), .A2(n622), .ZN(n353) );
  NOR2_X1 U524 ( .A1(n621), .A2(n622), .ZN(n354) );
  XOR2_X1 U525 ( .A(KEYINPUT23), .B(KEYINPUT75), .Z(n355) );
  NAND2_X1 U526 ( .A1(n426), .A2(KEYINPUT69), .ZN(n356) );
  NAND2_X1 U527 ( .A1(n518), .A2(n485), .ZN(n357) );
  OR2_X1 U528 ( .A1(n605), .A2(n607), .ZN(n358) );
  OR2_X1 U529 ( .A1(n348), .A2(n651), .ZN(n359) );
  INV_X1 U530 ( .A(n623), .ZN(n481) );
  AND2_X1 U531 ( .A1(n441), .A2(n440), .ZN(n360) );
  XOR2_X1 U532 ( .A(KEYINPUT72), .B(KEYINPUT22), .Z(n361) );
  XNOR2_X1 U533 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n362) );
  INV_X1 U534 ( .A(KEYINPUT34), .ZN(n398) );
  INV_X1 U535 ( .A(KEYINPUT36), .ZN(n440) );
  XOR2_X1 U536 ( .A(KEYINPUT45), .B(KEYINPUT82), .Z(n363) );
  XOR2_X1 U537 ( .A(n729), .B(n728), .Z(n364) );
  XOR2_X1 U538 ( .A(n554), .B(KEYINPUT62), .Z(n365) );
  XOR2_X1 U539 ( .A(n731), .B(n517), .Z(n366) );
  INV_X1 U540 ( .A(n740), .ZN(n467) );
  XOR2_X1 U541 ( .A(n654), .B(KEYINPUT112), .Z(n367) );
  XOR2_X1 U542 ( .A(KEYINPUT60), .B(KEYINPUT68), .Z(n368) );
  XOR2_X1 U543 ( .A(KEYINPUT84), .B(KEYINPUT56), .Z(n369) );
  XOR2_X1 U544 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n370) );
  INV_X1 U545 ( .A(KEYINPUT2), .ZN(n424) );
  XNOR2_X1 U546 ( .A(n652), .B(KEYINPUT73), .ZN(n403) );
  NAND2_X1 U547 ( .A1(n372), .A2(n371), .ZN(n375) );
  INV_X1 U548 ( .A(n769), .ZN(n372) );
  XNOR2_X2 U549 ( .A(n380), .B(n470), .ZN(n502) );
  XNOR2_X2 U550 ( .A(n383), .B(KEYINPUT105), .ZN(n621) );
  NOR2_X1 U551 ( .A1(n601), .A2(n383), .ZN(n602) );
  NAND2_X1 U552 ( .A1(n710), .A2(n383), .ZN(n712) );
  NAND2_X1 U553 ( .A1(n600), .A2(n383), .ZN(n663) );
  OR2_X4 U554 ( .A1(n472), .A2(n471), .ZN(n383) );
  XNOR2_X2 U555 ( .A(n384), .B(n519), .ZN(n587) );
  XNOR2_X1 U556 ( .A(n384), .B(n559), .ZN(n446) );
  XNOR2_X2 U557 ( .A(n493), .B(G143), .ZN(n384) );
  XNOR2_X2 U558 ( .A(n385), .B(n432), .ZN(n769) );
  NAND2_X1 U559 ( .A1(n650), .A2(n632), .ZN(n385) );
  NAND2_X1 U560 ( .A1(n387), .A2(n404), .ZN(n388) );
  NOR2_X1 U561 ( .A1(n741), .A2(n424), .ZN(n386) );
  INV_X1 U562 ( .A(n756), .ZN(n387) );
  AND2_X1 U563 ( .A1(n388), .A2(n370), .ZN(n683) );
  NAND2_X1 U564 ( .A1(n390), .A2(n389), .ZN(n393) );
  INV_X1 U565 ( .A(n699), .ZN(n390) );
  NAND2_X1 U566 ( .A1(n391), .A2(n394), .ZN(n596) );
  NAND2_X1 U567 ( .A1(n699), .A2(KEYINPUT34), .ZN(n394) );
  NAND2_X1 U568 ( .A1(n459), .A2(KEYINPUT34), .ZN(n396) );
  INV_X1 U569 ( .A(KEYINPUT15), .ZN(n399) );
  NOR2_X4 U570 ( .A1(n405), .A2(n401), .ZN(n736) );
  AND2_X2 U571 ( .A1(n402), .A2(n424), .ZN(n401) );
  NAND2_X1 U572 ( .A1(n404), .A2(n403), .ZN(n402) );
  INV_X1 U573 ( .A(n741), .ZN(n404) );
  NOR2_X1 U574 ( .A1(n597), .A2(n598), .ZN(n406) );
  NAND2_X1 U575 ( .A1(n410), .A2(n407), .ZN(n483) );
  NAND2_X1 U576 ( .A1(n414), .A2(n408), .ZN(n407) );
  NAND2_X1 U577 ( .A1(n597), .A2(n598), .ZN(n409) );
  NAND2_X1 U578 ( .A1(n413), .A2(KEYINPUT44), .ZN(n412) );
  INV_X1 U579 ( .A(n414), .ZN(n413) );
  XNOR2_X1 U580 ( .A(n465), .B(KEYINPUT88), .ZN(n414) );
  XNOR2_X2 U581 ( .A(n634), .B(n562), .ZN(n641) );
  NOR2_X1 U582 ( .A1(n655), .A2(n359), .ZN(n416) );
  NOR2_X1 U583 ( .A1(n593), .A2(n705), .ZN(n594) );
  XNOR2_X2 U584 ( .A(n444), .B(n361), .ZN(n593) );
  OR2_X2 U585 ( .A1(n587), .A2(n507), .ZN(n511) );
  NAND2_X1 U586 ( .A1(n621), .A2(n506), .ZN(n505) );
  NAND2_X1 U587 ( .A1(n512), .A2(n587), .ZN(n510) );
  XNOR2_X1 U588 ( .A(n505), .B(n504), .ZN(n626) );
  NAND2_X1 U589 ( .A1(n425), .A2(KEYINPUT36), .ZN(n435) );
  NAND2_X1 U590 ( .A1(n633), .A2(n441), .ZN(n425) );
  XNOR2_X1 U591 ( .A(n426), .B(G122), .ZN(n766) );
  XNOR2_X2 U592 ( .A(n596), .B(KEYINPUT35), .ZN(n426) );
  XNOR2_X2 U593 ( .A(n427), .B(G469), .ZN(n625) );
  XNOR2_X1 U594 ( .A(n536), .B(n352), .ZN(n727) );
  NAND2_X1 U595 ( .A1(n705), .A2(n706), .ZN(n601) );
  NAND2_X1 U596 ( .A1(n621), .A2(n691), .ZN(n433) );
  AND2_X1 U597 ( .A1(n633), .A2(n360), .ZN(n439) );
  NAND2_X1 U598 ( .A1(n675), .A2(KEYINPUT36), .ZN(n437) );
  NAND2_X1 U599 ( .A1(n439), .A2(n632), .ZN(n438) );
  NAND2_X1 U600 ( .A1(n632), .A2(n633), .ZN(n644) );
  INV_X1 U601 ( .A(n634), .ZN(n441) );
  NOR2_X2 U602 ( .A1(n603), .A2(n347), .ZN(n444) );
  NAND2_X1 U603 ( .A1(n484), .A2(n486), .ZN(n603) );
  XNOR2_X2 U604 ( .A(n532), .B(n531), .ZN(n556) );
  XNOR2_X1 U605 ( .A(n453), .B(n368), .ZN(G60) );
  NAND2_X1 U606 ( .A1(n455), .A2(n467), .ZN(n453) );
  XNOR2_X1 U607 ( .A(n454), .B(n367), .ZN(G57) );
  NAND2_X1 U608 ( .A1(n466), .A2(n467), .ZN(n454) );
  NAND2_X1 U609 ( .A1(n692), .A2(n691), .ZN(n695) );
  XNOR2_X1 U610 ( .A(n732), .B(n366), .ZN(n455) );
  XNOR2_X1 U611 ( .A(n594), .B(KEYINPUT106), .ZN(n595) );
  NAND2_X1 U612 ( .A1(n515), .A2(n516), .ZN(n509) );
  XNOR2_X1 U613 ( .A(n460), .B(n369), .ZN(G51) );
  NAND2_X1 U614 ( .A1(n660), .A2(n467), .ZN(n460) );
  XNOR2_X2 U615 ( .A(n625), .B(n537), .ZN(n705) );
  XNOR2_X1 U616 ( .A(n462), .B(n461), .ZN(G54) );
  NAND2_X1 U617 ( .A1(n468), .A2(n467), .ZN(n462) );
  XNOR2_X1 U618 ( .A(n653), .B(n365), .ZN(n466) );
  XNOR2_X1 U619 ( .A(n730), .B(n364), .ZN(n468) );
  NOR2_X2 U620 ( .A1(n593), .A2(n591), .ZN(n611) );
  NOR2_X2 U621 ( .A1(n640), .A2(n641), .ZN(n503) );
  NOR2_X1 U622 ( .A1(n554), .A2(n474), .ZN(n471) );
  NAND2_X1 U623 ( .A1(n554), .A2(n477), .ZN(n473) );
  XNOR2_X2 U624 ( .A(n536), .B(n530), .ZN(n554) );
  INV_X1 U625 ( .A(n555), .ZN(n477) );
  NAND2_X1 U626 ( .A1(n482), .A2(n478), .ZN(n637) );
  NOR2_X1 U627 ( .A1(n618), .A2(n481), .ZN(n478) );
  NAND2_X1 U628 ( .A1(n692), .A2(n623), .ZN(n480) );
  OR2_X1 U629 ( .A1(n641), .A2(n357), .ZN(n484) );
  NAND2_X1 U630 ( .A1(n641), .A2(KEYINPUT0), .ZN(n489) );
  XNOR2_X2 U631 ( .A(G128), .B(KEYINPUT65), .ZN(n493) );
  NAND2_X1 U632 ( .A1(n502), .A2(n501), .ZN(n500) );
  AND2_X1 U633 ( .A1(n682), .A2(KEYINPUT83), .ZN(n501) );
  INV_X1 U634 ( .A(n630), .ZN(n506) );
  NAND2_X1 U635 ( .A1(n559), .A2(G137), .ZN(n508) );
  NAND2_X2 U636 ( .A1(n511), .A2(n510), .ZN(n753) );
  XNOR2_X1 U637 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U638 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n517) );
  AND2_X1 U639 ( .A1(n619), .A2(n567), .ZN(n518) );
  XNOR2_X1 U640 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U641 ( .A(n547), .B(n546), .ZN(n738) );
  NOR2_X1 U642 ( .A1(G952), .A2(n748), .ZN(n740) );
  XNOR2_X2 U643 ( .A(n753), .B(G146), .ZN(n536) );
  XNOR2_X1 U644 ( .A(n524), .B(KEYINPUT74), .ZN(n573) );
  NAND2_X1 U645 ( .A1(G210), .A2(n573), .ZN(n525) );
  XOR2_X1 U646 ( .A(n527), .B(n526), .Z(n528) );
  XOR2_X1 U647 ( .A(n572), .B(KEYINPUT91), .Z(n534) );
  NAND2_X1 U648 ( .A1(G227), .A2(n748), .ZN(n533) );
  XNOR2_X1 U649 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U650 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n537) );
  INV_X1 U651 ( .A(n705), .ZN(n612) );
  XNOR2_X1 U652 ( .A(n538), .B(KEYINPUT24), .ZN(n539) );
  NAND2_X1 U653 ( .A1(n748), .A2(G234), .ZN(n541) );
  NAND2_X1 U654 ( .A1(G221), .A2(n583), .ZN(n545) );
  XNOR2_X1 U655 ( .A(n543), .B(n542), .ZN(n544) );
  NOR2_X1 U656 ( .A1(G902), .A2(n738), .ZN(n553) );
  XOR2_X1 U657 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n551) );
  INV_X1 U658 ( .A(n651), .ZN(n548) );
  NAND2_X1 U659 ( .A1(G234), .A2(n548), .ZN(n549) );
  XNOR2_X1 U660 ( .A(KEYINPUT20), .B(n549), .ZN(n589) );
  NAND2_X1 U661 ( .A1(G217), .A2(n589), .ZN(n550) );
  XNOR2_X1 U662 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U663 ( .A(G472), .B(KEYINPUT96), .ZN(n555) );
  INV_X1 U664 ( .A(n631), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G210), .A2(n561), .ZN(n560) );
  NAND2_X1 U666 ( .A1(G214), .A2(n561), .ZN(n691) );
  XNOR2_X1 U667 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n562) );
  NAND2_X1 U668 ( .A1(G234), .A2(G237), .ZN(n563) );
  XNOR2_X1 U669 ( .A(n563), .B(KEYINPUT14), .ZN(n690) );
  NOR2_X1 U670 ( .A1(G902), .A2(n748), .ZN(n565) );
  NOR2_X1 U671 ( .A1(G953), .A2(G952), .ZN(n564) );
  NOR2_X1 U672 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U673 ( .A1(n690), .A2(n566), .ZN(n619) );
  NAND2_X1 U674 ( .A1(G898), .A2(G953), .ZN(n567) );
  XOR2_X1 U675 ( .A(KEYINPUT13), .B(KEYINPUT100), .Z(n569) );
  XNOR2_X1 U676 ( .A(KEYINPUT99), .B(G475), .ZN(n568) );
  INV_X1 U677 ( .A(n570), .ZN(n571) );
  NAND2_X1 U678 ( .A1(n573), .A2(G214), .ZN(n579) );
  XOR2_X1 U679 ( .A(KEYINPUT11), .B(G104), .Z(n575) );
  XNOR2_X1 U680 ( .A(G113), .B(G122), .ZN(n574) );
  XNOR2_X1 U681 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U682 ( .A(G143), .B(KEYINPUT12), .ZN(n577) );
  XNOR2_X1 U683 ( .A(n579), .B(n578), .ZN(n580) );
  NAND2_X1 U684 ( .A1(G217), .A2(n583), .ZN(n584) );
  XNOR2_X1 U685 ( .A(n585), .B(n584), .ZN(n586) );
  NOR2_X1 U686 ( .A1(G902), .A2(n734), .ZN(n588) );
  NAND2_X1 U687 ( .A1(n605), .A2(n607), .ZN(n694) );
  NAND2_X1 U688 ( .A1(G221), .A2(n589), .ZN(n590) );
  XNOR2_X1 U689 ( .A(n590), .B(KEYINPUT21), .ZN(n701) );
  INV_X1 U690 ( .A(KEYINPUT44), .ZN(n598) );
  NAND2_X1 U691 ( .A1(n625), .A2(n706), .ZN(n618) );
  NOR2_X1 U692 ( .A1(n459), .A2(n618), .ZN(n599) );
  XNOR2_X1 U693 ( .A(KEYINPUT94), .B(n599), .ZN(n600) );
  XNOR2_X1 U694 ( .A(KEYINPUT97), .B(n602), .ZN(n711) );
  NOR2_X1 U695 ( .A1(n711), .A2(n459), .ZN(n604) );
  XNOR2_X1 U696 ( .A(n604), .B(KEYINPUT31), .ZN(n677) );
  NAND2_X1 U697 ( .A1(n663), .A2(n677), .ZN(n610) );
  NOR2_X1 U698 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U699 ( .A(KEYINPUT103), .B(n609), .ZN(n678) );
  NAND2_X1 U700 ( .A1(n675), .A2(n678), .ZN(n642) );
  NAND2_X1 U701 ( .A1(n610), .A2(n642), .ZN(n616) );
  XNOR2_X1 U702 ( .A(n611), .B(KEYINPUT86), .ZN(n613) );
  NAND2_X1 U703 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U704 ( .A(n614), .B(KEYINPUT87), .ZN(n615) );
  NAND2_X1 U705 ( .A1(n615), .A2(n622), .ZN(n661) );
  NAND2_X1 U706 ( .A1(n616), .A2(n661), .ZN(n617) );
  NAND2_X1 U707 ( .A1(n619), .A2(n760), .ZN(n620) );
  XOR2_X1 U708 ( .A(KEYINPUT78), .B(n620), .Z(n623) );
  NAND2_X1 U709 ( .A1(n624), .A2(n623), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n640) );
  NOR2_X1 U711 ( .A1(n694), .A2(n695), .ZN(n628) );
  XOR2_X1 U712 ( .A(KEYINPUT41), .B(KEYINPUT109), .Z(n627) );
  XNOR2_X1 U713 ( .A(n628), .B(n627), .ZN(n717) );
  NOR2_X1 U714 ( .A1(n640), .A2(n717), .ZN(n629) );
  NOR2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n633) );
  INV_X1 U716 ( .A(n636), .ZN(n647) );
  NOR2_X1 U717 ( .A1(n647), .A2(n637), .ZN(n638) );
  XOR2_X1 U718 ( .A(KEYINPUT108), .B(n638), .Z(n639) );
  NOR2_X1 U719 ( .A1(n358), .A2(n639), .ZN(n671) );
  INV_X1 U720 ( .A(n642), .ZN(n696) );
  NOR2_X1 U721 ( .A1(n705), .A2(n644), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n645), .A2(n691), .ZN(n646) );
  XNOR2_X1 U723 ( .A(KEYINPUT43), .B(n646), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n682) );
  INV_X1 U725 ( .A(n678), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n681) );
  NAND2_X1 U727 ( .A1(n736), .A2(G472), .ZN(n653) );
  INV_X1 U728 ( .A(KEYINPUT63), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n736), .A2(G210), .ZN(n659) );
  XOR2_X1 U730 ( .A(KEYINPUT89), .B(KEYINPUT55), .Z(n657) );
  XNOR2_X1 U731 ( .A(n655), .B(KEYINPUT54), .ZN(n656) );
  XNOR2_X1 U732 ( .A(G101), .B(n661), .ZN(G3) );
  NOR2_X1 U733 ( .A1(n675), .A2(n663), .ZN(n662) );
  XOR2_X1 U734 ( .A(G104), .B(n662), .Z(G6) );
  NOR2_X1 U735 ( .A1(n663), .A2(n678), .ZN(n667) );
  XOR2_X1 U736 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n665) );
  XNOR2_X1 U737 ( .A(G107), .B(KEYINPUT113), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(G9) );
  XOR2_X1 U740 ( .A(n668), .B(G110), .Z(G12) );
  NOR2_X1 U741 ( .A1(n678), .A2(n673), .ZN(n670) );
  XNOR2_X1 U742 ( .A(G128), .B(KEYINPUT29), .ZN(n669) );
  XNOR2_X1 U743 ( .A(n670), .B(n669), .ZN(G30) );
  XOR2_X1 U744 ( .A(G143), .B(n671), .Z(n672) );
  XNOR2_X1 U745 ( .A(KEYINPUT114), .B(n672), .ZN(G45) );
  NOR2_X1 U746 ( .A1(n675), .A2(n673), .ZN(n674) );
  XOR2_X1 U747 ( .A(G146), .B(n674), .Z(G48) );
  NOR2_X1 U748 ( .A1(n675), .A2(n677), .ZN(n676) );
  XOR2_X1 U749 ( .A(G113), .B(n676), .Z(G15) );
  NOR2_X1 U750 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U751 ( .A(G116), .B(n679), .Z(G18) );
  XOR2_X1 U752 ( .A(G134), .B(KEYINPUT115), .Z(n680) );
  XNOR2_X1 U753 ( .A(n681), .B(n680), .ZN(G36) );
  XNOR2_X1 U754 ( .A(G140), .B(n682), .ZN(G42) );
  XNOR2_X1 U755 ( .A(KEYINPUT79), .B(n683), .ZN(n685) );
  NAND2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n717), .A2(n699), .ZN(n686) );
  XNOR2_X1 U758 ( .A(KEYINPUT120), .B(n686), .ZN(n687) );
  NOR2_X1 U759 ( .A1(G953), .A2(n687), .ZN(n688) );
  NAND2_X1 U760 ( .A1(n689), .A2(n688), .ZN(n725) );
  NAND2_X1 U761 ( .A1(G952), .A2(n690), .ZN(n722) );
  NOR2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n700) );
  NOR2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n719) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U768 ( .A(n703), .B(KEYINPUT116), .ZN(n704) );
  XNOR2_X1 U769 ( .A(KEYINPUT49), .B(n704), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U771 ( .A(KEYINPUT50), .B(n707), .ZN(n708) );
  NOR2_X1 U772 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n715) );
  XOR2_X1 U774 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n713) );
  XNOR2_X1 U775 ( .A(KEYINPUT51), .B(n713), .ZN(n714) );
  XNOR2_X1 U776 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U777 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U778 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U779 ( .A(n720), .B(KEYINPUT52), .ZN(n721) );
  NOR2_X1 U780 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U781 ( .A(KEYINPUT119), .B(n723), .Z(n724) );
  NOR2_X1 U782 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U783 ( .A(KEYINPUT53), .B(n726), .ZN(G75) );
  XNOR2_X1 U784 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n729) );
  XNOR2_X1 U785 ( .A(n727), .B(KEYINPUT57), .ZN(n728) );
  NAND2_X1 U786 ( .A1(n736), .A2(G469), .ZN(n730) );
  NAND2_X1 U787 ( .A1(n736), .A2(G475), .ZN(n732) );
  NAND2_X1 U788 ( .A1(G478), .A2(n736), .ZN(n733) );
  XNOR2_X1 U789 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U790 ( .A1(n740), .A2(n735), .ZN(G63) );
  NAND2_X1 U791 ( .A1(G217), .A2(n736), .ZN(n737) );
  XNOR2_X1 U792 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U793 ( .A1(n740), .A2(n739), .ZN(G66) );
  NOR2_X1 U794 ( .A1(G953), .A2(n741), .ZN(n742) );
  XNOR2_X1 U795 ( .A(n742), .B(KEYINPUT125), .ZN(n747) );
  NAND2_X1 U796 ( .A1(G224), .A2(G953), .ZN(n743) );
  XNOR2_X1 U797 ( .A(n743), .B(KEYINPUT124), .ZN(n744) );
  XNOR2_X1 U798 ( .A(KEYINPUT61), .B(n744), .ZN(n745) );
  NAND2_X1 U799 ( .A1(n745), .A2(G898), .ZN(n746) );
  NAND2_X1 U800 ( .A1(n747), .A2(n746), .ZN(n752) );
  OR2_X1 U801 ( .A1(n748), .A2(G898), .ZN(n750) );
  NAND2_X1 U802 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U803 ( .A(n752), .B(n751), .Z(G69) );
  BUF_X1 U804 ( .A(n753), .Z(n754) );
  XNOR2_X1 U805 ( .A(n755), .B(n754), .ZN(n758) );
  XNOR2_X1 U806 ( .A(n758), .B(n756), .ZN(n757) );
  NOR2_X1 U807 ( .A1(G953), .A2(n757), .ZN(n762) );
  XOR2_X1 U808 ( .A(G227), .B(n758), .Z(n759) );
  NOR2_X1 U809 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U810 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U811 ( .A(KEYINPUT126), .B(n763), .ZN(G72) );
  XNOR2_X1 U812 ( .A(n764), .B(G125), .ZN(n765) );
  XNOR2_X1 U813 ( .A(n765), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U814 ( .A(n766), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U815 ( .A(n767), .B(G137), .Z(G39) );
  XOR2_X1 U816 ( .A(n768), .B(G119), .Z(G21) );
  XOR2_X1 U817 ( .A(n769), .B(G131), .Z(G33) );
endmodule

