//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n191), .A2(G140), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n193), .A2(new_n194), .A3(G146), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(KEYINPUT70), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT69), .B(G140), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(new_n191), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n200), .A2(KEYINPUT69), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(KEYINPUT69), .ZN(new_n202));
  OAI211_X1 g016(.A(KEYINPUT70), .B(G125), .C1(new_n201), .C2(new_n202), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n199), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n196), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G953), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT68), .A2(G237), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT68), .A2(G237), .ZN(new_n209));
  OAI211_X1 g023(.A(G214), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(KEYINPUT81), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(G237), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G214), .A4(new_n207), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT82), .B1(new_n217), .B2(new_n211), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n219));
  AOI211_X1 g033(.A(new_n219), .B(G143), .C1(new_n213), .C2(new_n216), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n212), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(KEYINPUT18), .A2(G131), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n206), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n221), .A2(G131), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(KEYINPUT18), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n199), .A2(KEYINPUT19), .A3(new_n203), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT19), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n193), .B2(new_n194), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n205), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT83), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n199), .A2(KEYINPUT16), .A3(new_n203), .ZN(new_n232));
  OR3_X1    g046(.A1(new_n191), .A2(KEYINPUT16), .A3(G140), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(G146), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT83), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n229), .A2(new_n235), .A3(new_n205), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n231), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n221), .A2(G131), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n239), .B(new_n212), .C1(new_n218), .C2(new_n220), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n190), .B1(new_n225), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n221), .A2(KEYINPUT18), .A3(G131), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(new_n206), .C1(new_n221), .C2(new_n222), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT17), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n238), .A2(new_n245), .A3(new_n240), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n221), .A2(KEYINPUT17), .A3(G131), .ZN(new_n247));
  AOI21_X1  g061(.A(G146), .B1(new_n232), .B2(new_n233), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n234), .B1(new_n248), .B2(KEYINPUT71), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n250));
  AOI211_X1 g064(.A(new_n250), .B(G146), .C1(new_n232), .C2(new_n233), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n244), .B(new_n189), .C1(new_n246), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n242), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n256));
  NOR2_X1   g070(.A1(G475), .A2(G902), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT84), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n257), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT20), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT84), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n255), .A2(new_n262), .A3(new_n256), .A4(new_n257), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  INV_X1    g079(.A(new_n254), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n238), .A2(new_n245), .A3(new_n240), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n247), .A3(new_n252), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n189), .B1(new_n268), .B2(new_n244), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n265), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G475), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT14), .ZN(new_n273));
  INV_X1    g087(.A(G116), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(G122), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(G122), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(KEYINPUT14), .B2(new_n276), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n211), .A2(G128), .ZN(new_n279));
  INV_X1    g093(.A(G128), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G143), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n281), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G134), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n278), .A2(G107), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G122), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G116), .ZN(new_n288));
  INV_X1    g102(.A(G107), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n276), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(KEYINPUT85), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n280), .A2(G143), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(KEYINPUT13), .B2(new_n281), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n293), .A2(KEYINPUT13), .ZN(new_n295));
  OAI21_X1  g109(.A(G134), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n288), .A2(new_n276), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G107), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n290), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n283), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT9), .B(G234), .ZN(new_n301));
  INV_X1    g115(.A(G217), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n301), .A2(new_n302), .A3(G953), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n292), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n292), .B2(new_n300), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G902), .ZN(new_n307));
  INV_X1    g121(.A(G478), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(KEYINPUT15), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(KEYINPUT15), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n313), .B1(new_n306), .B2(G902), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(G234), .A2(G237), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(G952), .A3(new_n207), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(G902), .A3(G953), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT21), .B(G898), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n289), .A2(G104), .ZN(new_n327));
  AND2_X1   g141(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT76), .B(G101), .Z(new_n330));
  NAND2_X1  g144(.A1(new_n188), .A2(G107), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n188), .A2(G107), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n329), .A2(new_n330), .A3(new_n331), .A4(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n289), .A2(G104), .ZN(new_n336));
  OAI21_X1  g150(.A(G101), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n205), .A2(G143), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n211), .A2(G146), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(KEYINPUT1), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(G128), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n339), .B(new_n340), .C1(KEYINPUT1), .C2(new_n280), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OR3_X1    g159(.A1(new_n338), .A2(KEYINPUT10), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT10), .B1(new_n338), .B2(new_n345), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT66), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT11), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n282), .B2(G137), .ZN(new_n351));
  INV_X1    g165(.A(G137), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT11), .A3(G134), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n282), .A2(G137), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G131), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n351), .A2(new_n353), .A3(new_n239), .A4(new_n354), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n349), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n349), .A3(new_n357), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G101), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n336), .B1(new_n333), .B2(new_n332), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(new_n329), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n366));
  NOR2_X1   g180(.A1(KEYINPUT0), .A2(G128), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT0), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(new_n280), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n341), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n339), .B(new_n340), .C1(new_n368), .C2(new_n280), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n365), .A2(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n331), .B1(new_n326), .B2(new_n327), .ZN(new_n373));
  NAND2_X1  g187(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n333), .B1(new_n332), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G101), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT4), .A3(new_n335), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n372), .A2(KEYINPUT77), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT77), .B1(new_n372), .B2(new_n377), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n348), .B(new_n362), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n345), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n335), .A3(new_n337), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n338), .A2(new_n345), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n356), .A2(new_n357), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(KEYINPUT12), .A3(new_n385), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n382), .A2(new_n383), .B1(new_n359), .B2(new_n360), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(KEYINPUT12), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n380), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G110), .B(G140), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n207), .A2(G227), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n390), .B(new_n391), .Z(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n348), .B1(new_n378), .B2(new_n379), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n361), .ZN(new_n395));
  INV_X1    g209(.A(new_n392), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n380), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G469), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n397), .A3(new_n398), .A4(new_n265), .ZN(new_n399));
  NAND2_X1  g213(.A1(G469), .A2(G902), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n389), .A2(new_n396), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n395), .A2(new_n380), .A3(new_n392), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n399), .B(new_n400), .C1(new_n398), .C2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G221), .B1(new_n301), .B2(G902), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n405), .B(KEYINPUT74), .Z(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G224), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(G953), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n343), .A2(new_n191), .A3(new_n344), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n191), .B1(new_n370), .B2(new_n371), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT7), .B(new_n410), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n413), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n410), .A2(KEYINPUT7), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT8), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n335), .A2(new_n337), .ZN(new_n420));
  XNOR2_X1  g234(.A(G116), .B(G119), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT5), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n274), .A2(KEYINPUT5), .A3(G119), .ZN(new_n423));
  INV_X1    g237(.A(G113), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(KEYINPUT2), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT2), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G113), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n430), .A2(new_n421), .A3(KEYINPUT65), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT65), .B1(new_n430), .B2(new_n421), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n419), .B1(new_n420), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT65), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n427), .A2(new_n429), .ZN(new_n436));
  XOR2_X1   g250(.A(G116), .B(G119), .Z(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n430), .A2(new_n421), .A3(KEYINPUT65), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n422), .A2(KEYINPUT79), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT79), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n421), .A2(new_n442), .A3(KEYINPUT5), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n443), .A3(new_n425), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n338), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n414), .B(new_n417), .C1(new_n434), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n365), .A2(new_n366), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n436), .A2(new_n437), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n431), .B2(new_n432), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n377), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n440), .A2(new_n335), .A3(new_n337), .A4(new_n426), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n450), .A2(new_n451), .A3(new_n418), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n265), .B1(new_n446), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT80), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n450), .A2(new_n451), .ZN(new_n456));
  INV_X1    g270(.A(new_n418), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n451), .A3(new_n418), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(KEYINPUT6), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n412), .A2(new_n413), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(new_n409), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n456), .A2(new_n463), .A3(new_n457), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n460), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT80), .B(new_n265), .C1(new_n446), .C2(new_n452), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n455), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G210), .B1(G237), .B2(G902), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n455), .A2(new_n465), .A3(new_n468), .A4(new_n466), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G214), .B1(G237), .B2(G902), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT78), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n407), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n272), .A2(KEYINPUT87), .A3(new_n325), .A4(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n476), .A2(new_n264), .A3(new_n271), .A4(new_n325), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT22), .B(G137), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n207), .A2(G221), .A3(G234), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n280), .A2(G119), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n280), .A2(KEYINPUT23), .A3(G119), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT23), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n280), .A2(G119), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G110), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n485), .A2(new_n489), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G110), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n249), .B2(new_n251), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT72), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(new_n496), .C1(new_n249), .C2(new_n251), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n490), .A2(new_n491), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n493), .A2(new_n494), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n195), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n504), .A2(new_n234), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n484), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n505), .B(new_n483), .C1(new_n498), .C2(new_n500), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n265), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT25), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n302), .B1(G234), .B2(new_n265), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT25), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n512), .B(new_n265), .C1(new_n507), .C2(new_n508), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n507), .ZN(new_n515));
  INV_X1    g329(.A(new_n508), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n511), .A2(G902), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT73), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G472), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n370), .A2(new_n371), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n356), .A2(new_n349), .A3(new_n357), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n358), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n354), .A2(KEYINPUT64), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n352), .A2(G134), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n352), .A2(KEYINPUT64), .A3(G134), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n239), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n357), .ZN(new_n532));
  OR3_X1    g346(.A1(new_n531), .A2(new_n345), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n523), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n531), .A2(new_n345), .A3(new_n532), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n356), .A2(new_n357), .B1(new_n370), .B2(new_n371), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n535), .A2(KEYINPUT30), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n449), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n214), .A2(G210), .A3(new_n207), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT27), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT26), .B(G101), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT67), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n449), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n440), .A2(KEYINPUT67), .A3(new_n448), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n526), .A2(new_n533), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n538), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n547), .A2(KEYINPUT31), .ZN(new_n548));
  INV_X1    g362(.A(new_n542), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT28), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n449), .B1(new_n535), .B2(new_n536), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n550), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n535), .B1(new_n361), .B2(new_n524), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n545), .A2(new_n544), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT28), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n549), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT31), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n538), .A2(new_n558), .A3(new_n542), .A4(new_n546), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n522), .B(new_n265), .C1(new_n548), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT32), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n547), .A2(KEYINPUT31), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n559), .A3(new_n557), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT32), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n522), .A4(new_n265), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n538), .A2(new_n546), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n549), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT29), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n552), .A2(new_n556), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(new_n549), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n526), .A2(new_n533), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n554), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n546), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n556), .B1(new_n574), .B2(KEYINPUT28), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n549), .A2(new_n569), .ZN(new_n576));
  AOI21_X1  g390(.A(G902), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n562), .A2(new_n566), .B1(G472), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n521), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n477), .A2(new_n480), .A3(new_n580), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(new_n330), .Z(G3));
  INV_X1    g396(.A(KEYINPUT88), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n470), .B1(new_n583), .B2(new_n471), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n471), .A2(new_n583), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n473), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT89), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n455), .A2(new_n465), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n590), .A2(KEYINPUT88), .A3(new_n468), .A4(new_n466), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(new_n470), .A3(new_n585), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(KEYINPUT89), .A3(new_n473), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(new_n324), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n265), .A2(G478), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n305), .A2(KEYINPUT90), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  OR3_X1    g412(.A1(new_n306), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n306), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT91), .B1(new_n307), .B2(G478), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(KEYINPUT91), .B2(new_n601), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n272), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n564), .A2(new_n265), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(G472), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n608), .A2(new_n561), .ZN(new_n609));
  INV_X1    g423(.A(new_n407), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n521), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n595), .A2(new_n606), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  XNOR2_X1  g429(.A(new_n324), .B(KEYINPUT93), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n594), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT92), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n268), .A2(new_n244), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n190), .ZN(new_n620));
  AOI21_X1  g434(.A(G902), .B1(new_n620), .B2(new_n254), .ZN(new_n621));
  INV_X1    g435(.A(G475), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n270), .A2(KEYINPUT92), .A3(G475), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n317), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n617), .A2(new_n612), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NAND2_X1  g446(.A1(new_n501), .A2(new_n506), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n484), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT94), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n633), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n519), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n514), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n477), .A2(new_n480), .A3(new_n609), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT37), .B(G110), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT95), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(G12));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n320), .B1(new_n322), .B2(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n625), .A2(new_n628), .A3(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n592), .A2(KEYINPUT89), .A3(new_n473), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT89), .B1(new_n592), .B2(new_n473), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n578), .A2(G472), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n562), .A2(new_n566), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n649), .A2(new_n650), .B1(new_n514), .B2(new_n637), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n645), .A2(new_n648), .A3(new_n610), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT96), .B(G128), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G30));
  INV_X1    g468(.A(new_n317), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n264), .B2(new_n271), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n644), .B(KEYINPUT39), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n610), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT99), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n472), .B(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n522), .B1(new_n574), .B2(new_n549), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n547), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n522), .A2(new_n265), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT98), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n562), .B2(new_n566), .ZN(new_n672));
  INV_X1    g486(.A(new_n473), .ZN(new_n673));
  NOR4_X1   g487(.A1(new_n665), .A2(new_n672), .A3(new_n638), .A4(new_n673), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n662), .B(new_n674), .C1(new_n661), .C2(new_n660), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  AOI211_X1 g490(.A(new_n605), .B(new_n644), .C1(new_n264), .C2(new_n271), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n677), .A2(new_n610), .A3(new_n648), .A4(new_n651), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  NAND2_X1  g493(.A1(new_n393), .A2(new_n397), .ZN(new_n680));
  OAI21_X1  g494(.A(G469), .B1(new_n680), .B2(G902), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n399), .A3(new_n405), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n521), .A2(new_n579), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n595), .A2(new_n606), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NAND3_X1  g500(.A1(new_n617), .A2(new_n629), .A3(new_n683), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n650), .A2(new_n649), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(new_n589), .A3(new_n638), .A4(new_n593), .ZN(new_n691));
  INV_X1    g505(.A(new_n682), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n264), .A2(new_n271), .A3(new_n325), .A4(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n689), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n693), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n695), .A2(KEYINPUT100), .A3(new_n648), .A4(new_n651), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  OAI211_X1 g512(.A(new_n563), .B(new_n559), .C1(new_n542), .C2(new_n575), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n522), .A2(new_n265), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT101), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n607), .A2(G472), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n521), .A2(new_n682), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n617), .A2(new_n656), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NOR3_X1   g520(.A1(new_n646), .A2(new_n647), .A3(new_n682), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n703), .B1(new_n514), .B2(new_n637), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n677), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT102), .B(G125), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G27));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n264), .A2(new_n271), .ZN(new_n713));
  INV_X1    g527(.A(new_n605), .ZN(new_n714));
  INV_X1    g528(.A(new_n644), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n513), .A2(new_n511), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n717), .A2(new_n510), .B1(new_n519), .B2(new_n517), .ZN(new_n718));
  AND4_X1   g532(.A1(new_n405), .A2(new_n470), .A3(new_n471), .A4(new_n473), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n402), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n395), .A2(KEYINPUT103), .A3(new_n380), .A4(new_n392), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n401), .A3(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n399), .B(new_n400), .C1(new_n723), .C2(new_n398), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n718), .A2(new_n690), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n712), .B1(new_n716), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n719), .A2(new_n724), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n521), .A2(new_n579), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n677), .A2(new_n729), .A3(KEYINPUT42), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n645), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  INV_X1    g548(.A(new_n405), .ZN(new_n735));
  INV_X1    g549(.A(new_n399), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n398), .B1(new_n403), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n723), .B2(new_n737), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n739), .A2(new_n400), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(KEYINPUT46), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n736), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n742), .B1(new_n740), .B2(KEYINPUT46), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(KEYINPUT46), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n735), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n472), .A2(new_n673), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n658), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n713), .A2(new_n605), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(KEYINPUT105), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n713), .B2(new_n605), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n609), .B1(new_n514), .B2(new_n637), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT44), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(KEYINPUT44), .A3(new_n756), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  XNOR2_X1  g578(.A(new_n747), .B(KEYINPUT47), .ZN(new_n765));
  INV_X1    g579(.A(new_n748), .ZN(new_n766));
  NOR4_X1   g580(.A1(new_n716), .A2(new_n718), .A3(new_n690), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT107), .B(G140), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G42));
  AND2_X1   g584(.A1(new_n755), .A2(new_n320), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n681), .A2(new_n399), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n766), .A2(new_n735), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n708), .ZN(new_n775));
  INV_X1    g589(.A(new_n672), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n521), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n320), .A3(new_n773), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n272), .A2(new_n605), .ZN(new_n779));
  OAI22_X1  g593(.A1(new_n774), .A2(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n772), .B(KEYINPUT108), .Z(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n406), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n765), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n521), .A2(new_n703), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n771), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n766), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n780), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n682), .B2(new_n473), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n692), .A2(KEYINPUT111), .A3(new_n673), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n665), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n771), .A2(new_n785), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n788), .A2(KEYINPUT51), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT51), .B1(new_n788), .B2(new_n795), .ZN(new_n797));
  INV_X1    g611(.A(new_n707), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n786), .A2(KEYINPUT112), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n606), .ZN(new_n800));
  OAI211_X1 g614(.A(G952), .B(new_n207), .C1(new_n778), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n771), .A2(new_n580), .A3(new_n773), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT48), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT112), .B1(new_n786), .B2(new_n798), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OR3_X1    g620(.A1(new_n796), .A2(new_n797), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n735), .A2(new_n644), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n514), .A2(new_n637), .A3(new_n724), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n648), .A2(new_n810), .A3(new_n776), .A4(new_n656), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n678), .A2(new_n709), .A3(new_n652), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n812), .A2(KEYINPUT52), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(KEYINPUT52), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT110), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n475), .A2(new_n616), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n264), .A2(new_n271), .A3(new_n317), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n817), .A2(KEYINPUT109), .B1(new_n713), .B2(new_n714), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n713), .A2(KEYINPUT109), .A3(new_n714), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n612), .B(new_n816), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n697), .A2(new_n820), .A3(new_n639), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n702), .A2(new_n719), .A3(new_n724), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n713), .A2(new_n822), .A3(new_n714), .A4(new_n715), .ZN(new_n823));
  INV_X1    g637(.A(new_n625), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n261), .A2(new_n258), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n317), .A2(new_n644), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n470), .A3(new_n471), .A4(new_n473), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n407), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n824), .A2(new_n690), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n638), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n731), .A2(new_n831), .A3(new_n733), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n581), .A2(new_n684), .A3(new_n687), .A4(new_n705), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n821), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n709), .A2(new_n652), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n836), .A3(new_n678), .A4(new_n811), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n812), .A2(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n709), .A2(new_n652), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT110), .B1(new_n839), .B2(KEYINPUT52), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n815), .A2(KEYINPUT53), .A3(new_n834), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n697), .A2(new_n820), .A3(new_n639), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n731), .A2(new_n733), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n581), .A2(new_n684), .A3(new_n687), .A4(new_n705), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n844), .A2(new_n846), .A3(new_n847), .A4(new_n831), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n837), .A2(new_n838), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n843), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n842), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n815), .A2(new_n843), .A3(new_n834), .A4(new_n841), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n848), .A2(new_n849), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n855), .B(KEYINPUT54), .C1(new_n843), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n807), .A2(new_n858), .B1(G952), .B2(G953), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n781), .B(KEYINPUT49), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n665), .A2(new_n406), .A3(new_n474), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n750), .A3(new_n777), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(G75));
  NAND3_X1  g677(.A1(new_n851), .A2(G210), .A3(G902), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n460), .A2(new_n464), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT113), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n462), .B(KEYINPUT55), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n870), .B2(new_n871), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n207), .A2(G952), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G51));
  NAND3_X1  g690(.A1(new_n852), .A2(KEYINPUT114), .A3(new_n853), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n851), .B2(KEYINPUT54), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n400), .B(KEYINPUT57), .Z(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n680), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n739), .B(KEYINPUT115), .Z(new_n886));
  NAND3_X1  g700(.A1(new_n851), .A2(G902), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n875), .B1(new_n885), .B2(new_n887), .ZN(G54));
  INV_X1    g702(.A(new_n875), .ZN(new_n889));
  AND4_X1   g703(.A1(KEYINPUT58), .A2(new_n851), .A3(G475), .A4(G902), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(new_n255), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n255), .B2(new_n890), .ZN(G60));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT59), .Z(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n854), .B2(new_n857), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n599), .A2(new_n600), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n889), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n599), .B2(new_n600), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n881), .B2(new_n898), .ZN(G63));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT117), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT60), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n851), .A2(new_n636), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT118), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n851), .A2(new_n902), .ZN(new_n905));
  INV_X1    g719(.A(new_n517), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n851), .A2(new_n908), .A3(new_n636), .A4(new_n902), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n904), .A2(new_n907), .A3(new_n889), .A4(new_n909), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n910), .A2(KEYINPUT116), .A3(KEYINPUT61), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT61), .B1(new_n910), .B2(KEYINPUT116), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(G66));
  NOR3_X1   g727(.A1(new_n323), .A2(new_n408), .A3(new_n207), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n844), .A2(new_n847), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT119), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n916), .B2(new_n207), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n869), .B1(G898), .B2(new_n207), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT121), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT120), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n917), .B(new_n920), .ZN(G69));
  AOI21_X1  g735(.A(new_n207), .B1(G227), .B2(G900), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT123), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n534), .A2(new_n537), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n229), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n846), .A2(KEYINPUT125), .ZN(new_n927));
  INV_X1    g741(.A(new_n580), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n928), .A2(new_n657), .A3(new_n594), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n747), .A2(new_n658), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n768), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(KEYINPUT125), .B2(new_n846), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n835), .A2(new_n678), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n763), .A2(KEYINPUT124), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT124), .B1(new_n763), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n926), .B1(new_n936), .B2(new_n207), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n926), .A2(new_n207), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n933), .A2(new_n675), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT62), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n818), .A2(new_n819), .ZN(new_n941));
  NOR4_X1   g755(.A1(new_n941), .A2(new_n928), .A3(new_n659), .A4(new_n766), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n765), .B2(new_n767), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n763), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  OR3_X1    g759(.A1(new_n940), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n940), .B2(new_n944), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n938), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n923), .B1(new_n937), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(G227), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n643), .B1(new_n926), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n207), .B2(new_n951), .ZN(G72));
  NAND2_X1  g766(.A1(new_n567), .A2(new_n542), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n946), .A2(new_n916), .A3(new_n947), .ZN(new_n954));
  XNOR2_X1  g768(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n669), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n932), .B(new_n916), .C1(new_n935), .C2(new_n934), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n542), .B(new_n567), .C1(new_n958), .C2(new_n956), .ZN(new_n959));
  INV_X1    g773(.A(new_n956), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n568), .B2(new_n547), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n855), .B(new_n961), .C1(new_n856), .C2(new_n843), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n889), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n957), .A2(new_n959), .A3(new_n963), .ZN(G57));
endmodule


