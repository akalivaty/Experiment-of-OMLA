//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n555, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(G137), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n466), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n475), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n463), .A2(new_n465), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT69), .ZN(new_n483));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n471), .C2(G112), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n480), .A2(new_n471), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n466), .A2(G138), .A3(new_n471), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n489), .B(new_n491), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n466), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n493));
  INV_X1    g068(.A(G102), .ZN(new_n494));
  OAI22_X1  g069(.A1(new_n493), .A2(new_n467), .B1(new_n494), .B2(new_n474), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  NAND2_X1  g072(.A1(G75), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n506), .B(KEYINPUT71), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n509), .A2(new_n511), .A3(new_n500), .A4(new_n502), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n509), .A2(new_n511), .A3(G543), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(G88), .B1(new_n515), .B2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n507), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NOR2_X1   g093(.A1(new_n501), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT72), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n500), .A2(new_n502), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n513), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n515), .A2(G51), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n525), .A2(new_n526), .A3(new_n528), .A4(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n521), .B2(new_n523), .ZN(new_n533));
  AND2_X1   g108(.A1(G77), .A2(G543), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n513), .A2(G90), .B1(new_n515), .B2(G52), .ZN(new_n538));
  OAI211_X1 g113(.A(KEYINPUT73), .B(G651), .C1(new_n533), .C2(new_n534), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(G171));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  INV_X1    g117(.A(G43), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n512), .A2(new_n542), .B1(new_n514), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n500), .A2(new_n502), .A3(new_n522), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n522), .B1(new_n500), .B2(new_n502), .ZN(new_n546));
  OAI21_X1  g121(.A(G56), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n544), .B1(new_n549), .B2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT74), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n514), .B2(new_n560), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n503), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(G651), .A2(new_n565), .B1(new_n513), .B2(G91), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n515), .A2(KEYINPUT76), .A3(G53), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n540), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n537), .A2(KEYINPUT77), .A3(new_n538), .A4(new_n539), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G301));
  OAI21_X1  g149(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n513), .A2(G87), .B1(new_n515), .B2(G49), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n503), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n513), .A2(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n515), .A2(G48), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n508), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n512), .A2(new_n587), .B1(new_n514), .B2(new_n588), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n586), .A2(KEYINPUT78), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT78), .B1(new_n586), .B2(new_n589), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n512), .A2(KEYINPUT10), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT10), .B1(new_n512), .B2(new_n593), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n503), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(new_n515), .B2(G54), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G301), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n603), .ZN(G284));
  XOR2_X1   g181(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n562), .A2(new_n566), .ZN(new_n609));
  INV_X1    g184(.A(new_n569), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n608), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n608), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(new_n602), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  INV_X1    g191(.A(new_n544), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n508), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n603), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n614), .A2(new_n615), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT80), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n620), .B1(new_n622), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g199(.A1(new_n480), .A2(new_n474), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  AOI22_X1  g203(.A1(G123), .A2(new_n485), .B1(new_n481), .B2(G135), .ZN(new_n629));
  OAI221_X1 g204(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n471), .C2(G111), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(new_n632), .ZN(G156));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT82), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2430), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  OAI21_X1  g223(.A(new_n634), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G14), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n647), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n642), .B(new_n645), .ZN(new_n652));
  INV_X1    g227(.A(new_n648), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT83), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2096), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  AOI21_X1  g241(.A(KEYINPUT18), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n674), .A2(KEYINPUT84), .ZN(new_n675));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(KEYINPUT84), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n671), .A2(new_n673), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n679), .A2(new_n680), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(new_n674), .ZN(new_n684));
  OAI221_X1 g259(.A(new_n682), .B1(new_n680), .B2(new_n679), .C1(new_n677), .C2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1986), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT85), .B(G1981), .Z(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(G229));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G35), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G162), .B2(new_n693), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G2090), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT99), .Z(new_n698));
  AND2_X1   g273(.A1(KEYINPUT30), .A2(G28), .ZN(new_n699));
  NOR2_X1   g274(.A1(KEYINPUT30), .A2(G28), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n693), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT31), .B(G11), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n701), .B(new_n702), .C1(new_n631), .C2(new_n693), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT97), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT27), .B(G1996), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n693), .A2(G32), .ZN(new_n706));
  AOI22_X1  g281(.A1(G129), .A2(new_n485), .B1(new_n481), .B2(G141), .ZN(new_n707));
  NAND3_X1  g282(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT26), .Z(new_n709));
  INV_X1    g284(.A(G105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n707), .B(new_n709), .C1(new_n710), .C2(new_n474), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT95), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT96), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n706), .B1(new_n713), .B2(new_n693), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n698), .B(new_n704), .C1(new_n705), .C2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n696), .A2(G2090), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT98), .Z(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G4), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n614), .B2(new_n718), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1348), .Z(new_n721));
  NAND2_X1  g296(.A1(G168), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G16), .B2(G21), .ZN(new_n723));
  INV_X1    g298(.A(G1966), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G34), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(new_n693), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G160), .B2(new_n693), .ZN(new_n728));
  OAI22_X1  g303(.A1(new_n723), .A2(new_n724), .B1(new_n728), .B2(G2084), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n724), .B2(new_n723), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n717), .A2(new_n721), .A3(new_n730), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n728), .A2(G2084), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n481), .A2(G139), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT92), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n734), .B(new_n737), .C1(new_n471), .C2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT93), .ZN(new_n740));
  MUX2_X1   g315(.A(G33), .B(new_n740), .S(G29), .Z(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(G2072), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n693), .A2(G26), .ZN(new_n743));
  INV_X1    g318(.A(new_n481), .ZN(new_n744));
  INV_X1    g319(.A(G140), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(G2104), .B1(new_n471), .B2(G116), .ZN(new_n747));
  NOR2_X1   g322(.A1(G104), .A2(G2105), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(KEYINPUT90), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(KEYINPUT90), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n746), .B(new_n751), .C1(G128), .C2(new_n485), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n743), .B1(new_n752), .B2(new_n693), .ZN(new_n753));
  MUX2_X1   g328(.A(new_n743), .B(new_n753), .S(KEYINPUT28), .Z(new_n754));
  INV_X1    g329(.A(G2067), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n718), .A2(KEYINPUT23), .A3(G20), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT23), .ZN(new_n758));
  INV_X1    g333(.A(G20), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G16), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n760), .C1(new_n611), .C2(new_n718), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1956), .ZN(new_n762));
  NAND2_X1  g337(.A1(G171), .A2(G16), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G5), .B2(G16), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n762), .B1(G1961), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n714), .A2(new_n705), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n742), .A2(new_n756), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n715), .A2(new_n731), .A3(new_n732), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n693), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n693), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G2078), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n718), .A2(G22), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G166), .B2(new_n718), .ZN(new_n774));
  INV_X1    g349(.A(G1971), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G6), .B(G305), .S(G16), .Z(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT32), .B(G1981), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT87), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n777), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G16), .A2(G23), .ZN(new_n781));
  INV_X1    g356(.A(G288), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT33), .B(G1976), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n776), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G24), .B(G290), .S(G16), .Z(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1986), .Z(new_n790));
  AOI22_X1  g365(.A1(G119), .A2(new_n485), .B1(new_n481), .B2(G131), .ZN(new_n791));
  OAI221_X1 g366(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n471), .C2(G107), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G25), .B(new_n793), .S(G29), .Z(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT35), .B(G1991), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n788), .A2(new_n790), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n799));
  OR2_X1    g374(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n798), .A2(new_n799), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n769), .A2(new_n772), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n765), .A2(G1961), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G19), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n550), .B2(G16), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT89), .B(G1341), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n803), .A2(new_n804), .A3(new_n809), .ZN(G311));
  INV_X1    g385(.A(G311), .ZN(G150));
  OAI21_X1  g386(.A(G67), .B1(new_n545), .B2(new_n546), .ZN(new_n812));
  NAND2_X1  g387(.A1(G80), .A2(G543), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n508), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT100), .ZN(new_n815));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  INV_X1    g391(.A(G55), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n512), .A2(new_n816), .B1(new_n514), .B2(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n814), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G67), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n521), .B2(new_n523), .ZN(new_n821));
  INV_X1    g396(.A(new_n813), .ZN(new_n822));
  OAI21_X1  g397(.A(G651), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n818), .ZN(new_n824));
  AOI21_X1  g399(.A(KEYINPUT100), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n614), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT39), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n619), .B1(new_n819), .B2(new_n825), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n550), .B1(new_n814), .B2(new_n818), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n815), .B1(new_n814), .B2(new_n818), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n823), .A2(KEYINPUT100), .A3(new_n824), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n550), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n812), .A2(new_n813), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n818), .B1(new_n839), .B2(G651), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n619), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n838), .A2(KEYINPUT101), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n831), .B(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n828), .B1(new_n844), .B2(G860), .ZN(G145));
  NAND2_X1  g420(.A1(new_n740), .A2(new_n712), .ZN(new_n846));
  INV_X1    g421(.A(new_n713), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(new_n740), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n752), .B(new_n496), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n849), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n846), .B(new_n851), .C1(new_n847), .C2(new_n740), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n626), .B(new_n793), .Z(new_n854));
  OAI221_X1 g429(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n471), .C2(G118), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n485), .A2(G130), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n481), .A2(KEYINPUT103), .A3(G142), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT103), .B1(new_n481), .B2(G142), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n854), .B(new_n859), .Z(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n850), .A2(new_n860), .A3(new_n852), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(G160), .B(KEYINPUT102), .Z(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(new_n631), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n487), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n863), .A2(KEYINPUT104), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n850), .A2(new_n872), .A3(new_n860), .A4(new_n852), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n871), .A2(new_n862), .A3(new_n867), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n870), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  NAND4_X1  g451(.A1(new_n567), .A2(new_n597), .A3(new_n569), .A4(new_n601), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n601), .ZN(new_n879));
  OAI22_X1  g454(.A1(new_n609), .A2(new_n610), .B1(new_n879), .B2(new_n596), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT41), .B1(new_n878), .B2(new_n881), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n833), .A2(new_n832), .A3(new_n834), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT101), .B1(new_n838), .B2(new_n841), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n622), .B(new_n889), .ZN(new_n890));
  MUX2_X1   g465(.A(new_n882), .B(new_n886), .S(new_n890), .Z(new_n891));
  OR2_X1    g466(.A1(new_n891), .A2(KEYINPUT42), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(KEYINPUT42), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G290), .B(G305), .ZN(new_n895));
  XNOR2_X1  g470(.A(G303), .B(new_n782), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n892), .A2(new_n897), .A3(new_n893), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(G868), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n826), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT105), .B1(new_n902), .B2(G868), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n904), .B1(new_n905), .B2(new_n901), .ZN(G295));
  OAI21_X1  g481(.A(new_n904), .B1(new_n905), .B2(new_n901), .ZN(G331));
  NAND4_X1  g482(.A1(new_n537), .A2(G286), .A3(new_n538), .A4(new_n539), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(G301), .B2(G168), .ZN(new_n911));
  AOI211_X1 g486(.A(KEYINPUT106), .B(G286), .C1(new_n572), .C2(new_n573), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n843), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(G301), .A2(new_n909), .A3(G168), .ZN(new_n914));
  AOI21_X1  g489(.A(G286), .B1(new_n572), .B2(new_n573), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n889), .B(new_n914), .C1(new_n915), .C2(new_n910), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n913), .A2(new_n916), .A3(new_n882), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n885), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n877), .A2(new_n880), .A3(KEYINPUT108), .A4(new_n884), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n919), .A2(new_n883), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n913), .B2(new_n916), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n897), .B1(new_n917), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT109), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n925), .B(new_n897), .C1(new_n917), .C2(new_n922), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n913), .A2(new_n916), .A3(KEYINPUT107), .A4(new_n882), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n913), .A2(new_n916), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n931), .B2(new_n886), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n898), .B(new_n929), .C1(new_n932), .C2(new_n917), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n927), .A2(new_n928), .A3(new_n870), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n870), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n913), .A2(new_n916), .A3(new_n882), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n913), .A2(new_n916), .B1(new_n885), .B2(new_n883), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(new_n930), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n898), .B1(new_n938), .B2(new_n929), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n934), .A2(new_n940), .A3(KEYINPUT110), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  INV_X1    g517(.A(new_n935), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n928), .A4(new_n927), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n941), .A2(KEYINPUT111), .A3(new_n942), .A4(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OR3_X1    g525(.A1(new_n935), .A2(KEYINPUT43), .A3(new_n939), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n935), .B1(new_n924), .B2(new_n926), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n951), .B(KEYINPUT44), .C1(new_n928), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(G397));
  INV_X1    g529(.A(KEYINPUT120), .ZN(new_n955));
  XNOR2_X1  g530(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  XOR2_X1   g532(.A(KEYINPUT58), .B(G1341), .Z(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n492), .B2(new_n495), .ZN(new_n960));
  NAND2_X1  g535(.A1(G160), .A2(G40), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT118), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n961), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(G1996), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n957), .B1(new_n969), .B2(new_n550), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n550), .A3(new_n957), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT61), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n967), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1956), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(G299), .B(KEYINPUT57), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT56), .B(G2072), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n964), .A2(new_n966), .A3(new_n967), .A4(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n981), .B1(new_n979), .B2(new_n983), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n974), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n986), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(KEYINPUT61), .A3(new_n984), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n955), .B1(new_n973), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n972), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(new_n970), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(KEYINPUT120), .A3(new_n987), .A4(new_n989), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n960), .A2(new_n961), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n755), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n975), .A2(new_n967), .A3(new_n976), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n997), .B2(G1348), .ZN(new_n998));
  OR3_X1    g573(.A1(new_n998), .A2(KEYINPUT60), .A3(new_n602), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n998), .A2(new_n614), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n998), .A2(new_n614), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT60), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n991), .A2(new_n994), .A3(new_n999), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n984), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n988), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n968), .A2(new_n724), .ZN(new_n1007));
  INV_X1    g582(.A(G2084), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n975), .A2(new_n1008), .A3(new_n967), .A4(new_n976), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G168), .A2(new_n1006), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT51), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT121), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1014), .B(KEYINPUT51), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT122), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n1010), .A2(new_n1016), .B1(new_n1006), .B2(G168), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1013), .B(new_n1015), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n1011), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n997), .A2(G1961), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n968), .B2(G2078), .ZN(new_n1026));
  OR3_X1    g601(.A1(new_n968), .A2(new_n1025), .A3(G2078), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G171), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1024), .A2(G301), .A3(new_n1027), .A4(new_n1026), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1030), .A2(KEYINPUT54), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1021), .A2(new_n1023), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT124), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G303), .A2(G8), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT55), .ZN(new_n1035));
  INV_X1    g610(.A(G2090), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n997), .A2(new_n1036), .B1(new_n968), .B2(new_n775), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1037), .B2(new_n1006), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n968), .A2(new_n775), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(G2090), .B2(new_n977), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1035), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(G8), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n995), .A2(new_n1006), .ZN(new_n1043));
  XNOR2_X1  g618(.A(G305), .B(KEYINPUT49), .ZN(new_n1044));
  INV_X1    g619(.A(G1981), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n581), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1043), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n782), .A2(G1976), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1043), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1052), .B(G8), .C1(new_n960), .C2(new_n961), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT52), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1051), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1038), .A2(new_n1042), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1028), .A2(new_n605), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1030), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1032), .A2(new_n1033), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1033), .B1(new_n1032), .B2(new_n1063), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1005), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1058), .A2(G8), .A3(new_n1041), .A4(new_n1040), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1051), .A2(new_n1053), .A3(new_n782), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G305), .A2(G1981), .ZN(new_n1069));
  XOR2_X1   g644(.A(new_n1069), .B(KEYINPUT115), .Z(new_n1070));
  OAI21_X1  g645(.A(new_n1043), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n1006), .B(G286), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1038), .A2(new_n1042), .A3(new_n1072), .A4(new_n1058), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1073), .A2(KEYINPUT116), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1073), .B2(KEYINPUT116), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1067), .B(new_n1071), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(KEYINPUT117), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1059), .B1(new_n1079), .B2(KEYINPUT62), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1060), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1080), .B(new_n1081), .C1(KEYINPUT62), .C2(new_n1079), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1066), .A2(new_n1078), .A3(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n966), .A2(new_n961), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n712), .A2(new_n1084), .A3(G1996), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT112), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n752), .B(G2067), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n847), .B2(G1996), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1086), .B1(new_n1088), .B2(new_n1084), .ZN(new_n1089));
  XOR2_X1   g664(.A(new_n1089), .B(KEYINPUT113), .Z(new_n1090));
  INV_X1    g665(.A(new_n1084), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n793), .B(new_n796), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(G290), .B(G1986), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1084), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1083), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1090), .A2(new_n796), .A3(new_n791), .A4(new_n792), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n752), .A2(new_n755), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1091), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1091), .A2(G1986), .A3(G290), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(KEYINPUT125), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT48), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1093), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n712), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1091), .B1(new_n1104), .B2(new_n1087), .ZN(new_n1105));
  OR3_X1    g680(.A1(new_n1091), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT46), .B1(new_n1091), .B2(G1996), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT47), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1099), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1096), .A2(new_n1110), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g686(.A1(new_n655), .A2(G319), .A3(new_n668), .ZN(new_n1113));
  OR2_X1    g687(.A1(new_n1113), .A2(KEYINPUT126), .ZN(new_n1114));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT126), .ZN(new_n1115));
  AOI21_X1  g689(.A(G229), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g690(.A1(new_n941), .A2(new_n875), .A3(new_n945), .A4(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g691(.A(new_n1117), .B(KEYINPUT127), .ZN(G308));
  INV_X1    g692(.A(KEYINPUT127), .ZN(new_n1119));
  XNOR2_X1  g693(.A(new_n1117), .B(new_n1119), .ZN(G225));
endmodule


