//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n202), .B1(new_n205), .B2(KEYINPUT90), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(G1gat), .B2(new_n203), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI221_X1 g007(.A(new_n205), .B1(KEYINPUT90), .B2(new_n202), .C1(G1gat), .C2(new_n203), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT92), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT89), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n215), .A2(new_n216), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n213), .B(KEYINPUT14), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT89), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G43gat), .B(G50gat), .Z(new_n221));
  INV_X1    g020(.A(KEYINPUT15), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n218), .B1(new_n222), .B2(new_n221), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n220), .A2(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT93), .B1(new_n211), .B2(new_n226), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n231), .B(KEYINPUT13), .Z(new_n232));
  NAND3_X1  g031(.A1(new_n212), .A2(KEYINPUT93), .A3(new_n227), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n210), .B(KEYINPUT91), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n226), .A2(KEYINPUT17), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n226), .A2(KEYINPUT17), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n228), .A2(new_n231), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n228), .A2(KEYINPUT18), .A3(new_n238), .A4(new_n231), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n234), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(G169gat), .B(G197gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(new_n249), .Z(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n250), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n234), .A2(new_n241), .A3(new_n252), .A4(new_n242), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G78gat), .B(G106gat), .Z(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT81), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT31), .B(G50gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n257), .B(new_n258), .Z(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G141gat), .B(G148gat), .Z(new_n261));
  NAND2_X1  g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT2), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT76), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT76), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n262), .A2(new_n265), .A3(KEYINPUT2), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n261), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  OR3_X1    g066(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n268), .A2(new_n269), .B1(G155gat), .B2(G162gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  OR2_X1    g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n262), .B1(new_n272), .B2(KEYINPUT2), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n261), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n276));
  INV_X1    g075(.A(G211gat), .ZN(new_n277));
  INV_X1    g076(.A(G218gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT72), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G218gat), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n276), .B1(new_n282), .B2(KEYINPUT22), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT22), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT72), .B(G218gat), .ZN(new_n285));
  OAI211_X1 g084(.A(KEYINPUT73), .B(new_n284), .C1(new_n285), .C2(new_n277), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G197gat), .B(G204gat), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G211gat), .B(G218gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(new_n289), .A3(new_n291), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT29), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n275), .B1(new_n295), .B2(KEYINPUT3), .ZN(new_n296));
  INV_X1    g095(.A(G22gat), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n291), .B1(new_n287), .B2(new_n289), .ZN(new_n298));
  AOI211_X1 g097(.A(new_n288), .B(new_n292), .C1(new_n283), .C2(new_n286), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n267), .A2(new_n270), .B1(new_n261), .B2(new_n273), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n296), .A2(new_n297), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n304), .B1(new_n298), .B2(new_n299), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n301), .B1(new_n308), .B2(new_n302), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n305), .A2(new_n294), .A3(new_n293), .ZN(new_n310));
  OAI21_X1  g109(.A(G22gat), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G228gat), .A2(G233gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n307), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n307), .B2(new_n311), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n260), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT82), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT82), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n318), .B(new_n260), .C1(new_n314), .C2(new_n315), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n297), .B1(new_n296), .B2(new_n306), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n309), .A2(new_n310), .A3(G22gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n312), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n311), .A3(new_n313), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n259), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT83), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT83), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n323), .A2(new_n324), .A3(new_n327), .A4(new_n259), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT69), .ZN(new_n331));
  INV_X1    g130(.A(G169gat), .ZN(new_n332));
  INV_X1    g131(.A(G176gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT23), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(G169gat), .B2(G176gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n334), .B(new_n336), .C1(new_n332), .C2(new_n333), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT25), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT65), .ZN(new_n340));
  INV_X1    g139(.A(G183gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G190gat), .ZN(new_n342));
  INV_X1    g141(.A(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G183gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT24), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(G183gat), .A3(G190gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n340), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n342), .B2(new_n344), .ZN(new_n350));
  INV_X1    g149(.A(new_n348), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n350), .A2(KEYINPUT65), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n339), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G183gat), .B(G190gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n348), .B1(new_n354), .B2(new_n347), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n338), .B1(new_n355), .B2(new_n337), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT64), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT64), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n358), .B(new_n338), .C1(new_n355), .C2(new_n337), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n332), .A2(new_n333), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT26), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(G169gat), .B2(G176gat), .ZN(new_n364));
  OAI22_X1  g163(.A1(new_n361), .A2(new_n362), .B1(new_n341), .B2(new_n343), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n341), .A2(KEYINPUT27), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G183gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n369), .A3(new_n343), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT66), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT28), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT66), .A4(new_n343), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n372), .A2(KEYINPUT67), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n367), .A2(new_n369), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(KEYINPUT28), .A3(new_n343), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT28), .B1(new_n370), .B2(new_n371), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT67), .B1(new_n379), .B2(new_n374), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n366), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G113gat), .B(G120gat), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT68), .B(G127gat), .C1(new_n382), .C2(KEYINPUT1), .ZN(new_n383));
  INV_X1    g182(.A(G120gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G113gat), .ZN(new_n385));
  INV_X1    g184(.A(G113gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G120gat), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT1), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G127gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G134gat), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n383), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n383), .B2(new_n390), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n360), .A2(new_n381), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n394), .B1(new_n360), .B2(new_n381), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G227gat), .ZN(new_n398));
  INV_X1    g197(.A(G233gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n331), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n360), .A2(new_n381), .ZN(new_n402));
  NAND2_X1  g201(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n388), .A2(new_n403), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n382), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n405));
  OAI21_X1  g204(.A(G134gat), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n383), .A2(new_n390), .A3(new_n391), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n360), .A2(new_n381), .A3(new_n394), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n409), .A2(new_n331), .A3(new_n400), .A4(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT32), .B1(new_n401), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n400), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(new_n395), .B2(new_n396), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT34), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT34), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n417), .B(new_n414), .C1(new_n395), .C2(new_n396), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(G71gat), .B(G99gat), .Z(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT71), .ZN(new_n422));
  XNOR2_X1  g221(.A(G15gat), .B(G43gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT70), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n422), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n400), .A3(new_n410), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT69), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n411), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT32), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n428), .B2(new_n411), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n420), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n431), .B1(new_n420), .B2(new_n435), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G8gat), .B(G36gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(G64gat), .B(G92gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(G226gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(new_n399), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n360), .A2(new_n381), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n444), .A2(KEYINPUT29), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n360), .B2(new_n381), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n446), .A2(new_n448), .A3(new_n300), .ZN(new_n449));
  INV_X1    g248(.A(new_n300), .ZN(new_n450));
  INV_X1    g249(.A(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n402), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n360), .A2(new_n381), .A3(new_n445), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n442), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n300), .B1(new_n446), .B2(new_n448), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n355), .A2(KEYINPUT65), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n346), .A2(new_n340), .A3(new_n348), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n459), .A2(new_n339), .B1(new_n356), .B2(KEYINPUT64), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n377), .A3(new_n375), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n359), .A2(new_n460), .B1(new_n464), .B2(new_n366), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n450), .B(new_n453), .C1(new_n465), .C2(new_n447), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n456), .A2(new_n466), .A3(new_n441), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT30), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n467), .A2(KEYINPUT74), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT74), .B1(new_n467), .B2(new_n470), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n455), .B(new_n469), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n474));
  NAND2_X1  g273(.A1(G225gat), .A2(G233gat), .ZN(new_n475));
  INV_X1    g274(.A(new_n303), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n406), .B(new_n407), .C1(new_n301), .C2(new_n302), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n474), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(KEYINPUT4), .B(new_n301), .C1(new_n392), .C2(new_n393), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT4), .B1(new_n408), .B2(new_n301), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT78), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT78), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n301), .B1(new_n392), .B2(new_n393), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n484), .B1(new_n487), .B2(new_n480), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n479), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n394), .A2(new_n490), .A3(new_n303), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n491), .A2(new_n487), .A3(new_n480), .A4(new_n475), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n275), .A2(new_n406), .A3(new_n407), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n475), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n474), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(G1gat), .B(G29gat), .Z(new_n498));
  XNOR2_X1  g297(.A(G57gat), .B(G85gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  NAND3_X1  g301(.A1(new_n489), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT79), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n502), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n492), .A2(new_n496), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT78), .B1(new_n481), .B2(new_n482), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n484), .A3(new_n480), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n478), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n508), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n503), .A2(KEYINPUT79), .A3(new_n504), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n507), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT6), .B(new_n508), .C1(new_n509), .C2(new_n512), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT80), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n489), .A2(new_n497), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(new_n508), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n473), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n330), .A2(new_n438), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT35), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n330), .A2(new_n438), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT86), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n513), .A2(new_n503), .A3(new_n504), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n518), .A2(new_n527), .A3(new_n520), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n528), .B2(new_n473), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n455), .B1(new_n470), .B2(new_n467), .ZN(new_n530));
  INV_X1    g329(.A(new_n471), .ZN(new_n531));
  INV_X1    g330(.A(new_n472), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n527), .A3(new_n520), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT86), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  OAI22_X1  g335(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT37), .B1(new_n449), .B2(new_n454), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(KEYINPUT85), .A3(new_n442), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT85), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n456), .B2(new_n466), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n542), .B2(new_n441), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n456), .A2(new_n466), .A3(new_n541), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT38), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT38), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n542), .A2(new_n441), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n468), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n528), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n513), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n491), .B1(new_n483), .B2(new_n488), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT39), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n495), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n494), .A2(new_n495), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(new_n554), .ZN(new_n557));
  INV_X1    g356(.A(new_n491), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(new_n510), .B2(new_n511), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n557), .B1(new_n559), .B2(new_n475), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n555), .A2(new_n560), .A3(new_n502), .ZN(new_n561));
  NOR2_X1   g360(.A1(KEYINPUT84), .A2(KEYINPUT40), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n552), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n473), .B(new_n563), .C1(new_n562), .C2(new_n561), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n330), .A2(new_n551), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n436), .B2(new_n437), .ZN(new_n567));
  INV_X1    g366(.A(new_n431), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n413), .A2(new_n419), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n433), .A2(new_n434), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n420), .A2(new_n431), .A3(new_n435), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(KEYINPUT36), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n317), .A2(new_n319), .B1(new_n326), .B2(new_n328), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n518), .A2(new_n520), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n552), .B1(new_n505), .B2(new_n506), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(new_n514), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n575), .B1(new_n578), .B2(new_n473), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n565), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n255), .B1(new_n537), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n583));
  INV_X1    g382(.A(G64gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(KEYINPUT97), .A2(G57gat), .A3(G64gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n587), .A2(G71gat), .A3(G78gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n585), .B(new_n586), .C1(new_n588), .C2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(KEYINPUT95), .B(G57gat), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(G64gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT95), .B(G57gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n584), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n589), .A2(new_n587), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n590), .A2(KEYINPUT94), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n590), .A2(KEYINPUT94), .ZN(new_n599));
  NOR2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n597), .A2(KEYINPUT96), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT96), .B1(new_n597), .B2(new_n601), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n591), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n211), .B1(new_n582), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n605), .B(KEYINPUT98), .Z(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  INV_X1    g406(.A(G155gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n604), .A2(new_n582), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(new_n389), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G183gat), .B(G211gat), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n389), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n618), .B1(new_n616), .B2(new_n619), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n611), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n620), .A3(new_n610), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(G85gat), .A3(G92gat), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT7), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g437(.A1(G99gat), .A2(G106gat), .ZN(new_n639));
  INV_X1    g438(.A(G85gat), .ZN(new_n640));
  INV_X1    g439(.A(G92gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(KEYINPUT8), .A2(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n637), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G99gat), .B(G106gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n633), .B1(new_n226), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n236), .A2(new_n237), .A3(new_n645), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT99), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n648), .B2(new_n649), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n630), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n648), .A2(new_n649), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n651), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n653), .A3(new_n629), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n604), .A2(new_n645), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT10), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n643), .A2(new_n644), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n643), .A2(new_n644), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n665), .B(new_n591), .C1(new_n603), .C2(new_n602), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n604), .A2(new_n662), .A3(new_n645), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(G230gat), .A2(G233gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(KEYINPUT102), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n661), .A2(new_n666), .ZN(new_n676));
  INV_X1    g475(.A(new_n670), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(G120gat), .B(G148gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(G176gat), .B(G204gat), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n680), .B(new_n681), .Z(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n671), .A2(new_n678), .A3(new_n682), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n626), .A2(new_n660), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n581), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT103), .Z(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n578), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT104), .B(G1gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1324gat));
  XOR2_X1   g491(.A(KEYINPUT16), .B(G8gat), .Z(new_n693));
  AND3_X1   g492(.A1(new_n689), .A2(new_n473), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n202), .B1(new_n689), .B2(new_n473), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT42), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n689), .A2(new_n473), .A3(new_n693), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(G1325gat));
  INV_X1    g499(.A(G15gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n689), .A2(new_n701), .A3(new_n438), .ZN(new_n702));
  INV_X1    g501(.A(new_n574), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n689), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n704), .B2(new_n701), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n575), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(new_n685), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n679), .B2(new_n683), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n626), .A2(new_n660), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT105), .Z(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n581), .ZN(new_n713));
  INV_X1    g512(.A(new_n578), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n713), .A2(G29gat), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT45), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n571), .A2(new_n572), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n575), .A2(new_n717), .A3(KEYINPUT35), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n529), .A2(new_n535), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n330), .A2(new_n438), .A3(new_n522), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n718), .A2(new_n719), .B1(new_n720), .B2(KEYINPUT35), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n565), .A2(new_n574), .A3(new_n579), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n660), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT44), .B(new_n660), .C1(new_n721), .C2(new_n722), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n626), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(new_n255), .A3(new_n686), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n714), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n731), .ZN(G1328gat));
  NOR3_X1   g531(.A1(new_n713), .A2(G36gat), .A3(new_n533), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n730), .B2(new_n533), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1329gat));
  NOR2_X1   g535(.A1(new_n713), .A2(new_n717), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n703), .A2(G43gat), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n737), .A2(G43gat), .B1(new_n730), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g539(.A1(new_n727), .A2(new_n575), .A3(new_n729), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G50gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n330), .A2(G50gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n712), .A2(new_n581), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT48), .B1(new_n745), .B2(KEYINPUT106), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n747), .B(new_n748), .C1(new_n742), .C2(new_n744), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n746), .A2(new_n749), .ZN(G1331gat));
  NOR3_X1   g549(.A1(new_n626), .A2(new_n254), .A3(new_n660), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n686), .C1(new_n721), .C2(new_n722), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n714), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g553(.A(new_n752), .B(KEYINPUT107), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n473), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT49), .B(G64gat), .Z(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(G1333gat));
  NAND3_X1  g558(.A1(new_n755), .A2(G71gat), .A3(new_n703), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n752), .A2(new_n717), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(G71gat), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g562(.A1(new_n755), .A2(new_n575), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g564(.A(new_n254), .B1(new_n623), .B2(new_n625), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n766), .A2(new_n686), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n727), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768), .B2(new_n714), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n660), .B(new_n766), .C1(new_n721), .C2(new_n722), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT51), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n686), .A2(new_n578), .A3(new_n640), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(G1336gat));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n725), .A2(new_n473), .A3(new_n767), .A4(new_n726), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G92gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n771), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n710), .A2(G92gat), .A3(new_n533), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n774), .B(new_n776), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n779), .B(KEYINPUT108), .Z(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n785));
  INV_X1    g584(.A(new_n660), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n537), .B2(new_n580), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n787), .B2(new_n766), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n770), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n784), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n791), .A2(KEYINPUT110), .B1(G92gat), .B2(new_n775), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n784), .C1(new_n788), .C2(new_n790), .ZN(new_n794));
  AOI211_X1 g593(.A(new_n783), .B(new_n774), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(KEYINPUT110), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n794), .A3(new_n776), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT111), .B1(new_n797), .B2(KEYINPUT52), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n782), .B1(new_n795), .B2(new_n798), .ZN(G1337gat));
  OAI21_X1  g598(.A(G99gat), .B1(new_n768), .B2(new_n574), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n717), .A2(G99gat), .A3(new_n710), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n771), .B2(new_n801), .ZN(G1338gat));
  NAND4_X1  g601(.A1(new_n725), .A2(new_n575), .A3(new_n767), .A4(new_n726), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G106gat), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n330), .A2(G106gat), .A3(new_n710), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n804), .B(new_n805), .C1(new_n771), .C2(new_n806), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n803), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n788), .A2(new_n790), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n806), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT113), .B1(new_n803), .B2(G106gat), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n807), .B1(new_n812), .B2(new_n805), .ZN(G1339gat));
  NOR4_X1   g612(.A1(new_n626), .A2(new_n254), .A3(new_n660), .A4(new_n686), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n673), .A2(new_n816), .A3(new_n674), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n669), .B2(new_n670), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n667), .A2(new_n668), .A3(new_n677), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n682), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n660), .A2(new_n685), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n232), .B1(new_n230), .B2(new_n233), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n231), .B1(new_n228), .B2(new_n238), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n248), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n253), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n817), .A2(new_n820), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT114), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n831), .B(KEYINPUT55), .C1(new_n817), .C2(new_n820), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n822), .B(new_n827), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n830), .A2(new_n832), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n836), .A2(KEYINPUT115), .A3(new_n827), .A4(new_n822), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n686), .A2(KEYINPUT116), .A3(new_n827), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n710), .B2(new_n826), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n830), .A2(new_n832), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n254), .A2(new_n685), .A3(new_n821), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n838), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n835), .A2(new_n837), .B1(new_n843), .B2(new_n786), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n815), .B1(new_n844), .B2(new_n728), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n575), .A2(new_n717), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n714), .A2(new_n473), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n254), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n849), .A2(new_n850), .A3(G113gat), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n849), .B2(G113gat), .ZN(new_n852));
  OAI22_X1  g651(.A1(new_n851), .A2(new_n852), .B1(G113gat), .B2(new_n849), .ZN(G1340gat));
  NAND2_X1  g652(.A1(new_n847), .A2(new_n848), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n710), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(new_n384), .ZN(G1341gat));
  NOR2_X1   g655(.A1(new_n854), .A2(new_n626), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(new_n389), .ZN(G1342gat));
  NAND2_X1  g657(.A1(new_n847), .A2(new_n578), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n533), .A2(new_n660), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  XOR2_X1   g660(.A(KEYINPUT68), .B(G134gat), .Z(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT56), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n859), .B2(new_n860), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n859), .A2(KEYINPUT56), .A3(new_n863), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR4_X1   g667(.A1(new_n859), .A2(KEYINPUT118), .A3(KEYINPUT56), .A4(new_n863), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n864), .B(new_n865), .C1(new_n868), .C2(new_n869), .ZN(G1343gat));
  NAND2_X1  g669(.A1(new_n835), .A2(new_n837), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT55), .B1(new_n817), .B2(new_n820), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n842), .A2(new_n872), .B1(new_n710), .B2(new_n826), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n786), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n814), .B1(new_n875), .B2(new_n626), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT57), .B1(new_n876), .B2(new_n330), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n845), .A2(new_n878), .A3(new_n575), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n574), .A2(new_n578), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n473), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n877), .A2(new_n254), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n882), .A2(G141gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n843), .A2(new_n786), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n728), .B1(new_n871), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n814), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n330), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n881), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n255), .A2(G141gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT58), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n882), .A2(G141gat), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n892), .B(new_n893), .C1(new_n888), .C2(new_n889), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(G1344gat));
  OR2_X1    g694(.A1(new_n710), .A2(G148gat), .ZN(new_n896));
  OR3_X1    g695(.A1(new_n888), .A2(KEYINPUT119), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT119), .B1(new_n888), .B2(new_n896), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT57), .B1(new_n886), .B2(new_n330), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n822), .B1(new_n830), .B2(new_n832), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT120), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(KEYINPUT120), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n827), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n728), .B1(new_n905), .B2(new_n874), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n878), .B(new_n575), .C1(new_n906), .C2(new_n814), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n901), .A2(new_n686), .A3(new_n907), .A4(new_n881), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n900), .B1(new_n908), .B2(G148gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n877), .A2(new_n879), .A3(new_n881), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n710), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n900), .A2(G148gat), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n899), .B1(new_n909), .B2(new_n913), .ZN(G1345gat));
  OAI21_X1  g713(.A(G155gat), .B1(new_n910), .B2(new_n626), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n728), .A2(new_n608), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n888), .B2(new_n916), .ZN(G1346gat));
  OAI21_X1  g716(.A(G162gat), .B1(new_n910), .B2(new_n786), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n880), .A2(G162gat), .A3(new_n860), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n887), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1347gat));
  NAND2_X1  g720(.A1(new_n846), .A2(new_n473), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT121), .B1(new_n886), .B2(new_n578), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n845), .A2(new_n924), .A3(new_n714), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n922), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n255), .A2(G169gat), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n926), .A2(KEYINPUT122), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT122), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  INV_X1    g728(.A(new_n922), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n714), .B(new_n930), .C1(new_n885), .C2(new_n814), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n845), .A2(KEYINPUT123), .A3(new_n714), .A4(new_n930), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n254), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n935), .A2(new_n936), .A3(G169gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n935), .B2(G169gat), .ZN(new_n938));
  OAI22_X1  g737(.A1(new_n928), .A2(new_n929), .B1(new_n937), .B2(new_n938), .ZN(G1348gat));
  NAND3_X1  g738(.A1(new_n926), .A2(new_n333), .A3(new_n686), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n933), .A2(new_n686), .A3(new_n934), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n333), .B2(new_n941), .ZN(G1349gat));
  NAND3_X1  g741(.A1(new_n933), .A2(new_n728), .A3(new_n934), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(G183gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n923), .A2(new_n925), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n728), .A2(new_n376), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(new_n930), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT60), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n944), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1350gat));
  NAND3_X1  g751(.A1(new_n926), .A2(new_n343), .A3(new_n660), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n933), .A2(new_n660), .A3(new_n934), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n954), .A2(new_n955), .A3(G190gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n954), .B2(G190gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(G1351gat));
  NAND3_X1  g757(.A1(new_n574), .A2(new_n714), .A3(new_n473), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT125), .Z(new_n960));
  NAND3_X1  g759(.A1(new_n901), .A2(new_n907), .A3(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(G197gat), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n961), .A2(new_n962), .A3(new_n255), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n703), .A2(new_n533), .A3(new_n330), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n254), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n963), .B1(new_n962), .B2(new_n965), .ZN(G1352gat));
  NOR2_X1   g765(.A1(new_n710), .A2(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n945), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n945), .A2(new_n970), .A3(new_n964), .A4(new_n967), .ZN(new_n971));
  OAI21_X1  g770(.A(G204gat), .B1(new_n961), .B2(new_n710), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(G1353gat));
  NAND4_X1  g772(.A1(new_n945), .A2(new_n277), .A3(new_n728), .A4(new_n964), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n959), .A2(new_n626), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n901), .A2(new_n907), .A3(new_n975), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n961), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n786), .A2(new_n285), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT127), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n961), .A2(new_n980), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n945), .A2(new_n660), .A3(new_n964), .ZN(new_n986));
  AOI22_X1  g785(.A1(new_n984), .A2(new_n985), .B1(new_n278), .B2(new_n986), .ZN(G1355gat));
endmodule


