

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U324 ( .A(n397), .B(n396), .ZN(n535) );
  XOR2_X1 U325 ( .A(n360), .B(n359), .Z(n292) );
  XOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT123), .Z(n293) );
  INV_X1 U327 ( .A(KEYINPUT9), .ZN(n350) );
  XNOR2_X1 U328 ( .A(n351), .B(n350), .ZN(n352) );
  INV_X1 U329 ( .A(KEYINPUT116), .ZN(n395) );
  XNOR2_X1 U330 ( .A(n408), .B(n352), .ZN(n353) );
  XNOR2_X1 U331 ( .A(n395), .B(KEYINPUT48), .ZN(n396) );
  XNOR2_X1 U332 ( .A(n361), .B(n292), .ZN(n362) );
  XNOR2_X1 U333 ( .A(n363), .B(n362), .ZN(n560) );
  NOR2_X1 U334 ( .A1(n457), .A2(n539), .ZN(n565) );
  XOR2_X1 U335 ( .A(n456), .B(n455), .Z(n527) );
  XNOR2_X1 U336 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n459) );
  XNOR2_X1 U337 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XNOR2_X1 U338 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n294), .B(KEYINPUT88), .ZN(n295) );
  XOR2_X1 U340 ( .A(n295), .B(KEYINPUT19), .Z(n297) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(G183GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n446) );
  XOR2_X1 U343 ( .A(G8GAT), .B(KEYINPUT80), .Z(n366) );
  XOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .Z(n354) );
  XOR2_X1 U345 ( .A(n366), .B(n354), .Z(n299) );
  NAND2_X1 U346 ( .A1(G226GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U348 ( .A(KEYINPUT98), .B(G92GAT), .Z(n301) );
  XNOR2_X1 U349 ( .A(G218GAT), .B(G204GAT), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U351 ( .A(n303), .B(n302), .Z(n309) );
  XOR2_X1 U352 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n305) );
  XNOR2_X1 U353 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U355 ( .A(G197GAT), .B(n306), .Z(n413) );
  INV_X1 U356 ( .A(n413), .ZN(n307) );
  XOR2_X1 U357 ( .A(G176GAT), .B(G64GAT), .Z(n330) );
  XOR2_X1 U358 ( .A(n307), .B(n330), .Z(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n446), .B(n310), .ZN(n525) );
  XOR2_X1 U361 ( .A(G197GAT), .B(G22GAT), .Z(n312) );
  XNOR2_X1 U362 ( .A(G50GAT), .B(G36GAT), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U364 ( .A(n313), .B(G15GAT), .Z(n315) );
  XOR2_X1 U365 ( .A(G113GAT), .B(G1GAT), .Z(n427) );
  XNOR2_X1 U366 ( .A(G169GAT), .B(n427), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n321) );
  XOR2_X1 U368 ( .A(G29GAT), .B(G43GAT), .Z(n317) );
  XNOR2_X1 U369 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n358) );
  XOR2_X1 U371 ( .A(n358), .B(KEYINPUT67), .Z(n319) );
  NAND2_X1 U372 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(n321), .B(n320), .Z(n329) );
  XOR2_X1 U375 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n323) );
  XNOR2_X1 U376 ( .A(G141GAT), .B(KEYINPUT66), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U378 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n325) );
  XNOR2_X1 U379 ( .A(KEYINPUT65), .B(G8GAT), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U382 ( .A(n329), .B(n328), .Z(n510) );
  INV_X1 U383 ( .A(n510), .ZN(n571) );
  XOR2_X1 U384 ( .A(G120GAT), .B(G71GAT), .Z(n441) );
  XNOR2_X1 U385 ( .A(n441), .B(n330), .ZN(n345) );
  XOR2_X1 U386 ( .A(G85GAT), .B(G92GAT), .Z(n332) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G106GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n357) );
  XOR2_X1 U389 ( .A(n357), .B(KEYINPUT33), .Z(n334) );
  NAND2_X1 U390 ( .A1(G230GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U392 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n336) );
  XNOR2_X1 U393 ( .A(KEYINPUT32), .B(KEYINPUT71), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U395 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U396 ( .A(G78GAT), .B(G148GAT), .Z(n340) );
  XNOR2_X1 U397 ( .A(KEYINPUT72), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n407) );
  XNOR2_X1 U399 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n341), .B(KEYINPUT13), .ZN(n370) );
  XNOR2_X1 U401 ( .A(n407), .B(n370), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U403 ( .A(n345), .B(n344), .Z(n575) );
  XOR2_X1 U404 ( .A(n575), .B(KEYINPUT41), .Z(n554) );
  NAND2_X1 U405 ( .A1(n571), .A2(n554), .ZN(n347) );
  XOR2_X1 U406 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n384) );
  XOR2_X1 U408 ( .A(G162GAT), .B(KEYINPUT75), .Z(n349) );
  XNOR2_X1 U409 ( .A(G50GAT), .B(G218GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n408) );
  NAND2_X1 U411 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n353), .B(KEYINPUT77), .ZN(n356) );
  XOR2_X1 U413 ( .A(n354), .B(KEYINPUT76), .Z(n355) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n361) );
  XOR2_X1 U416 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n360) );
  XNOR2_X1 U417 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n359) );
  XOR2_X1 U418 ( .A(G78GAT), .B(G211GAT), .Z(n365) );
  XNOR2_X1 U419 ( .A(G183GAT), .B(G71GAT), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n367) );
  XOR2_X1 U421 ( .A(n367), .B(n366), .Z(n369) );
  XNOR2_X1 U422 ( .A(G1GAT), .B(G64GAT), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n371) );
  XOR2_X1 U424 ( .A(n371), .B(n370), .Z(n373) );
  XOR2_X1 U425 ( .A(G15GAT), .B(G127GAT), .Z(n450) );
  XOR2_X1 U426 ( .A(G22GAT), .B(G155GAT), .Z(n401) );
  XNOR2_X1 U427 ( .A(n450), .B(n401), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U429 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n375) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U432 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U433 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n379) );
  XNOR2_X1 U434 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n380), .B(KEYINPUT84), .ZN(n381) );
  XOR2_X1 U437 ( .A(n382), .B(n381), .Z(n465) );
  INV_X1 U438 ( .A(n465), .ZN(n579) );
  NOR2_X1 U439 ( .A1(n560), .A2(n579), .ZN(n383) );
  NAND2_X1 U440 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n385), .B(KEYINPUT47), .ZN(n394) );
  INV_X1 U442 ( .A(KEYINPUT79), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n386), .B(n560), .ZN(n458) );
  XNOR2_X1 U444 ( .A(KEYINPUT36), .B(n458), .ZN(n581) );
  NAND2_X1 U445 ( .A1(n581), .A2(n579), .ZN(n389) );
  XOR2_X1 U446 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n387) );
  XNOR2_X1 U447 ( .A(KEYINPUT64), .B(n387), .ZN(n388) );
  XOR2_X1 U448 ( .A(n389), .B(n388), .Z(n390) );
  NOR2_X1 U449 ( .A1(n575), .A2(n390), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n391), .B(KEYINPUT115), .ZN(n392) );
  NOR2_X1 U451 ( .A1(n392), .A2(n571), .ZN(n393) );
  NOR2_X1 U452 ( .A1(n394), .A2(n393), .ZN(n397) );
  NAND2_X1 U453 ( .A1(n525), .A2(n535), .ZN(n398) );
  XOR2_X1 U454 ( .A(n293), .B(n398), .Z(n568) );
  XOR2_X1 U455 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n400) );
  XNOR2_X1 U456 ( .A(G141GAT), .B(KEYINPUT93), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n426) );
  XOR2_X1 U458 ( .A(n426), .B(KEYINPUT23), .Z(n403) );
  XNOR2_X1 U459 ( .A(G106GAT), .B(n401), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n412) );
  XOR2_X1 U461 ( .A(KEYINPUT94), .B(KEYINPUT24), .Z(n405) );
  NAND2_X1 U462 ( .A1(G228GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U464 ( .A(n406), .B(KEYINPUT22), .Z(n410) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U468 ( .A(n414), .B(n413), .Z(n476) );
  XOR2_X1 U469 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n416) );
  XNOR2_X1 U470 ( .A(KEYINPUT5), .B(KEYINPUT95), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n435) );
  XOR2_X1 U472 ( .A(G85GAT), .B(G155GAT), .Z(n418) );
  XNOR2_X1 U473 ( .A(G120GAT), .B(G127GAT), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U475 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n420) );
  XNOR2_X1 U476 ( .A(G148GAT), .B(G57GAT), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U478 ( .A(n422), .B(n421), .Z(n433) );
  XNOR2_X1 U479 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n423), .B(KEYINPUT85), .ZN(n442) );
  XOR2_X1 U481 ( .A(KEYINPUT4), .B(n442), .Z(n425) );
  NAND2_X1 U482 ( .A1(G225GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n431) );
  XOR2_X1 U484 ( .A(n426), .B(G162GAT), .Z(n429) );
  XNOR2_X1 U485 ( .A(G29GAT), .B(n427), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n523) );
  INV_X1 U490 ( .A(n523), .ZN(n567) );
  AND2_X1 U491 ( .A1(n476), .A2(n567), .ZN(n436) );
  NAND2_X1 U492 ( .A1(n568), .A2(n436), .ZN(n438) );
  XOR2_X1 U493 ( .A(KEYINPUT55), .B(KEYINPUT124), .Z(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n457) );
  XOR2_X1 U495 ( .A(G176GAT), .B(KEYINPUT90), .Z(n440) );
  XNOR2_X1 U496 ( .A(G113GAT), .B(KEYINPUT89), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n456) );
  XOR2_X1 U498 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n454) );
  XOR2_X1 U502 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n448) );
  XNOR2_X1 U503 ( .A(G190GAT), .B(KEYINPUT87), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U505 ( .A(n449), .B(G99GAT), .Z(n452) );
  XNOR2_X1 U506 ( .A(G43GAT), .B(n450), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n455) );
  INV_X1 U509 ( .A(n527), .ZN(n539) );
  NAND2_X1 U510 ( .A1(n565), .A2(n458), .ZN(n460) );
  XOR2_X1 U511 ( .A(KEYINPUT109), .B(n554), .Z(n542) );
  NAND2_X1 U512 ( .A1(n565), .A2(n542), .ZN(n464) );
  XOR2_X1 U513 ( .A(G176GAT), .B(KEYINPUT57), .Z(n462) );
  XOR2_X1 U514 ( .A(KEYINPUT125), .B(KEYINPUT56), .Z(n461) );
  XNOR2_X1 U515 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n464), .B(n463), .ZN(G1349GAT) );
  NOR2_X1 U517 ( .A1(n458), .A2(n465), .ZN(n466) );
  XNOR2_X1 U518 ( .A(n466), .B(KEYINPUT16), .ZN(n482) );
  NAND2_X1 U519 ( .A1(n527), .A2(n525), .ZN(n467) );
  NAND2_X1 U520 ( .A1(n476), .A2(n467), .ZN(n468) );
  XNOR2_X1 U521 ( .A(KEYINPUT25), .B(n468), .ZN(n472) );
  XNOR2_X1 U522 ( .A(KEYINPUT27), .B(n525), .ZN(n474) );
  NOR2_X1 U523 ( .A1(n476), .A2(n527), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT26), .ZN(n569) );
  NAND2_X1 U525 ( .A1(n474), .A2(n569), .ZN(n470) );
  XNOR2_X1 U526 ( .A(KEYINPUT101), .B(n470), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n472), .A2(n471), .ZN(n473) );
  NOR2_X1 U528 ( .A1(n523), .A2(n473), .ZN(n480) );
  NAND2_X1 U529 ( .A1(n523), .A2(n474), .ZN(n475) );
  XNOR2_X1 U530 ( .A(n475), .B(KEYINPUT99), .ZN(n534) );
  XOR2_X1 U531 ( .A(KEYINPUT28), .B(n476), .Z(n531) );
  INV_X1 U532 ( .A(n531), .ZN(n537) );
  NAND2_X1 U533 ( .A1(n534), .A2(n537), .ZN(n477) );
  NOR2_X1 U534 ( .A1(n527), .A2(n477), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(KEYINPUT100), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n493) );
  INV_X1 U537 ( .A(n493), .ZN(n481) );
  NAND2_X1 U538 ( .A1(n482), .A2(n481), .ZN(n511) );
  OR2_X1 U539 ( .A1(n575), .A2(n510), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(KEYINPUT74), .ZN(n498) );
  NOR2_X1 U541 ( .A1(n511), .A2(n498), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n484), .B(KEYINPUT102), .ZN(n491) );
  NAND2_X1 U543 ( .A1(n491), .A2(n523), .ZN(n487) );
  XOR2_X1 U544 ( .A(G1GAT), .B(KEYINPUT103), .Z(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT34), .B(n485), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U547 ( .A1(n491), .A2(n525), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U550 ( .A1(n527), .A2(n491), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U552 ( .A1(n491), .A2(n531), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .Z(n501) );
  XOR2_X1 U555 ( .A(KEYINPUT37), .B(KEYINPUT106), .Z(n497) );
  NOR2_X1 U556 ( .A1(n579), .A2(n493), .ZN(n494) );
  XOR2_X1 U557 ( .A(KEYINPUT105), .B(n494), .Z(n495) );
  NAND2_X1 U558 ( .A1(n495), .A2(n581), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n522) );
  NOR2_X1 U560 ( .A1(n522), .A2(n498), .ZN(n499) );
  XNOR2_X1 U561 ( .A(KEYINPUT38), .B(n499), .ZN(n508) );
  NAND2_X1 U562 ( .A1(n508), .A2(n523), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(KEYINPUT104), .B(n502), .ZN(G1328GAT) );
  XOR2_X1 U565 ( .A(G36GAT), .B(KEYINPUT107), .Z(n504) );
  NAND2_X1 U566 ( .A1(n508), .A2(n525), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1329GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n506) );
  NAND2_X1 U569 ( .A1(n527), .A2(n508), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U571 ( .A(G43GAT), .B(n507), .Z(G1330GAT) );
  NAND2_X1 U572 ( .A1(n531), .A2(n508), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(n509), .ZN(G1331GAT) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n514) );
  NAND2_X1 U575 ( .A1(n510), .A2(n542), .ZN(n521) );
  NOR2_X1 U576 ( .A1(n511), .A2(n521), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT110), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n523), .A2(n518), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  XOR2_X1 U580 ( .A(G64GAT), .B(KEYINPUT111), .Z(n516) );
  NAND2_X1 U581 ( .A1(n518), .A2(n525), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n518), .A2(n527), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U586 ( .A1(n518), .A2(n531), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n530), .A2(n523), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n525), .A2(n530), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(KEYINPUT112), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n532), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(KEYINPUT118), .ZN(n541) );
  NAND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(KEYINPUT117), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n537), .A2(n551), .ZN(n538) );
  NOR2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n571), .A2(n548), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U607 ( .A1(n548), .A2(n542), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U609 ( .A(G120GAT), .B(n545), .Z(G1341GAT) );
  NAND2_X1 U610 ( .A1(n548), .A2(n579), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U614 ( .A1(n548), .A2(n458), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  AND2_X1 U616 ( .A1(n551), .A2(n569), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n571), .A2(n561), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT120), .B(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n556) );
  NAND2_X1 U621 ( .A1(n561), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT53), .Z(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n579), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n571), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n579), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n573) );
  AND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n570) );
  AND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n582) );
  NAND2_X1 U637 ( .A1(n582), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n582), .A2(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n584) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

