//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(G127gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n209));
  XNOR2_X1  g008(.A(G113gat), .B(G120gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n211));
  INV_X1    g010(.A(G134gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213));
  INV_X1    g012(.A(G113gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(G120gat), .ZN(new_n215));
  INV_X1    g014(.A(G120gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G113gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n213), .B(new_n208), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n211), .A2(new_n212), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n212), .B1(new_n211), .B2(new_n218), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT72), .A2(G148gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT72), .A2(G148gat), .ZN(new_n223));
  OAI21_X1  g022(.A(G141gat), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G141gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G148gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  INV_X1    g027(.A(G155gat), .ZN(new_n229));
  INV_X1    g028(.A(G162gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n224), .A2(new_n226), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n230), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n227), .ZN(new_n234));
  INV_X1    g033(.A(G148gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G141gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n226), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n234), .B1(new_n228), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT3), .B1(new_n232), .B2(new_n238), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n221), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n244), .B(new_n239), .C1(new_n219), .C2(new_n220), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n209), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n216), .A2(G113gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n214), .A2(G120gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n247), .B1(new_n250), .B2(new_n213), .ZN(new_n251));
  AOI211_X1 g050(.A(KEYINPUT1), .B(G127gat), .C1(new_n248), .C2(new_n249), .ZN(new_n252));
  OAI21_X1  g051(.A(G134gat), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n211), .A2(new_n212), .A3(new_n218), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n244), .B1(new_n255), .B2(new_n239), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n207), .B(new_n243), .C1(new_n246), .C2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT5), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n239), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(new_n253), .A3(new_n254), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n239), .B1(new_n219), .B2(new_n220), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n207), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(KEYINPUT4), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n242), .A2(new_n253), .A3(new_n254), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n264), .A2(new_n245), .B1(new_n265), .B2(new_n241), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n263), .B1(new_n266), .B2(new_n207), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n206), .B(new_n259), .C1(new_n267), .C2(new_n258), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT73), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n206), .ZN(new_n271));
  INV_X1    g070(.A(new_n263), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n258), .B1(new_n257), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT5), .B1(new_n266), .B2(new_n207), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n268), .A3(new_n269), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n273), .A2(new_n274), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT6), .A4(new_n206), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n270), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  AND2_X1   g080(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(KEYINPUT28), .B(new_n281), .C1(new_n282), .C2(new_n283), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR3_X1   g091(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296));
  NOR2_X1   g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  AND4_X1   g099(.A1(new_n296), .A2(new_n298), .A3(new_n300), .A4(new_n291), .ZN(new_n301));
  INV_X1    g100(.A(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n281), .ZN(new_n303));
  NAND3_X1  g102(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT24), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n288), .A2(new_n295), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT64), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n303), .B(new_n304), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n300), .A3(new_n291), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT25), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n309), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G226gat), .ZN(new_n319));
  INV_X1    g118(.A(G233gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT69), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT69), .ZN(new_n323));
  INV_X1    g122(.A(new_n321), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n307), .A2(KEYINPUT64), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n305), .A2(new_n325), .A3(new_n313), .ZN(new_n326));
  INV_X1    g125(.A(new_n316), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n296), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n294), .B1(new_n286), .B2(new_n287), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n307), .A2(new_n303), .A3(new_n304), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n330), .A2(new_n316), .A3(KEYINPUT25), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n323), .B(new_n324), .C1(new_n332), .C2(KEYINPUT29), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n324), .B1(new_n309), .B2(new_n317), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI211_X1 g135(.A(KEYINPUT70), .B(new_n324), .C1(new_n309), .C2(new_n317), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n322), .B(new_n333), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(G197gat), .A2(G204gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(G197gat), .A2(G204gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT22), .ZN(new_n341));
  NAND2_X1  g140(.A1(G211gat), .A2(G218gat), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n339), .A2(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(G211gat), .A2(G218gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n342), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n345), .B2(new_n342), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n349), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(new_n343), .A3(new_n347), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n288), .A2(new_n295), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n301), .A2(new_n308), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n317), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n321), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n359), .A2(new_n353), .A3(new_n334), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT71), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n338), .B2(new_n353), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n369), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n364), .A2(KEYINPUT30), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT30), .B1(new_n364), .B2(new_n371), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n280), .A2(new_n370), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT74), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n364), .A2(new_n365), .ZN(new_n377));
  AOI211_X1 g176(.A(KEYINPUT71), .B(new_n360), .C1(new_n338), .C2(new_n353), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n377), .A2(new_n378), .A3(new_n371), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n354), .A2(new_n361), .A3(new_n371), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n364), .A2(KEYINPUT30), .A3(new_n371), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT74), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n280), .ZN(new_n387));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT66), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n357), .A2(new_n221), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n255), .A2(new_n317), .A3(new_n309), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n357), .B2(new_n221), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT32), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT67), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT32), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT66), .B1(new_n332), .B2(new_n255), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n392), .A3(new_n391), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n400), .B2(new_n389), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT67), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n395), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n397), .A2(new_n403), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n401), .B1(new_n408), .B2(new_n407), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n399), .A2(new_n388), .A3(new_n392), .A4(new_n391), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n412), .B(KEYINPUT34), .Z(new_n413));
  AND3_X1   g212(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n410), .B2(new_n411), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n241), .A2(new_n358), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n353), .ZN(new_n417));
  AND2_X1   g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n350), .A2(new_n358), .A3(new_n352), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n419), .A2(new_n239), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n417), .A2(new_n242), .A3(new_n418), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(KEYINPUT76), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT76), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n350), .A2(new_n352), .A3(new_n423), .A4(new_n358), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n240), .A3(new_n424), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n425), .A2(new_n260), .B1(new_n353), .B2(new_n416), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n421), .B1(new_n426), .B2(new_n418), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT77), .B(G22gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n428), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n430), .B(new_n421), .C1(new_n426), .C2(new_n418), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT31), .B(G50gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n435), .B(KEYINPUT75), .Z(new_n436));
  AND2_X1   g235(.A1(new_n431), .A2(new_n435), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n427), .A2(G22gat), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n432), .A2(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n414), .A2(new_n415), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n376), .A2(new_n387), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT35), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT80), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n275), .A2(new_n269), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n273), .B2(new_n274), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT79), .B(new_n259), .C1(new_n267), .C2(new_n258), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n444), .B1(new_n206), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n270), .A2(new_n279), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n374), .A2(new_n370), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n443), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n271), .B1(new_n446), .B2(new_n447), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n279), .B(new_n270), .C1(new_n454), .C2(new_n444), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n385), .A2(KEYINPUT80), .A3(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(KEYINPUT81), .B(KEYINPUT35), .Z(new_n457));
  NAND4_X1  g256(.A1(new_n453), .A2(new_n440), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n377), .A2(new_n378), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n371), .B1(new_n364), .B2(new_n459), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT38), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n353), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n338), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n359), .A2(new_n334), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n459), .B1(new_n466), .B2(new_n353), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT38), .B(new_n371), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n364), .A2(new_n459), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n468), .A2(new_n469), .B1(new_n364), .B2(new_n371), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT40), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n261), .A2(KEYINPUT78), .A3(new_n207), .A4(new_n262), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT39), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT78), .B1(new_n266), .B2(new_n207), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n261), .A2(new_n207), .A3(new_n262), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n243), .B1(new_n246), .B2(new_n256), .ZN(new_n478));
  INV_X1    g277(.A(new_n207), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n271), .B1(new_n480), .B2(KEYINPUT39), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n472), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n474), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT78), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n478), .B2(new_n479), .ZN(new_n485));
  INV_X1    g284(.A(new_n476), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n266), .A2(new_n207), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT39), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n206), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(KEYINPUT40), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(new_n454), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n439), .B1(new_n452), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n410), .A2(new_n411), .ZN(new_n495));
  INV_X1    g294(.A(new_n413), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(KEYINPUT36), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n414), .B2(new_n415), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n471), .A2(new_n494), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n386), .B1(new_n385), .B2(new_n280), .ZN(new_n503));
  AND4_X1   g302(.A1(new_n386), .A2(new_n280), .A3(new_n370), .A4(new_n374), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n439), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n442), .A2(new_n458), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G183gat), .B(G211gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n507), .B(new_n508), .Z(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT9), .ZN(new_n512));
  NAND2_X1  g311(.A1(G71gat), .A2(G78gat), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G71gat), .B(G78gat), .Z(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n516), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(new_n208), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G155gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G231gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(new_n320), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT16), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G1gat), .B2(new_n527), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n531), .A2(G8gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(G8gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(KEYINPUT84), .A3(new_n533), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n519), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT90), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n541), .A2(KEYINPUT90), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT89), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n544), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT89), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n547), .A3(new_n542), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n526), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n548), .A3(new_n526), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n524), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  NOR3_X1   g352(.A1(new_n553), .A2(new_n549), .A3(new_n523), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n510), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT7), .ZN(new_n556));
  INV_X1    g355(.A(G92gat), .ZN(new_n557));
  OAI211_X1 g356(.A(KEYINPUT91), .B(new_n556), .C1(new_n203), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n203), .A2(new_n557), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n560));
  OAI211_X1 g359(.A(G85gat), .B(G92gat), .C1(new_n560), .C2(KEYINPUT7), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n556), .A2(KEYINPUT91), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n558), .B(new_n559), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(KEYINPUT92), .A2(G99gat), .A3(G106gat), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n566), .A2(KEYINPUT8), .A3(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G99gat), .B(G106gat), .Z(new_n569));
  OR3_X1    g368(.A1(new_n563), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n563), .B2(new_n568), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT93), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT14), .ZN(new_n574));
  INV_X1    g373(.A(G29gat), .ZN(new_n575));
  INV_X1    g374(.A(G36gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n577), .A2(new_n578), .B1(G29gat), .B2(G36gat), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n580));
  XNOR2_X1  g379(.A(G43gat), .B(G50gat), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n573), .B1(KEYINPUT17), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n585), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT83), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT83), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n586), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n573), .A2(new_n587), .B1(KEYINPUT41), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G134gat), .B(G162gat), .Z(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n594), .A2(KEYINPUT41), .ZN(new_n599));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n596), .A2(new_n597), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n598), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n550), .A2(new_n551), .A3(new_n524), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n523), .B1(new_n553), .B2(new_n549), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n608), .A3(new_n509), .ZN(new_n609));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT95), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n572), .A2(KEYINPUT94), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n519), .B1(new_n572), .B2(KEYINPUT94), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT10), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n573), .A2(KEYINPUT10), .A3(new_n539), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n612), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n616), .A2(new_n611), .A3(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n555), .A2(new_n606), .A3(new_n609), .A4(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n534), .B1(new_n585), .B2(KEYINPUT17), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n592), .B2(new_n589), .ZN(new_n634));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n587), .A2(new_n536), .A3(new_n537), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT18), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n634), .A2(KEYINPUT18), .A3(new_n635), .A4(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n538), .A2(new_n585), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n636), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n635), .B(KEYINPUT13), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT86), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n643), .A2(KEYINPUT86), .A3(new_n644), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n641), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n641), .A2(new_n647), .A3(KEYINPUT85), .A4(new_n648), .ZN(new_n651));
  XNOR2_X1  g450(.A(G113gat), .B(G141gat), .ZN(new_n652));
  INV_X1    g451(.A(G197gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT11), .B(G169gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT12), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n651), .B(new_n658), .C1(new_n640), .C2(new_n649), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT87), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n660), .A2(KEYINPUT87), .A3(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n506), .A2(new_n632), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n280), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n452), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n671), .A2(G8gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT16), .B(G8gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT42), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(KEYINPUT42), .B2(new_n674), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT96), .ZN(G1325gat));
  NOR2_X1   g476(.A1(new_n414), .A2(new_n415), .ZN(new_n678));
  AOI21_X1  g477(.A(G15gat), .B1(new_n667), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n501), .A2(new_n499), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n679), .B1(new_n667), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n439), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  NOR2_X1   g485(.A1(new_n506), .A2(new_n606), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n687), .A2(KEYINPUT97), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(KEYINPUT44), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(KEYINPUT44), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n555), .A2(new_n609), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n631), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n660), .A2(new_n661), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G29gat), .B1(new_n696), .B2(new_n280), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n693), .A2(new_n666), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n687), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n699), .A2(G29gat), .A3(new_n280), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT45), .Z(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n699), .A2(G36gat), .A3(new_n385), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT98), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n704), .B2(new_n703), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n452), .A3(new_n695), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT99), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n708), .B2(new_n709), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(G1329gat));
  INV_X1    g511(.A(new_n678), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n699), .A2(G43gat), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n689), .A2(new_n681), .A3(new_n690), .A4(new_n695), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G43gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT47), .B(new_n714), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(G43gat), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n720), .A2(new_n714), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(KEYINPUT47), .B2(new_n721), .ZN(G1330gat));
  INV_X1    g521(.A(new_n439), .ZN(new_n723));
  OAI21_X1  g522(.A(G50gat), .B1(new_n696), .B2(new_n723), .ZN(new_n724));
  OR3_X1    g523(.A1(new_n699), .A2(G50gat), .A3(new_n723), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n724), .A2(KEYINPUT48), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1331gat));
  INV_X1    g529(.A(new_n692), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n606), .A3(new_n630), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(new_n506), .A3(new_n662), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n668), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT102), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT101), .B(G57gat), .Z(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1332gat));
  NAND2_X1  g536(.A1(new_n733), .A2(new_n452), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT49), .B(G64gat), .Z(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n738), .B2(new_n740), .ZN(G1333gat));
  NAND3_X1  g540(.A1(new_n733), .A2(G71gat), .A3(new_n681), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n678), .B(KEYINPUT103), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n733), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n744), .B2(G71gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g545(.A1(new_n733), .A2(new_n439), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g547(.A1(new_n731), .A2(new_n631), .A3(new_n662), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n691), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n280), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n506), .B2(new_n606), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n731), .A2(new_n662), .ZN(new_n754));
  INV_X1    g553(.A(new_n606), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n456), .A2(new_n440), .A3(new_n457), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n756), .A2(new_n453), .B1(new_n441), .B2(KEYINPUT35), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT38), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n363), .A2(KEYINPUT37), .A3(new_n366), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n461), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n468), .A2(new_n469), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n380), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n760), .A2(new_n455), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n448), .A2(new_n206), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(new_n491), .A3(new_n482), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n723), .B1(new_n385), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n680), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n723), .B1(new_n376), .B2(new_n387), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(KEYINPUT104), .B(new_n755), .C1(new_n757), .C2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n753), .A2(new_n770), .A3(KEYINPUT51), .A4(new_n754), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(KEYINPUT105), .A3(new_n774), .ZN(new_n775));
  OR3_X1    g574(.A1(new_n771), .A2(KEYINPUT105), .A3(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT106), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n280), .A2(G85gat), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n778), .A2(new_n630), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n751), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n751), .A2(new_n782), .A3(KEYINPUT107), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1336gat));
  NAND4_X1  g586(.A1(new_n689), .A2(new_n452), .A3(new_n690), .A4(new_n749), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G92gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n630), .A2(new_n452), .A3(new_n557), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT108), .ZN(new_n791));
  INV_X1    g590(.A(new_n774), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n771), .A2(KEYINPUT109), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n753), .A2(new_n770), .A3(new_n794), .A4(new_n754), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n792), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n793), .A2(KEYINPUT111), .A3(new_n795), .A4(new_n796), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n791), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n789), .B1(new_n801), .B2(KEYINPUT112), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n803));
  AOI211_X1 g602(.A(new_n803), .B(new_n791), .C1(new_n799), .C2(new_n800), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n789), .B(new_n806), .C1(new_n777), .C2(new_n790), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1337gat));
  XOR2_X1   g607(.A(KEYINPUT113), .B(G99gat), .Z(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n750), .B2(new_n680), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n713), .A2(new_n809), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n778), .A2(new_n630), .A3(new_n780), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1338gat));
  NAND3_X1  g612(.A1(new_n691), .A2(new_n439), .A3(new_n749), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT53), .B1(new_n814), .B2(G106gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n631), .A2(G106gat), .A3(new_n723), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n777), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n799), .B2(new_n800), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(G106gat), .B2(new_n814), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(G1339gat));
  NOR2_X1   g621(.A1(new_n632), .A2(new_n662), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n647), .A2(new_n648), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n825), .A2(new_n639), .A3(new_n641), .A4(new_n657), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n635), .B1(new_n634), .B2(new_n636), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n643), .A2(new_n644), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n656), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n604), .A3(new_n605), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT10), .ZN(new_n833));
  INV_X1    g632(.A(new_n617), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n614), .A2(new_n615), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n611), .B1(new_n836), .B2(new_n619), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n628), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n611), .A3(new_n619), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n621), .A2(new_n840), .A3(KEYINPUT54), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n841), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n629), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n832), .A2(new_n846), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n694), .A2(new_n846), .B1(new_n631), .B2(new_n830), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n606), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n824), .B1(new_n849), .B2(new_n731), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n385), .A2(new_n668), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n713), .A2(new_n851), .A3(new_n439), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G113gat), .B1(new_n854), .B2(new_n666), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n214), .A3(new_n662), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1340gat));
  NAND2_X1  g656(.A1(new_n853), .A2(new_n630), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g658(.A1(new_n853), .A2(new_n731), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g660(.A1(new_n854), .A2(new_n606), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n212), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT65), .B(G134gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(KEYINPUT56), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(KEYINPUT56), .B2(new_n865), .ZN(G1343gat));
  NOR2_X1   g666(.A1(new_n681), .A2(new_n851), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n606), .ZN(new_n869));
  INV_X1    g668(.A(new_n847), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n692), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n723), .B1(new_n872), .B2(new_n824), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT114), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n850), .A2(new_n439), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n846), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n844), .A2(KEYINPUT116), .A3(new_n629), .A4(new_n845), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n664), .A2(new_n881), .A3(new_n665), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT115), .B1(new_n831), .B2(new_n630), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n830), .A2(new_n631), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n755), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n692), .B1(new_n888), .B2(new_n847), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n877), .B(new_n723), .C1(new_n889), .C2(new_n824), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n868), .B1(new_n879), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G141gat), .B1(new_n891), .B2(new_n666), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n873), .A2(new_n868), .ZN(new_n893));
  INV_X1    g692(.A(new_n666), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n225), .A3(new_n894), .ZN(new_n895));
  XOR2_X1   g694(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G141gat), .B1(new_n891), .B2(new_n694), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n895), .B(KEYINPUT117), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(G1344gat));
  OR2_X1    g701(.A1(new_n222), .A2(new_n223), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(KEYINPUT59), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n891), .B2(new_n631), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT119), .B(new_n904), .C1(new_n891), .C2(new_n631), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n731), .B1(new_n869), .B2(new_n870), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT57), .B(new_n439), .C1(new_n909), .C2(new_n823), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT120), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n850), .A2(new_n912), .A3(KEYINPUT57), .A4(new_n439), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n894), .A2(new_n632), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n889), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT57), .B1(new_n916), .B2(new_n439), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n630), .B(new_n868), .C1(new_n914), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G148gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT59), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n907), .A2(new_n908), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n893), .A2(new_n903), .A3(new_n630), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1345gat));
  NOR3_X1   g722(.A1(new_n891), .A2(new_n229), .A3(new_n692), .ZN(new_n924));
  AOI21_X1  g723(.A(G155gat), .B1(new_n893), .B2(new_n731), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1346gat));
  OAI21_X1  g725(.A(G162gat), .B1(new_n891), .B2(new_n606), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n893), .A2(new_n230), .A3(new_n755), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1347gat));
  AOI21_X1  g728(.A(new_n668), .B1(new_n872), .B2(new_n824), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n743), .A2(new_n723), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n452), .A3(new_n931), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G169gat), .B1(new_n935), .B2(new_n666), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n452), .A3(new_n440), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n694), .A2(G169gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G1348gat));
  INV_X1    g738(.A(new_n937), .ZN(new_n940));
  AOI21_X1  g739(.A(G176gat), .B1(new_n940), .B2(new_n630), .ZN(new_n941));
  INV_X1    g740(.A(new_n935), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n630), .A2(G176gat), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G1349gat));
  OAI211_X1 g743(.A(new_n940), .B(new_n731), .C1(new_n283), .C2(new_n282), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n935), .A2(new_n692), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n302), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT60), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n949), .B(new_n945), .C1(new_n946), .C2(new_n302), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n940), .A2(new_n281), .A3(new_n755), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n942), .A2(new_n755), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(G190gat), .ZN(new_n955));
  AOI211_X1 g754(.A(KEYINPUT61), .B(new_n281), .C1(new_n942), .C2(new_n755), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1351gat));
  NOR3_X1   g756(.A1(new_n681), .A2(new_n668), .A3(new_n385), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n894), .B(new_n958), .C1(new_n914), .C2(new_n917), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G197gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n680), .A2(new_n452), .A3(new_n439), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT122), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n930), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n653), .A3(new_n662), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT123), .Z(G1352gat));
  NOR2_X1   g765(.A1(new_n631), .A2(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n930), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT124), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n930), .A2(new_n970), .A3(new_n962), .A4(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT62), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n914), .A2(new_n917), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n974), .A2(new_n630), .A3(new_n958), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G204gat), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n973), .A2(new_n976), .A3(KEYINPUT125), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1353gat));
  INV_X1    g780(.A(G211gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n982), .A3(new_n731), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n731), .B(new_n958), .C1(new_n914), .C2(new_n917), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(KEYINPUT126), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n989), .B(new_n983), .C1(new_n985), .C2(new_n986), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n990), .ZN(G1354gat));
  AOI21_X1  g790(.A(G218gat), .B1(new_n963), .B2(new_n755), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n974), .A2(new_n958), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n755), .A2(G218gat), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT127), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n992), .B1(new_n993), .B2(new_n995), .ZN(G1355gat));
endmodule


