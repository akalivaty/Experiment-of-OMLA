//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT64), .Z(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n214), .B1(new_n217), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n220), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n242), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(KEYINPUT67), .B1(new_n253), .B2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(new_n209), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G77), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n252), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n261), .A2(KEYINPUT11), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(KEYINPUT11), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n265));
  OR3_X1    g0065(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n266));
  INV_X1    g0066(.A(new_n264), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n251), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n220), .B1(new_n208), .B2(G20), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n265), .A2(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n262), .A2(new_n263), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(G274), .ZN(new_n277));
  INV_X1    g0077(.A(new_n274), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n276), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n279), .B2(new_n221), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G226), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G232), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n282), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G97), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n276), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT13), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n281), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT70), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT13), .B1(new_n280), .B2(new_n290), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n281), .A2(new_n291), .A3(KEYINPUT70), .A4(new_n292), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(G169), .A3(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n298), .A2(KEYINPUT14), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT14), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n296), .A2(new_n300), .A3(G169), .A4(new_n297), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n293), .A2(KEYINPUT71), .A3(G179), .A4(new_n295), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n293), .A2(G179), .A3(new_n295), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT71), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n301), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n271), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n295), .A2(G190), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n271), .B1(new_n293), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n296), .A2(G200), .A3(new_n297), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n254), .B2(new_n256), .ZN(new_n314));
  INV_X1    g0114(.A(G150), .ZN(new_n315));
  INV_X1    g0115(.A(new_n259), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n315), .A2(new_n316), .B1(new_n201), .B2(new_n209), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n251), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n243), .B1(new_n208), .B2(G20), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n268), .A2(new_n319), .B1(new_n243), .B2(new_n267), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT9), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n277), .B1(new_n279), .B2(new_n283), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G223), .A2(G1698), .ZN(new_n324));
  INV_X1    g0124(.A(G222), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(G1698), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n282), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n202), .B2(new_n282), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT66), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n276), .B1(new_n328), .B2(KEYINPUT66), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G190), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n322), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n331), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G200), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT69), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n333), .B(new_n335), .C1(new_n336), .C2(KEYINPUT10), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n322), .A3(new_n332), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n322), .A2(new_n336), .A3(new_n332), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT10), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n268), .ZN(new_n343));
  INV_X1    g0143(.A(new_n313), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n208), .A2(G20), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n343), .A2(new_n346), .B1(new_n264), .B2(new_n344), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT72), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G33), .ZN(new_n351));
  AOI21_X1  g0151(.A(G20), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n348), .B1(new_n352), .B2(KEYINPUT7), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n209), .A2(KEYINPUT7), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n282), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  OAI211_X1 g0157(.A(KEYINPUT72), .B(new_n357), .C1(new_n282), .C2(G20), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G68), .ZN(new_n360));
  AND2_X1   g0160(.A1(G58), .A2(G68), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G58), .A2(G68), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n259), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n252), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT73), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n350), .B2(G33), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n253), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n351), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n354), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n357), .B1(new_n282), .B2(G20), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n220), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n366), .B1(new_n376), .B2(new_n365), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n347), .B1(new_n368), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n283), .A2(G1698), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n282), .B(new_n379), .C1(G223), .C2(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n276), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n277), .B1(new_n279), .B2(new_n286), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G169), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n382), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT18), .B1(new_n378), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n349), .A2(new_n351), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT7), .B1(new_n391), .B2(new_n209), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n355), .B1(new_n392), .B2(KEYINPUT72), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n220), .B1(new_n393), .B2(new_n353), .ZN(new_n394));
  INV_X1    g0194(.A(new_n367), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n377), .B(new_n251), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n347), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n384), .A2(G179), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n385), .B2(new_n384), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n380), .A2(new_n381), .ZN(new_n403));
  INV_X1    g0203(.A(new_n276), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n383), .ZN(new_n406));
  INV_X1    g0206(.A(G190), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G200), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n382), .B2(new_n383), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n396), .A2(new_n397), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT17), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n396), .A2(KEYINPUT17), .A3(new_n411), .A4(new_n397), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n390), .A2(new_n402), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n321), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n334), .B2(new_n385), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G179), .B2(new_n334), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n282), .A2(new_n284), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n420), .A2(new_n286), .B1(new_n205), .B2(new_n282), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n391), .A2(new_n221), .A3(new_n284), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n404), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n277), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n404), .A2(new_n274), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n424), .B1(G244), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n387), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT68), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n257), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n344), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n252), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n268), .A2(G77), .A3(new_n345), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(G77), .B2(new_n264), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n427), .A2(new_n385), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n429), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n427), .A2(G200), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n435), .A2(new_n437), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(new_n442), .C1(new_n407), .C2(new_n427), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n419), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NOR4_X1   g0244(.A1(new_n312), .A2(new_n342), .A3(new_n416), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n272), .A3(KEYINPUT5), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT5), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(KEYINPUT76), .B2(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n273), .A2(G1), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n276), .A2(G274), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(G264), .A3(new_n276), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n282), .A2(G257), .A3(G1698), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G294), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n457), .C1(new_n420), .C2(new_n223), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n404), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT81), .B1(new_n460), .B2(G190), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT81), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n455), .A2(new_n459), .A3(new_n462), .A4(new_n407), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n409), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n282), .A2(new_n209), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT22), .B1(new_n466), .B2(new_n222), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT22), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n282), .A2(new_n468), .A3(new_n209), .A4(G87), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT23), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(G20), .B2(new_n205), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n209), .A2(KEYINPUT23), .A3(G107), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G116), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G20), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT79), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR4_X1   g0278(.A1(new_n472), .A2(new_n473), .A3(new_n475), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n476), .A2(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n470), .A2(new_n476), .A3(new_n477), .A4(new_n479), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n252), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n208), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n264), .A2(new_n486), .A3(new_n215), .A4(new_n250), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n487), .A2(KEYINPUT74), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(KEYINPUT74), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G107), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n264), .A2(G107), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT25), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n465), .A2(new_n485), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT19), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n209), .B1(new_n289), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(G87), .B2(new_n206), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n466), .B2(new_n220), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT19), .B1(new_n257), .B2(G97), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n251), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n430), .B(KEYINPUT68), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n267), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n488), .A2(G87), .A3(new_n489), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n282), .A2(G244), .A3(G1698), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n282), .A2(G238), .A3(new_n284), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(new_n474), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n404), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n276), .B(G250), .C1(G1), .C2(new_n273), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n276), .A2(G274), .A3(new_n450), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT77), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(KEYINPUT77), .A3(new_n513), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n511), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G200), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(new_n513), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT77), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(new_n515), .B1(new_n510), .B2(new_n404), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G190), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n507), .A2(new_n518), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n517), .A2(new_n385), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n522), .A2(new_n387), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n488), .A2(new_n489), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n502), .B(new_n504), .C1(new_n503), .C2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n460), .A2(KEYINPUT80), .A3(G169), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n455), .A2(new_n459), .A3(G179), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT80), .B1(new_n460), .B2(G169), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(new_n484), .B2(new_n494), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n496), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(new_n209), .C1(G33), .C2(new_n204), .ZN(new_n538));
  INV_X1    g0338(.A(G116), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G20), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n251), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT20), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n541), .B(new_n542), .ZN(new_n543));
  MUX2_X1   g0343(.A(new_n264), .B(new_n487), .S(G116), .Z(new_n544));
  AOI21_X1  g0344(.A(new_n385), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n282), .A2(G264), .A3(G1698), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n282), .A2(G257), .A3(new_n284), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n391), .A2(G303), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT78), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT78), .A4(new_n548), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n276), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n451), .A2(G270), .A3(new_n276), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n453), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n545), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT21), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT21), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n545), .B(new_n558), .C1(new_n553), .C2(new_n555), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n553), .A2(new_n555), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G190), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n543), .A2(new_n544), .ZN(new_n563));
  OAI21_X1  g0363(.A(G200), .B1(new_n553), .B2(new_n555), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OR4_X1    g0365(.A1(new_n387), .A2(new_n563), .A3(new_n553), .A4(new_n555), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n560), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n264), .A2(G97), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n490), .B2(G97), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT6), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n570), .A2(new_n204), .A3(G107), .ZN(new_n571));
  XNOR2_X1  g0371(.A(G97), .B(G107), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n573), .A2(new_n209), .B1(new_n202), .B2(new_n316), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n205), .B1(new_n374), .B2(new_n375), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n251), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n569), .A2(KEYINPUT75), .A3(new_n576), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n282), .A2(G250), .A3(G1698), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n282), .A2(G244), .A3(new_n284), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n537), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n391), .A2(G1698), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT4), .B1(new_n585), .B2(G244), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n404), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n451), .A2(G257), .A3(new_n276), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n453), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n407), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n585), .A2(KEYINPUT4), .A3(G244), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n582), .A2(new_n583), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n592), .A2(new_n537), .A3(new_n593), .A4(new_n581), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n589), .B1(new_n594), .B2(new_n404), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n591), .B1(new_n595), .B2(G200), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n579), .A2(new_n580), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(G179), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n587), .A2(new_n590), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G169), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n577), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n536), .A2(new_n567), .A3(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n445), .A2(new_n604), .ZN(G372));
  NAND2_X1  g0405(.A1(new_n390), .A2(new_n402), .ZN(new_n606));
  INV_X1    g0406(.A(new_n440), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n311), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n307), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n414), .A2(new_n415), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT83), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n342), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n337), .A2(new_n341), .A3(KEYINPUT83), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n419), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT84), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT84), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n618), .B(new_n419), .C1(new_n611), .C2(new_n615), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n535), .A2(new_n560), .A3(new_n566), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n506), .B1(G190), .B2(new_n522), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n518), .A2(KEYINPUT82), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT82), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n517), .B2(G200), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n622), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n496), .A2(new_n597), .A3(new_n626), .A4(new_n602), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n529), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n601), .A2(new_n524), .A3(new_n529), .A4(new_n577), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n579), .A2(new_n580), .B1(new_n600), .B2(new_n598), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(new_n529), .A3(new_n626), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n631), .B1(new_n633), .B2(new_n630), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n445), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n620), .A2(new_n636), .ZN(G369));
  INV_X1    g0437(.A(new_n567), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n563), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n638), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n560), .A2(new_n566), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n646), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n496), .A2(new_n535), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n644), .B1(new_n484), .B2(new_n494), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n535), .B2(new_n645), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n648), .A2(new_n644), .ZN(new_n657));
  INV_X1    g0457(.A(new_n535), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n657), .A2(new_n652), .B1(new_n658), .B2(new_n645), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT85), .ZN(G399));
  INV_X1    g0461(.A(new_n212), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n218), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT31), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n599), .A2(new_n553), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n511), .B(new_n554), .C1(new_n514), .C2(new_n516), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n532), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT30), .B1(new_n673), .B2(KEYINPUT86), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT86), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  AOI211_X1 g0476(.A(new_n675), .B(new_n676), .C1(new_n670), .C2(new_n672), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n599), .A2(new_n460), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT87), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n517), .A2(new_n387), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n561), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n522), .A2(G179), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n683), .B(KEYINPUT87), .C1(new_n555), .C2(new_n553), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n679), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(KEYINPUT88), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT88), .ZN(new_n687));
  AOI211_X1 g0487(.A(new_n687), .B(new_n679), .C1(new_n682), .C2(new_n684), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n678), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n669), .B1(new_n689), .B2(new_n645), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n645), .A2(new_n669), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n678), .B2(new_n685), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n496), .A2(new_n530), .A3(new_n535), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n597), .A2(new_n602), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(new_n638), .A3(new_n694), .A4(new_n645), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n690), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n535), .A2(new_n560), .A3(new_n566), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n694), .A2(new_n699), .A3(new_n496), .A4(new_n626), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n626), .A2(new_n529), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT89), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n632), .A3(new_n702), .A4(KEYINPUT26), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n629), .B2(new_n630), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n632), .A2(KEYINPUT26), .A3(new_n529), .A4(new_n626), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n700), .A2(new_n703), .A3(new_n706), .A4(new_n529), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n698), .B1(new_n707), .B2(new_n645), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n698), .B(new_n645), .C1(new_n628), .C2(new_n634), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n697), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n668), .B1(new_n712), .B2(G1), .ZN(G364));
  AND2_X1   g0513(.A1(new_n209), .A2(G13), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n208), .B1(new_n714), .B2(G45), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n663), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n215), .B1(G20), .B2(new_n385), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n209), .A2(new_n407), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n387), .A2(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n391), .B1(new_n724), .B2(G58), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n409), .A2(G179), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G87), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n209), .A2(G190), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n722), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n725), .B(new_n729), .C1(new_n202), .C2(new_n731), .ZN(new_n732));
  OR3_X1    g0532(.A1(new_n209), .A2(KEYINPUT91), .A3(G190), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT91), .B1(new_n209), .B2(G190), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n726), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n732), .B1(G107), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G179), .A2(G200), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n209), .B1(new_n738), .B2(G190), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n204), .ZN(new_n740));
  NAND3_X1  g0540(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n407), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n243), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n741), .A2(G190), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n740), .B(new_n744), .C1(G68), .C2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n733), .A2(new_n738), .A3(new_n734), .ZN(new_n747));
  INV_X1    g0547(.A(G159), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT32), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OR3_X1    g0549(.A1(new_n747), .A2(KEYINPUT32), .A3(new_n748), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n737), .A2(new_n746), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G322), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n723), .A2(new_n752), .B1(new_n731), .B2(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n282), .B(new_n754), .C1(G303), .C2(new_n728), .ZN(new_n755));
  INV_X1    g0555(.A(G326), .ZN(new_n756));
  INV_X1    g0556(.A(G294), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n743), .A2(new_n756), .B1(new_n739), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT33), .B(G317), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(new_n745), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n747), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G329), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n736), .A2(G283), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n755), .A2(new_n760), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n720), .B1(new_n751), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n719), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n662), .A2(new_n282), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G45), .B2(new_n218), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n248), .A2(new_n273), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n212), .A2(new_n282), .ZN(new_n774));
  INV_X1    g0574(.A(G355), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n774), .A2(new_n775), .B1(G116), .B2(new_n212), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n773), .B1(KEYINPUT90), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(KEYINPUT90), .B2(new_n776), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n718), .B(new_n765), .C1(new_n769), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n768), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n649), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n650), .A2(new_n718), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n649), .A2(G330), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT92), .Z(G396));
  NAND2_X1  g0585(.A1(new_n440), .A2(KEYINPUT96), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n438), .A2(KEYINPUT97), .A3(new_n644), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT97), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n442), .B2(new_n645), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT96), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n429), .A2(new_n438), .A3(new_n791), .A4(new_n439), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n786), .A2(new_n790), .A3(new_n443), .A4(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n645), .B(new_n794), .C1(new_n628), .C2(new_n634), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n635), .A2(new_n645), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n793), .B1(new_n440), .B2(new_n645), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n718), .B1(new_n798), .B2(new_n697), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n798), .A2(new_n697), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(KEYINPUT98), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(KEYINPUT98), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n720), .A2(new_n767), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n717), .B1(new_n803), .B2(G77), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n205), .A2(new_n727), .B1(new_n723), .B2(new_n757), .ZN(new_n805));
  INV_X1    g0605(.A(new_n731), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n282), .B(new_n805), .C1(G116), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G303), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n743), .A2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n740), .B(new_n809), .C1(G283), .C2(new_n745), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n761), .A2(G311), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n735), .A2(new_n222), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n807), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT34), .ZN(new_n815));
  XOR2_X1   g0615(.A(KEYINPUT93), .B(G143), .Z(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n724), .A2(new_n817), .B1(new_n806), .B2(G159), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  INV_X1    g0619(.A(new_n745), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(new_n743), .B2(new_n819), .C1(new_n315), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n736), .A2(G68), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n243), .B2(new_n727), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT94), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n815), .A2(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n815), .B2(new_n821), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n282), .B1(new_n747), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT95), .ZN(new_n830));
  INV_X1    g0630(.A(new_n739), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n829), .A2(new_n830), .B1(G58), .B2(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n830), .B2(new_n829), .C1(new_n824), .C2(new_n825), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n814), .B1(new_n827), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n804), .B1(new_n834), .B2(new_n719), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n797), .B2(new_n767), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n802), .A2(new_n836), .ZN(G384));
  INV_X1    g0637(.A(new_n573), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n838), .A2(KEYINPUT35), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(KEYINPUT35), .ZN(new_n840));
  NOR4_X1   g0640(.A1(new_n839), .A2(new_n840), .A3(new_n539), .A4(new_n217), .ZN(new_n841));
  XNOR2_X1  g0641(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n841), .B(new_n842), .ZN(new_n843));
  OR3_X1    g0643(.A1(new_n218), .A2(new_n361), .A3(new_n202), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n208), .B(G13), .C1(new_n844), .C2(new_n244), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G330), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT40), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT102), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n366), .B1(new_n394), .B2(new_n365), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n347), .B1(new_n850), .B2(new_n368), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n642), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n416), .A2(KEYINPUT100), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT100), .B1(new_n416), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n412), .B1(new_n851), .B2(new_n642), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n851), .A2(new_n389), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT37), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n412), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n389), .A2(new_n642), .B1(new_n396), .B2(new_n397), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT101), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT101), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT37), .B1(new_n378), .B2(new_n411), .ZN(new_n864));
  INV_X1    g0664(.A(new_n642), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n398), .B1(new_n401), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n858), .B1(new_n862), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT38), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n849), .B1(new_n855), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT101), .B1(new_n860), .B2(new_n861), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n864), .A2(new_n866), .A3(new_n863), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n871), .B1(new_n874), .B2(new_n858), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(KEYINPUT102), .C1(new_n854), .C2(new_n853), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n868), .B1(new_n853), .B2(new_n854), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n870), .A2(new_n876), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n271), .A2(new_n644), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n307), .A2(new_n311), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n307), .B2(new_n311), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n797), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n682), .A2(new_n684), .ZN(new_n883));
  INV_X1    g0683(.A(new_n679), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n687), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n673), .A2(KEYINPUT86), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n676), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n673), .A2(KEYINPUT86), .A3(KEYINPUT30), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n685), .A2(KEYINPUT88), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n892), .A2(new_n691), .B1(new_n604), .B2(new_n645), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n882), .B1(new_n690), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n848), .B1(new_n878), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n416), .A2(new_n852), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n416), .A2(KEYINPUT100), .A3(new_n852), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n875), .ZN(new_n902));
  XNOR2_X1  g0702(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n416), .A2(new_n398), .A3(new_n865), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n378), .A2(KEYINPUT104), .A3(new_n411), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT104), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n412), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n866), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n873), .A2(new_n872), .B1(new_n908), .B2(KEYINPUT37), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n903), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n848), .B1(new_n902), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n894), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n896), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n445), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n690), .B2(new_n893), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n847), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n913), .B2(new_n915), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n877), .A2(new_n871), .ZN(new_n918));
  INV_X1    g0718(.A(new_n876), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT102), .B1(new_n901), .B2(new_n875), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n880), .A2(new_n881), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n786), .A2(new_n792), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n645), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n795), .B2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n921), .A2(new_n925), .B1(new_n606), .B2(new_n642), .ZN(new_n926));
  OAI211_X1 g0726(.A(KEYINPUT39), .B(new_n918), .C1(new_n919), .C2(new_n920), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n307), .A2(new_n644), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT39), .B1(new_n902), .B2(new_n910), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n927), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n445), .B1(new_n708), .B2(new_n710), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n620), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n917), .A2(new_n936), .B1(new_n208), .B2(new_n714), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT105), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n917), .A2(new_n936), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n937), .B2(new_n938), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n846), .B1(new_n939), .B2(new_n941), .ZN(G367));
  NAND2_X1  g0742(.A1(new_n632), .A2(new_n644), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n645), .B1(new_n579), .B2(new_n580), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n603), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n659), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n659), .A2(new_n945), .ZN(new_n948));
  XOR2_X1   g0748(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n947), .A2(new_n656), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n656), .B1(new_n947), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n657), .A2(new_n652), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n655), .B2(new_n657), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n651), .B(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n712), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n712), .ZN(new_n958));
  XNOR2_X1  g0758(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n663), .B(new_n959), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n715), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n945), .B(KEYINPUT106), .Z(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n658), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(KEYINPUT107), .A3(new_n602), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n645), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT107), .B1(new_n965), .B2(new_n602), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n945), .A2(new_n657), .A3(new_n652), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT42), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n701), .B1(new_n507), .B2(new_n645), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n529), .A2(new_n507), .A3(new_n645), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT43), .Z(new_n976));
  NAND2_X1  g0776(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n978), .B(new_n971), .C1(new_n967), .C2(new_n968), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT108), .ZN(new_n980));
  INV_X1    g0780(.A(new_n656), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n964), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(KEYINPUT108), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n977), .A2(new_n980), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n977), .A2(new_n980), .A3(new_n984), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n982), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n963), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n769), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n770), .B2(new_n238), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n212), .B2(new_n503), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n717), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT111), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n728), .A2(G116), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT46), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n994), .A2(new_n995), .B1(new_n205), .B2(new_n739), .ZN(new_n996));
  INV_X1    g0796(.A(G317), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n204), .A2(new_n735), .B1(new_n747), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(G283), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n391), .B1(new_n731), .B2(new_n999), .C1(new_n808), .C2(new_n723), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n994), .A2(new_n995), .B1(new_n745), .B2(G294), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n753), .C2(new_n743), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT112), .Z(new_n1004));
  OAI22_X1  g0804(.A1(new_n743), .A2(new_n816), .B1(new_n220), .B2(new_n739), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n723), .A2(new_n315), .B1(new_n731), .B2(new_n243), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n391), .B(new_n1006), .C1(G58), .C2(new_n728), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n736), .A2(G77), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n819), .C2(new_n747), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1005), .B(new_n1009), .C1(G159), .C2(new_n745), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1011), .A2(KEYINPUT47), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n719), .B1(new_n1011), .B2(KEYINPUT47), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n993), .B1(new_n975), .B2(new_n780), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n988), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(KEYINPUT113), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1014), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n962), .A2(new_n715), .B1(new_n986), .B2(new_n982), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n985), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT113), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1016), .A2(new_n1021), .ZN(G387));
  OR2_X1    g0822(.A1(new_n655), .A2(new_n780), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n774), .A2(new_n665), .B1(G107), .B2(new_n212), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n235), .A2(G45), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n770), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n665), .ZN(new_n1027));
  AOI211_X1 g0827(.A(G45), .B(new_n1027), .C1(G68), .C2(G77), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n313), .A2(G50), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1026), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1024), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n717), .B1(new_n1032), .B2(new_n989), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n727), .A2(new_n202), .B1(new_n731), .B2(new_n220), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n391), .B(new_n1034), .C1(G50), .C2(new_n724), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n344), .A2(new_n745), .B1(G159), .B2(new_n742), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n432), .A2(new_n831), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G97), .A2(new_n736), .B1(new_n761), .B2(G150), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n727), .A2(new_n757), .B1(new_n739), .B2(new_n999), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G317), .A2(new_n724), .B1(new_n806), .B2(G303), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n743), .B2(new_n752), .C1(new_n753), .C2(new_n820), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT114), .Z(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(KEYINPUT49), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n391), .B1(new_n735), .B2(new_n539), .C1(new_n756), .C2(new_n747), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT115), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1046), .A2(KEYINPUT49), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1039), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1033), .B1(new_n1052), .B2(new_n719), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n956), .A2(new_n716), .B1(new_n1023), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n712), .A2(new_n956), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n663), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n712), .A2(new_n956), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(G393));
  OAI21_X1  g0858(.A(new_n1055), .B1(new_n951), .B2(new_n952), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n957), .A2(new_n663), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n953), .A2(new_n716), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n769), .B1(new_n204), .B2(new_n212), .C1(new_n1026), .C2(new_n242), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n717), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n739), .A2(new_n202), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n313), .B2(new_n731), .C1(new_n820), .C2(new_n243), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT116), .Z(new_n1067));
  AOI211_X1 g0867(.A(new_n391), .B(new_n812), .C1(G68), .C2(new_n728), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n743), .A2(new_n315), .B1(new_n723), .B2(new_n748), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1068), .B(new_n1070), .C1(new_n747), .C2(new_n816), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n724), .A2(G311), .B1(G317), .B2(new_n742), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n205), .A2(new_n735), .B1(new_n747), .B2(new_n752), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n391), .B1(new_n731), .B2(new_n757), .C1(new_n999), .C2(new_n727), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n820), .A2(new_n808), .B1(new_n739), .B2(new_n539), .ZN(new_n1076));
  OR3_X1    g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1067), .A2(new_n1071), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1063), .B1(new_n1078), .B2(new_n719), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n964), .B2(new_n780), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1060), .A2(new_n1061), .A3(new_n1080), .ZN(G390));
  INV_X1    g0881(.A(new_n882), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n691), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n695), .B1(new_n689), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT31), .B1(new_n892), .B2(new_n644), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1082), .B(G330), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n795), .A2(new_n924), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n922), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n929), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n927), .B2(new_n931), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n902), .A2(new_n910), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n928), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n707), .A2(new_n645), .A3(new_n794), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n924), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1087), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1094), .A2(new_n924), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n928), .B(new_n1092), .C1(new_n1098), .C2(new_n922), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n696), .A2(G330), .A3(new_n797), .A4(new_n1089), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n930), .B1(new_n878), .B2(KEYINPUT39), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1099), .B(new_n1100), .C1(new_n1101), .C2(new_n1090), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1097), .A2(new_n1102), .A3(new_n716), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n717), .B1(new_n803), .B2(new_n344), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G116), .A2(new_n724), .B1(new_n806), .B2(G97), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n822), .A2(new_n1105), .A3(new_n391), .A4(new_n729), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1065), .B1(new_n743), .B2(new_n999), .C1(new_n205), .C2(new_n820), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G294), .C2(new_n761), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1109), .A2(KEYINPUT118), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(KEYINPUT118), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n831), .A2(G159), .B1(G128), .B2(new_n742), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT53), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n727), .A2(new_n315), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G50), .A2(new_n736), .B1(new_n761), .B2(G125), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n282), .B1(new_n723), .B2(new_n828), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1117), .B1(new_n806), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1114), .A2(new_n1113), .B1(G137), .B2(new_n745), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1116), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1110), .B(new_n1111), .C1(new_n1115), .C2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1104), .B1(new_n1123), .B2(new_n719), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1101), .B2(new_n767), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1103), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT117), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n690), .A2(new_n893), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(G330), .A3(new_n445), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n620), .A2(new_n934), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n695), .A2(new_n692), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n797), .C1(new_n1085), .C2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n922), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1086), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1088), .ZN(new_n1137));
  OAI211_X1 g0937(.A(G330), .B(new_n797), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n922), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n1100), .A3(new_n1098), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1132), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1129), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1141), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1144));
  AND4_X1   g0944(.A1(new_n1128), .A2(new_n1143), .A3(new_n663), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n664), .B1(new_n1129), .B2(new_n1142), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1128), .B1(new_n1146), .B2(new_n1144), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1127), .B1(new_n1145), .B2(new_n1147), .ZN(G378));
  AOI21_X1  g0948(.A(KEYINPUT40), .B1(new_n921), .B2(new_n894), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n912), .A2(G330), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n613), .A2(new_n419), .A3(new_n614), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n417), .A2(new_n642), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1152), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n613), .A2(new_n419), .A3(new_n614), .A4(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1157), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1149), .A2(new_n1150), .A3(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1156), .B(new_n1158), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n847), .B1(new_n911), .B2(new_n894), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n896), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n933), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1161), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n896), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1167), .A2(new_n1168), .A3(new_n932), .A4(new_n926), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1132), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1144), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1172), .A3(KEYINPUT57), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1169), .A2(new_n1166), .B1(new_n1144), .B2(new_n1171), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n663), .C1(KEYINPUT57), .C2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1161), .A2(new_n766), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n717), .B1(new_n803), .B2(G50), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n282), .A2(G41), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n723), .B2(new_n205), .C1(new_n202), .C2(new_n727), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n432), .B2(new_n806), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n739), .A2(new_n220), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n743), .A2(new_n539), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G97), .C2(new_n745), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G58), .A2(new_n736), .B1(new_n761), .B2(G283), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT58), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n243), .B1(G33), .B2(G41), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n820), .A2(new_n828), .B1(new_n739), .B2(new_n315), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G128), .A2(new_n724), .B1(new_n728), .B2(new_n1119), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n819), .B2(new_n731), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(G125), .C2(new_n742), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n253), .B(new_n272), .C1(new_n735), .C2(new_n748), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G124), .B2(new_n761), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT59), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1195), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1186), .B1(new_n1178), .B2(new_n1187), .C1(new_n1193), .C2(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT119), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n720), .B1(new_n1198), .B2(KEYINPUT119), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1177), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1170), .A2(new_n716), .B1(new_n1176), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1175), .A2(new_n1202), .ZN(G375));
  AOI21_X1  g1003(.A(new_n715), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n922), .A2(new_n766), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n717), .B1(new_n803), .B2(G68), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n747), .A2(new_n808), .B1(new_n204), .B2(new_n727), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT120), .Z(new_n1209));
  OAI21_X1  g1009(.A(new_n391), .B1(new_n723), .B2(new_n999), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n820), .A2(new_n539), .B1(new_n743), .B2(new_n757), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(G107), .C2(new_n806), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1008), .A3(new_n1037), .A4(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT121), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n724), .A2(G137), .B1(new_n1119), .B2(new_n745), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n828), .B2(new_n743), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(KEYINPUT122), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(KEYINPUT122), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n282), .B1(new_n731), .B2(new_n315), .C1(new_n748), .C2(new_n727), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G50), .B2(new_n831), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G58), .A2(new_n736), .B1(new_n761), .B2(G128), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1217), .A2(new_n1218), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT123), .B1(new_n1214), .B2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(new_n720), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1214), .A2(KEYINPUT123), .A3(new_n1222), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1207), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1206), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1205), .A2(KEYINPUT124), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT124), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1227), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1229), .B1(new_n1204), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1137), .A2(new_n1140), .A3(new_n1132), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1142), .A2(new_n1233), .A3(new_n961), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(G381));
  AND2_X1   g1035(.A1(new_n1146), .A2(new_n1144), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(new_n1126), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G387), .A2(G375), .A3(new_n1238), .A4(new_n1240), .ZN(G407));
  NAND2_X1  g1041(.A1(new_n643), .A2(G213), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1237), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G407), .B(G213), .C1(G375), .C2(new_n1244), .ZN(G409));
  XNOR2_X1  g1045(.A(G393), .B(G396), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1019), .A2(KEYINPUT126), .A3(G390), .ZN(new_n1248));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1015), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT126), .B1(new_n1019), .B2(G390), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1247), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1016), .A2(new_n1021), .A3(new_n1249), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1247), .B1(new_n1019), .B2(G390), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(G378), .A2(new_n1202), .A3(new_n1175), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1174), .A2(new_n961), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1202), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1237), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1243), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1233), .B1(new_n1141), .B2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1137), .A2(new_n1140), .A3(KEYINPUT60), .A4(new_n1132), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n663), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1232), .A2(new_n1266), .A3(G384), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(G384), .B1(new_n1232), .B2(new_n1266), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1262), .A2(KEYINPUT63), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(new_n1242), .A3(new_n1270), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1243), .A2(G2897), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1268), .A2(new_n1269), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1232), .A2(new_n1266), .ZN(new_n1278));
  INV_X1    g1078(.A(G384), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1280), .A2(new_n1267), .B1(G2897), .B2(new_n1243), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT125), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1272), .A2(new_n1242), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1284), .A2(new_n1285), .A3(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1257), .A2(new_n1271), .A3(new_n1275), .A4(new_n1288), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1262), .B2(new_n1282), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1273), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1262), .A2(KEYINPUT62), .A3(new_n1270), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1292), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1290), .B1(new_n1296), .B2(KEYINPUT127), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1283), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1295), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT62), .B1(new_n1262), .B2(new_n1270), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1298), .B(KEYINPUT127), .C1(new_n1299), .C2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1289), .B1(new_n1297), .B2(new_n1302), .ZN(G405));
  NAND2_X1  g1103(.A1(G375), .A2(new_n1237), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1304), .A2(new_n1258), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1270), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1305), .B(new_n1306), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1290), .B(new_n1307), .ZN(G402));
endmodule


