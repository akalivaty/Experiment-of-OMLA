//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0002(.A(G50), .B1(G58), .B2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G1), .A2(G13), .ZN(new_n205));
  OR3_X1    g0005(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n206), .B(new_n210), .C1(new_n217), .C2(KEYINPUT1), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(KEYINPUT1), .B2(new_n217), .ZN(G361));
  XNOR2_X1  g0019(.A(G238), .B(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n220), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT2), .B(G226), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n222), .B(new_n223), .Z(new_n224));
  XNOR2_X1  g0024(.A(G250), .B(G257), .ZN(new_n225));
  XNOR2_X1  g0025(.A(G264), .B(G270), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n224), .B(new_n227), .Z(G358));
  XOR2_X1   g0028(.A(G50), .B(G58), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G68), .B(G77), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G87), .B(G97), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XOR2_X1   g0034(.A(G107), .B(G116), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G351));
  INV_X1    g0037(.A(G33), .ZN(new_n238));
  INV_X1    g0038(.A(G41), .ZN(new_n239));
  OAI211_X1 g0039(.A(G1), .B(G13), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G274), .ZN(new_n241));
  INV_X1    g0041(.A(G45), .ZN(new_n242));
  AOI21_X1  g0042(.A(G1), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n240), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(new_n243), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n245), .B1(G226), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(KEYINPUT67), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n238), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G222), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(new_n257), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n257), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT68), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT68), .B1(new_n257), .B2(G1698), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n261), .B1(new_n266), .B2(G223), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n248), .B1(new_n267), .B2(new_n240), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(G179), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n205), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT8), .B(G58), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n204), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G150), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI22_X1  g0076(.A1(new_n272), .A2(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G50), .A2(G58), .ZN(new_n278));
  INV_X1    g0078(.A(G68), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n204), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n271), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n271), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G50), .A3(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n281), .B(new_n287), .C1(G50), .C2(new_n283), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n268), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n269), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n268), .A2(G200), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n293), .B(new_n297), .C1(new_n298), .C2(new_n268), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n292), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G50), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n276), .A2(new_n303), .B1(new_n204), .B2(G68), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n273), .A2(new_n260), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n271), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT11), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n284), .A2(new_n279), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT12), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n285), .A2(G68), .A3(new_n286), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(KEYINPUT72), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT72), .B1(new_n309), .B2(new_n310), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT73), .A2(G169), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n257), .A2(G226), .A3(new_n258), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT70), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT70), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n257), .A2(new_n319), .A3(G226), .A4(new_n258), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n221), .B1(new_n251), .B2(new_n256), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n240), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n245), .B1(G238), .B2(new_n247), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT13), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n257), .A2(G232), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n258), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n320), .B2(new_n318), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n328), .B(new_n325), .C1(new_n332), .C2(new_n240), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n316), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n327), .A2(new_n333), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n334), .A2(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI211_X1 g0138(.A(KEYINPUT14), .B(new_n316), .C1(new_n327), .C2(new_n333), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n315), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n327), .A2(new_n333), .A3(G190), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT71), .B1(new_n336), .B2(G200), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT71), .ZN(new_n343));
  INV_X1    g0143(.A(G200), .ZN(new_n344));
  AOI211_X1 g0144(.A(new_n343), .B(new_n344), .C1(new_n327), .C2(new_n333), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n314), .B(new_n341), .C1(new_n342), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n245), .B1(G244), .B2(new_n247), .ZN(new_n349));
  OAI21_X1  g0149(.A(G238), .B1(new_n264), .B2(new_n265), .ZN(new_n350));
  INV_X1    g0150(.A(new_n257), .ZN(new_n351));
  AOI22_X1  g0151(.A1(G107), .A2(new_n351), .B1(new_n322), .B2(new_n258), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n337), .B(new_n349), .C1(new_n353), .C2(new_n240), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n240), .B1(new_n350), .B2(new_n352), .ZN(new_n355));
  INV_X1    g0155(.A(new_n349), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n289), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n272), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n275), .B1(G20), .B2(G77), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n273), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n271), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n285), .A2(G77), .A3(new_n286), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n362), .B(new_n363), .C1(G77), .C2(new_n283), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n354), .A2(new_n357), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n349), .B1(new_n353), .B2(new_n240), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n364), .B1(new_n366), .B2(G200), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n298), .B2(new_n366), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n302), .A2(new_n348), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G58), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(new_n279), .ZN(new_n371));
  NOR2_X1   g0171(.A1(G58), .A2(G68), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n275), .A2(G159), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  OR2_X1    g0177(.A1(KEYINPUT74), .A2(G33), .ZN(new_n378));
  NAND2_X1  g0178(.A1(KEYINPUT74), .A2(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n250), .B1(new_n380), .B2(KEYINPUT3), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(new_n381), .B2(new_n204), .ZN(new_n382));
  AND2_X1   g0182(.A1(KEYINPUT74), .A2(G33), .ZN(new_n383));
  NOR2_X1   g0183(.A1(KEYINPUT74), .A2(G33), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT3), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n385), .A2(new_n377), .A3(new_n204), .A4(new_n253), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G68), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n376), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n271), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT7), .A2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n251), .A2(new_n256), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n255), .A2(new_n204), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n383), .A2(new_n384), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n252), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n392), .B(G68), .C1(new_n395), .C2(new_n377), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n376), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT75), .B1(new_n397), .B2(new_n389), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT75), .ZN(new_n399));
  AOI211_X1 g0199(.A(new_n399), .B(KEYINPUT16), .C1(new_n396), .C2(new_n376), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n390), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n285), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n358), .A2(new_n286), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n402), .A2(new_n403), .B1(new_n283), .B2(new_n358), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT76), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n397), .A2(new_n389), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n399), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n270), .A2(new_n205), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n386), .A2(G68), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n385), .A2(new_n253), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT7), .B1(new_n410), .B2(G20), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n375), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n408), .B1(new_n412), .B2(KEYINPUT16), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n397), .A2(KEYINPUT75), .A3(new_n389), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n407), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT76), .ZN(new_n416));
  INV_X1    g0216(.A(new_n404), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(G223), .A2(G1698), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G226), .B2(new_n258), .ZN(new_n420));
  INV_X1    g0220(.A(G87), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n381), .A2(new_n420), .B1(new_n238), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n246), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n245), .B1(G232), .B2(new_n247), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n289), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n423), .A2(new_n424), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(G179), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n405), .A2(new_n418), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT18), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n405), .A2(new_n431), .A3(new_n418), .A4(new_n428), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n398), .A2(new_n400), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n404), .B1(new_n433), .B2(new_n413), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n344), .B1(new_n423), .B2(new_n424), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(G190), .B2(new_n426), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT17), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AND4_X1   g0237(.A1(KEYINPUT17), .A2(new_n415), .A3(new_n417), .A4(new_n436), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n430), .A2(new_n432), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n369), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G97), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n284), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n282), .A2(G33), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n408), .A2(new_n283), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n445), .B2(new_n442), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n392), .B(G107), .C1(new_n395), .C2(new_n377), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT77), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT7), .B1(new_n450), .B2(new_n393), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(KEYINPUT77), .A3(G107), .A4(new_n392), .ZN(new_n452));
  INV_X1    g0252(.A(G107), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(KEYINPUT6), .A3(G97), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n442), .A2(new_n453), .ZN(new_n455));
  NOR2_X1   g0255(.A1(G97), .A2(G107), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n457), .B2(KEYINPUT6), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(G20), .B1(G77), .B2(new_n275), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n449), .A2(new_n452), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n446), .B1(new_n460), .B2(new_n271), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n258), .A2(G244), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n385), .B2(new_n253), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n467), .B2(KEYINPUT4), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n246), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n242), .A2(G1), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n472), .A2(new_n240), .A3(G274), .A4(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n470), .B2(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n240), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G257), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n469), .A2(G190), .A3(new_n474), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n469), .A2(new_n474), .A3(new_n478), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n461), .B(new_n479), .C1(new_n481), .C2(new_n344), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n460), .A2(new_n271), .ZN(new_n483));
  INV_X1    g0283(.A(new_n446), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n480), .A2(new_n289), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n469), .A2(new_n337), .A3(new_n474), .A4(new_n478), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OR2_X1    g0288(.A1(G238), .A2(G1698), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(G244), .B2(new_n258), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n253), .B2(new_n385), .ZN(new_n491));
  INV_X1    g0291(.A(G116), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n394), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n246), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n282), .A2(G45), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n495), .A2(G250), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n240), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n241), .B2(new_n495), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G200), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n381), .A2(new_n490), .B1(new_n492), .B2(new_n394), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n498), .B1(new_n502), .B2(new_n246), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G190), .ZN(new_n504));
  AOI21_X1  g0304(.A(G20), .B1(new_n385), .B2(new_n253), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G68), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT19), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n204), .B1(new_n329), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n456), .A2(new_n421), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n204), .A2(G33), .A3(G97), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n508), .A2(new_n509), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n512), .A2(new_n271), .B1(new_n284), .B2(new_n360), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n408), .A2(new_n283), .A3(new_n444), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G87), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n501), .A2(new_n504), .A3(new_n513), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n512), .A2(new_n271), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n360), .A2(new_n284), .ZN(new_n518));
  INV_X1    g0318(.A(new_n360), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n503), .A2(new_n337), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n500), .A2(new_n289), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n482), .A2(new_n488), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n465), .B(new_n204), .C1(G33), .C2(new_n442), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT80), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n492), .A2(G20), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n271), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n271), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(KEYINPUT20), .B(new_n527), .C1(new_n530), .C2(new_n531), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n514), .A2(new_n537), .A3(G116), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT79), .B1(new_n445), .B2(new_n492), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n538), .A2(new_n539), .B1(new_n492), .B2(new_n284), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n289), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(G257), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n258), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n258), .A2(G264), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n410), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n251), .A2(new_n256), .A3(G303), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n240), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G270), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n474), .B1(new_n476), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT78), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(new_n546), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n246), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT78), .ZN(new_n553));
  INV_X1    g0353(.A(new_n549), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n541), .A2(new_n550), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n547), .A2(KEYINPUT78), .A3(new_n549), .ZN(new_n560));
  OAI21_X1  g0360(.A(G190), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n536), .A2(new_n540), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n555), .A2(new_n550), .A3(G200), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n547), .A2(new_n337), .A3(new_n549), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n541), .A2(KEYINPUT21), .A3(new_n550), .A4(new_n555), .ZN(new_n568));
  AND4_X1   g0368(.A1(new_n558), .A2(new_n565), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT24), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT22), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n505), .B2(G87), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n204), .A3(G87), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT81), .B1(new_n257), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT81), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n576), .B(new_n573), .C1(new_n251), .C2(new_n256), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n572), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n204), .B(G116), .C1(new_n383), .C2(new_n384), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT23), .B1(new_n204), .B2(G107), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT23), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n453), .A3(G20), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT82), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT82), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n579), .A2(new_n586), .A3(new_n581), .A4(new_n583), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(KEYINPUT83), .B(new_n570), .C1(new_n578), .C2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n575), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n252), .B1(new_n378), .B2(new_n379), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n204), .B(G87), .C1(new_n591), .C2(new_n250), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT22), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n257), .A2(KEYINPUT81), .A3(new_n574), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT83), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n585), .A2(new_n587), .B1(new_n596), .B2(KEYINPUT24), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n595), .B(new_n597), .C1(new_n596), .C2(KEYINPUT24), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n589), .A2(new_n598), .A3(new_n271), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n542), .A2(G1698), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(G250), .B2(G1698), .ZN(new_n601));
  INV_X1    g0401(.A(G294), .ZN(new_n602));
  OAI22_X1  g0402(.A1(new_n381), .A2(new_n601), .B1(new_n602), .B2(new_n394), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n475), .A2(G264), .A3(new_n240), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT86), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT86), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n475), .A2(new_n606), .A3(G264), .A4(new_n240), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n603), .A2(new_n246), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n344), .B1(new_n608), .B2(new_n474), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n607), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n601), .B1(new_n253), .B2(new_n385), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n394), .A2(new_n602), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n246), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n474), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(new_n298), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT25), .ZN(new_n618));
  AOI21_X1  g0418(.A(G107), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n284), .B(new_n619), .C1(new_n617), .C2(new_n618), .ZN(new_n620));
  OAI211_X1 g0420(.A(KEYINPUT84), .B(KEYINPUT25), .C1(new_n283), .C2(G107), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n621), .C1(new_n445), .C2(new_n453), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(KEYINPUT85), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n599), .A2(new_n616), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n289), .B1(new_n608), .B2(new_n474), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n614), .A2(new_n337), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT87), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n614), .A2(G169), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT87), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n629), .B(new_n630), .C1(new_n337), .C2(new_n614), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n595), .A2(new_n597), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n596), .A2(KEYINPUT24), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n408), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n623), .B1(new_n635), .B2(new_n598), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n625), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n441), .A2(new_n526), .A3(new_n569), .A4(new_n638), .ZN(G372));
  NAND2_X1  g0439(.A1(new_n526), .A2(new_n625), .ZN(new_n640));
  INV_X1    g0440(.A(new_n636), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n626), .B2(new_n627), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n558), .A2(new_n567), .A3(new_n568), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n516), .A2(new_n524), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n488), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n524), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n441), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n300), .A2(new_n301), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n415), .A2(new_n417), .A3(new_n436), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT17), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n434), .A2(KEYINPUT17), .A3(new_n436), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n365), .A2(KEYINPUT88), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT88), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n354), .A2(new_n357), .A3(new_n657), .A4(new_n364), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n346), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n655), .B1(new_n659), .B2(new_n340), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT18), .B1(new_n434), .B2(new_n427), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n428), .B(new_n431), .C1(new_n401), .C2(new_n404), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n650), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n291), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n649), .A2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n282), .A2(new_n204), .A3(G13), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n642), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n643), .A2(new_n673), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n638), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT89), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT89), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n558), .A2(new_n567), .A3(new_n568), .ZN(new_n680));
  INV_X1    g0480(.A(new_n673), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n563), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n569), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n632), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n641), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n636), .A2(new_n681), .ZN(new_n690));
  OAI22_X1  g0490(.A1(new_n689), .A2(new_n681), .B1(new_n637), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n679), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n208), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n509), .A2(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n203), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT90), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n566), .A2(new_n469), .A3(new_n478), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT92), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n610), .A2(new_n613), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(new_n500), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n608), .A2(new_n503), .A3(KEYINPUT92), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n702), .A2(new_n707), .A3(KEYINPUT30), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT30), .B1(new_n702), .B2(new_n707), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n503), .A2(G179), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n555), .A3(new_n550), .A4(new_n614), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n481), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n681), .ZN(new_n714));
  XNOR2_X1  g0514(.A(KEYINPUT91), .B(KEYINPUT31), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT93), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT93), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n714), .A2(new_n719), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n638), .A2(new_n569), .A3(new_n526), .A4(new_n681), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n714), .B1(new_n722), .B2(KEYINPUT31), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n681), .B1(new_n648), .B2(new_n644), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n680), .B1(new_n641), .B2(new_n688), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n647), .B(new_n524), .C1(new_n729), .C2(new_n640), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n728), .B1(new_n730), .B2(new_n681), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n701), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(G13), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n282), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n695), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n687), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G330), .B2(new_n685), .ZN(new_n741));
  INV_X1    g0541(.A(new_n739), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n204), .A2(G179), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G190), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G159), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT32), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n204), .A2(new_n337), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n750), .A2(new_n344), .A3(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n298), .A2(new_n344), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n749), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n751), .A2(G68), .B1(new_n754), .B2(G50), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n743), .A2(new_n298), .A3(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G107), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n749), .A2(new_n744), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G77), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n748), .A2(new_n755), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n750), .A2(new_n298), .A3(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G58), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n298), .A2(G179), .A3(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n204), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G97), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n752), .A2(new_n743), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G87), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n764), .A2(new_n768), .A3(new_n257), .A4(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n763), .A2(G322), .B1(G311), .B2(new_n760), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n773), .B(new_n351), .C1(new_n602), .C2(new_n766), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n745), .B(KEYINPUT95), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G329), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n751), .A2(new_n777), .B1(new_n754), .B2(G326), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G283), .A2(new_n757), .B1(new_n770), .B2(G303), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n762), .A2(new_n772), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n205), .B1(G20), .B2(new_n289), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n410), .A2(new_n694), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n203), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(new_n242), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n232), .B2(new_n242), .ZN(new_n788));
  INV_X1    g0588(.A(G355), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n257), .A2(new_n208), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT94), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n788), .B1(G116), .B2(new_n208), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n782), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n742), .B(new_n783), .C1(new_n792), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n795), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n685), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n741), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n364), .A2(new_n673), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n368), .A2(new_n365), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n656), .A2(new_n364), .A3(new_n658), .A4(new_n673), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT98), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n726), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n681), .B(new_n805), .C1(new_n648), .C2(new_n644), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(new_n725), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n725), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n812), .A2(new_n742), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n782), .A2(new_n793), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n742), .B1(new_n260), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n782), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n763), .A2(G143), .B1(new_n754), .B2(G137), .ZN(new_n818));
  INV_X1    g0618(.A(new_n751), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n274), .B2(new_n819), .C1(new_n746), .C2(new_n759), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n769), .A2(new_n303), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n756), .A2(new_n279), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(G58), .C2(new_n767), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n381), .B1(new_n775), .B2(G132), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT97), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n821), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n763), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n768), .B1(new_n828), .B2(new_n602), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT96), .Z(new_n830));
  AOI22_X1  g0630(.A1(new_n751), .A2(G283), .B1(G87), .B2(new_n757), .ZN(new_n831));
  INV_X1    g0631(.A(G303), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(new_n753), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n453), .A2(new_n769), .B1(new_n759), .B2(new_n492), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n833), .A2(new_n257), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G311), .ZN(new_n836));
  INV_X1    g0636(.A(new_n775), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n830), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n827), .A2(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n816), .B1(new_n817), .B2(new_n839), .C1(new_n805), .C2(new_n794), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n814), .A2(new_n840), .ZN(G384));
  NOR2_X1   g0641(.A1(new_n736), .A2(new_n282), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n365), .A2(new_n673), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n809), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n315), .A2(new_n673), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n340), .A2(new_n346), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(new_n340), .B2(new_n346), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n412), .A2(KEYINPUT16), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n417), .B1(new_n853), .B2(new_n390), .ZN(new_n854));
  INV_X1    g0654(.A(new_n671), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n655), .B1(KEYINPUT18), .B2(new_n429), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n432), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n405), .A2(new_n418), .A3(new_n855), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT37), .B1(new_n434), .B2(new_n436), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n429), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n428), .A2(new_n854), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(new_n651), .A3(new_n856), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n852), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n856), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n440), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n851), .A2(new_n871), .B1(new_n663), .B2(new_n671), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT39), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n867), .B2(new_n870), .ZN(new_n874));
  INV_X1    g0674(.A(new_n859), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n663), .B2(new_n655), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n429), .A2(new_n859), .A3(new_n860), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n415), .A2(new_n417), .A3(new_n436), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n427), .B1(new_n415), .B2(new_n417), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n878), .B1(new_n881), .B2(new_n859), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n876), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n852), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n870), .A2(new_n884), .A3(new_n873), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT100), .B1(new_n874), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n340), .A2(new_n673), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI221_X4 g0688(.A(new_n852), .B1(new_n861), .B2(new_n864), .C1(new_n440), .C2(new_n868), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n869), .B2(new_n865), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT39), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT100), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n870), .A2(new_n884), .A3(new_n873), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n886), .A2(new_n888), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n872), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n441), .B1(new_n727), .B2(new_n731), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n666), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n896), .B(new_n898), .Z(new_n899));
  OAI21_X1  g0699(.A(new_n715), .B1(new_n713), .B2(new_n681), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n709), .A2(new_n712), .ZN(new_n901));
  OAI211_X1 g0701(.A(KEYINPUT31), .B(new_n673), .C1(new_n901), .C2(new_n708), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n722), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(new_n805), .C1(new_n848), .C2(new_n849), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n870), .A2(new_n884), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT40), .B1(new_n867), .B2(new_n870), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n907), .A2(KEYINPUT40), .B1(new_n908), .B2(new_n905), .ZN(new_n909));
  INV_X1    g0709(.A(new_n441), .ZN(new_n910));
  INV_X1    g0710(.A(new_n903), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n889), .B2(new_n890), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(new_n904), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n913), .B1(new_n905), .B2(new_n906), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n441), .B(new_n903), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n912), .A2(new_n917), .A3(G330), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n842), .B1(new_n899), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n899), .B2(new_n918), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n205), .A2(new_n204), .A3(new_n492), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n458), .B(KEYINPUT99), .Z(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT35), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n924), .B2(new_n923), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT36), .Z(new_n927));
  NOR3_X1   g0727(.A1(new_n371), .A2(new_n203), .A3(new_n260), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n279), .A2(G50), .ZN(new_n929));
  OAI211_X1 g0729(.A(G1), .B(new_n735), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n920), .A2(new_n927), .A3(new_n930), .ZN(G367));
  NAND2_X1  g0731(.A1(new_n227), .A2(new_n784), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n782), .B(new_n795), .C1(new_n694), .C2(new_n519), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n742), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n513), .A2(new_n515), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n673), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n525), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n936), .A2(new_n524), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(KEYINPUT101), .A3(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n938), .A2(KEYINPUT101), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n756), .A2(new_n442), .ZN(new_n943));
  INV_X1    g0743(.A(G283), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n753), .A2(new_n836), .B1(new_n759), .B2(new_n944), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n943), .B(new_n945), .C1(G294), .C2(new_n751), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n767), .A2(G107), .ZN(new_n947));
  INV_X1    g0747(.A(G317), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n745), .A2(new_n948), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n410), .B(new_n949), .C1(G303), .C2(new_n763), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n770), .A2(G116), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT46), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n946), .A2(new_n947), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n766), .A2(new_n279), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G150), .B2(new_n763), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT108), .Z(new_n956));
  AOI22_X1  g0756(.A1(new_n751), .A2(G159), .B1(new_n754), .B2(G143), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n757), .A2(G77), .B1(new_n760), .B2(G50), .ZN(new_n958));
  INV_X1    g0758(.A(new_n745), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G58), .A2(new_n770), .B1(new_n959), .B2(G137), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n957), .A2(new_n958), .A3(new_n257), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n953), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT109), .Z(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n934), .B1(new_n942), .B2(new_n798), .C1(new_n964), .C2(new_n817), .ZN(new_n965));
  INV_X1    g0765(.A(new_n692), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n488), .B(new_n482), .C1(new_n461), .C2(new_n681), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n488), .A2(new_n681), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n679), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT45), .B1(new_n679), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT44), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n969), .B1(KEYINPUT106), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n677), .A2(new_n678), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(KEYINPUT106), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n966), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT107), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT107), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n980), .B(new_n966), .C1(new_n972), .C2(new_n977), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n675), .A2(new_n638), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n691), .B2(new_n675), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n686), .B(new_n983), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n725), .A2(new_n732), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n972), .ZN(new_n986));
  INV_X1    g0786(.A(new_n977), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n987), .A3(new_n692), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n979), .A2(new_n981), .A3(new_n985), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n733), .ZN(new_n990));
  XNOR2_X1  g0790(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n695), .B(new_n991), .Z(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n738), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n969), .A2(new_n675), .A3(new_n638), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n488), .B1(new_n967), .B2(new_n689), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n995), .A2(KEYINPUT42), .B1(new_n681), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(KEYINPUT42), .B2(new_n995), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n998), .B1(new_n999), .B2(new_n941), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT102), .Z(new_n1002));
  NOR2_X1   g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT104), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT103), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n969), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n692), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1007), .B(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n965), .B1(new_n994), .B2(new_n1011), .ZN(G387));
  NOR2_X1   g0812(.A1(new_n985), .A2(new_n696), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n984), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1013), .B1(new_n733), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n358), .A2(new_n303), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT50), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n697), .B(new_n242), .C1(new_n279), .C2(new_n260), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n784), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n224), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(G45), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n791), .A2(new_n697), .B1(G107), .B2(new_n208), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n796), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1023), .A2(new_n739), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n828), .A2(new_n948), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n819), .A2(new_n836), .B1(new_n759), .B2(new_n832), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(G322), .C2(new_n754), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1027), .A2(KEYINPUT48), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(KEYINPUT48), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n766), .A2(new_n944), .B1(new_n769), .B2(new_n602), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n757), .A2(G116), .B1(new_n959), .B2(G326), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1032), .A2(new_n381), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n769), .A2(new_n260), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n943), .A2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n279), .B2(new_n759), .C1(new_n746), .C2(new_n753), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n751), .A2(new_n358), .B1(G150), .B2(new_n959), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n303), .B2(new_n828), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n767), .A2(new_n519), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n410), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT110), .Z(new_n1044));
  AND2_X1   g0844(.A1(new_n1035), .A2(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1024), .B1(new_n691), .B2(new_n798), .C1(new_n1045), .C2(new_n817), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1015), .B(new_n1046), .C1(new_n737), .C2(new_n984), .ZN(G393));
  INV_X1    g0847(.A(KEYINPUT111), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n988), .A2(new_n978), .A3(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(KEYINPUT111), .B(new_n966), .C1(new_n972), .C2(new_n977), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n989), .B(new_n695), .C1(new_n1051), .C2(new_n985), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1008), .A2(new_n795), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n236), .A2(new_n785), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n796), .B1(new_n442), .B2(new_n208), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n739), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n758), .B1(new_n944), .B2(new_n769), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n257), .B(new_n1057), .C1(G322), .C2(new_n959), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT113), .Z(new_n1059));
  AOI22_X1  g0859(.A1(new_n763), .A2(G311), .B1(new_n754), .B2(G317), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT52), .Z(new_n1061));
  NAND2_X1  g0861(.A1(new_n767), .A2(G116), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n751), .A2(G303), .B1(G294), .B2(new_n760), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n751), .A2(G50), .B1(G87), .B2(new_n757), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n767), .A2(G77), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n410), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G68), .A2(new_n770), .B1(new_n959), .B2(G143), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n272), .B2(new_n759), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n763), .A2(G159), .B1(new_n754), .B2(G150), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1059), .A2(new_n1064), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1056), .B1(new_n1074), .B2(new_n782), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1051), .A2(new_n738), .B1(new_n1053), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1052), .A2(new_n1076), .ZN(G390));
  INV_X1    g0877(.A(KEYINPUT114), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n850), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n888), .B1(new_n845), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n886), .B2(new_n894), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n724), .A2(G330), .A3(new_n805), .A4(new_n1079), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n730), .A2(new_n681), .A3(new_n805), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n850), .B1(new_n1083), .B2(new_n844), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n906), .A2(new_n887), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1078), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1080), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1092));
  OAI211_X1 g0892(.A(G330), .B(new_n805), .C1(new_n721), .C2(new_n723), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(new_n850), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1091), .A2(KEYINPUT114), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1092), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1091), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n903), .A2(G330), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n847), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n347), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n340), .A2(new_n346), .A3(new_n847), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1102), .A2(new_n1103), .B1(new_n804), .B2(new_n803), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1087), .A2(new_n1096), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n793), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n815), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n739), .B1(new_n1109), .B2(new_n358), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT117), .Z(new_n1111));
  AOI22_X1  g0911(.A1(new_n751), .A2(G137), .B1(new_n754), .B2(G128), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n257), .C1(new_n746), .C2(new_n766), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n769), .A2(new_n274), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT53), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n757), .A2(G50), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n763), .A2(G132), .B1(new_n760), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1113), .B(new_n1120), .C1(G125), .C2(new_n775), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1122), .A2(KEYINPUT118), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n819), .A2(new_n453), .B1(new_n753), .B2(new_n944), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n828), .A2(new_n492), .B1(new_n759), .B2(new_n442), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n257), .B(new_n823), .C1(G87), .C2(new_n770), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n775), .A2(G294), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1126), .A2(new_n1066), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1122), .A2(KEYINPUT118), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1123), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1111), .B1(new_n1131), .B2(new_n782), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1107), .A2(new_n738), .B1(new_n1108), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT115), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1093), .A2(new_n850), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1105), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1083), .A2(new_n844), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n806), .A2(new_n1100), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n850), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1136), .A2(new_n845), .B1(new_n1082), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n897), .B(new_n666), .C1(new_n910), .C2(new_n1099), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1134), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1106), .B1(new_n1081), .B2(new_n1092), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1081), .A2(new_n1086), .A3(new_n1078), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT114), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1142), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n695), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT116), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1087), .A2(new_n1096), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1142), .B1(new_n1149), .B2(new_n1143), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n696), .B1(new_n1107), .B2(new_n1142), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1142), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT116), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1133), .B1(new_n1151), .B2(new_n1156), .ZN(G378));
  INV_X1    g0957(.A(KEYINPUT57), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT121), .ZN(new_n1159));
  INV_X1    g0959(.A(G330), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n881), .A2(new_n859), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT37), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n861), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT38), .B1(new_n1163), .B2(new_n876), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n889), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(KEYINPUT40), .B1(new_n1165), .B2(new_n904), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n871), .A2(new_n905), .A3(new_n913), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1160), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n288), .A2(new_n855), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n302), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1169), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1171), .B(new_n292), .C1(new_n300), .C2(new_n301), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1170), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1174), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n302), .A2(new_n1169), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n1172), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1159), .B1(new_n1168), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1179), .ZN(new_n1181));
  OAI211_X1 g0981(.A(KEYINPUT121), .B(new_n1181), .C1(new_n909), .C2(new_n1160), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(G330), .B(new_n1179), .C1(new_n915), .C2(new_n916), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(KEYINPUT122), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1168), .A2(new_n1186), .A3(new_n1179), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1183), .A2(new_n1188), .A3(new_n896), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n896), .B1(new_n1183), .B2(new_n1188), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1140), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1141), .B1(new_n1107), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1158), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1183), .A2(new_n1188), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n896), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1183), .A2(new_n1188), .A3(new_n896), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1149), .A2(new_n1143), .A3(new_n1192), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1141), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1199), .A2(new_n1202), .A3(KEYINPUT57), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1194), .A2(new_n695), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1181), .A2(new_n793), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n381), .A2(new_n239), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1206), .B(new_n303), .C1(G33), .C2(G41), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT119), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1036), .B(new_n954), .C1(G116), .C2(new_n754), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n763), .A2(G107), .B1(new_n519), .B2(new_n760), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n751), .A2(G97), .B1(G58), .B2(new_n757), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1206), .B(new_n1212), .C1(G283), .C2(new_n775), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1208), .B1(new_n1213), .B2(KEYINPUT58), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n238), .B(new_n239), .C1(new_n756), .C2(new_n746), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G124), .B2(new_n959), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n760), .A2(G137), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n763), .A2(G128), .B1(new_n754), .B2(G125), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n751), .A2(G132), .B1(new_n770), .B2(new_n1118), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n767), .A2(G150), .ZN(new_n1220));
  AND4_X1   g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT59), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1216), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1221), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1214), .B1(KEYINPUT58), .B2(new_n1213), .C1(new_n1223), .C2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n782), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT120), .Z(new_n1228));
  AOI211_X1 g1028(.A(new_n742), .B(new_n1228), .C1(new_n303), .C2(new_n815), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1205), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1191), .B2(new_n737), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1204), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(G375));
  NAND2_X1  g1034(.A1(new_n1192), .A2(new_n1201), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n993), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n739), .B1(new_n1109), .B2(G68), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1079), .A2(new_n794), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n751), .A2(G116), .B1(new_n754), .B2(G294), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n763), .A2(G283), .B1(G107), .B2(new_n760), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n837), .C2(new_n832), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G77), .A2(new_n757), .B1(new_n770), .B2(G97), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n351), .A3(new_n1041), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n775), .A2(G128), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n751), .A2(new_n1118), .B1(new_n754), .B2(G132), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n763), .A2(G137), .B1(G150), .B2(new_n760), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G58), .A2(new_n757), .B1(new_n770), .B2(G159), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n410), .C1(new_n303), .C2(new_n766), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n1242), .A2(new_n1244), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1238), .B(new_n1239), .C1(new_n782), .C2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1192), .B2(new_n738), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1237), .A2(new_n1253), .ZN(G381));
  NAND2_X1  g1054(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1133), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(G375), .A2(new_n1256), .ZN(new_n1257));
  OR3_X1    g1057(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(G387), .A2(new_n1258), .A3(G390), .A4(G381), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(G407));
  OAI21_X1  g1060(.A(new_n1257), .B1(new_n1259), .B2(new_n672), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(G213), .ZN(G409));
  INV_X1    g1062(.A(G390), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G387), .A2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(G393), .B(new_n800), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G390), .B(new_n965), .C1(new_n994), .C2(new_n1011), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1265), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(G378), .A2(new_n1204), .A3(new_n1232), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1191), .A2(new_n1193), .A3(new_n992), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1133), .B(new_n1255), .C1(new_n1272), .C2(new_n1231), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n672), .A2(G213), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1235), .A2(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1236), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n1141), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n695), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n814), .A2(KEYINPUT123), .A3(new_n840), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1280), .A2(new_n1253), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT123), .B1(new_n814), .B2(new_n840), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1283), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1279), .A2(new_n1281), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1274), .A2(new_n1275), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT62), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1271), .A2(new_n1273), .B1(G213), .B2(new_n672), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n672), .A2(G213), .A3(G2897), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1287), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1292), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1284), .A2(new_n1286), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1289), .B(new_n1290), .C1(new_n1291), .C2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT124), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1288), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1291), .A2(KEYINPUT124), .A3(new_n1287), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT62), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1270), .B1(new_n1297), .B2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1274), .A2(KEYINPUT63), .A3(new_n1275), .A4(new_n1287), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1269), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1290), .B1(new_n1291), .B2(new_n1296), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1299), .A2(new_n1307), .A3(new_n1300), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1306), .A2(KEYINPUT125), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT125), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1302), .B1(new_n1309), .B2(new_n1310), .ZN(G405));
  OAI21_X1  g1111(.A(new_n1271), .B1(new_n1233), .B2(new_n1256), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT126), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT127), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1315), .B(new_n1271), .C1(new_n1233), .C2(new_n1256), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1287), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1312), .A2(KEYINPUT126), .A3(new_n1318), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1314), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1317), .B1(new_n1314), .B2(new_n1319), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1270), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1314), .A2(new_n1319), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1317), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1314), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(new_n1269), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1322), .A2(new_n1327), .ZN(G402));
endmodule


