//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020;
  INV_X1    g000(.A(G64gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G57gat), .ZN(new_n203));
  INV_X1    g002(.A(G57gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G64gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n206), .A2(KEYINPUT9), .ZN(new_n207));
  XNOR2_X1  g006(.A(G71gat), .B(G78gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT100), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT101), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n204), .A2(KEYINPUT101), .A3(G64gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n203), .A3(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(G71gat), .A2(G78gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n213), .B(new_n208), .C1(KEYINPUT9), .C2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n208), .B1(KEYINPUT9), .B2(new_n206), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT100), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n209), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT21), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  AND2_X1   g024(.A1(G15gat), .A2(G22gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G15gat), .A2(G22gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT94), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n226), .B2(new_n227), .ZN(new_n230));
  INV_X1    g029(.A(G1gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI221_X1 g031(.A(new_n229), .B1(new_n225), .B2(G1gat), .C1(new_n226), .C2(new_n227), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT95), .B(G8gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT96), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(new_n233), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G8gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT96), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n232), .A2(new_n239), .A3(new_n233), .A4(new_n234), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n220), .B2(new_n219), .ZN(new_n242));
  INV_X1    g041(.A(G183gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G231gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n242), .B(G183gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n245), .ZN(new_n249));
  XNOR2_X1  g048(.A(G127gat), .B(G155gat), .ZN(new_n250));
  INV_X1    g049(.A(G211gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n247), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n253), .B1(new_n247), .B2(new_n249), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n224), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n248), .A2(new_n245), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n244), .A2(new_n246), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n252), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n247), .A2(new_n249), .A3(new_n253), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n223), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n263));
  INV_X1    g062(.A(G43gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(G50gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(G50gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT15), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT91), .ZN(new_n269));
  INV_X1    g068(.A(G50gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(KEYINPUT91), .A2(G50gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n264), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT15), .B1(new_n273), .B2(new_n266), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n268), .B1(new_n274), .B2(KEYINPUT92), .ZN(new_n275));
  INV_X1    g074(.A(G36gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT90), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT90), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G36gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n279), .A3(G29gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT14), .ZN(new_n281));
  OR3_X1    g080(.A1(new_n281), .A2(G29gat), .A3(G36gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n281), .B1(G29gat), .B2(G36gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n275), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT92), .ZN(new_n287));
  AOI211_X1 g086(.A(new_n287), .B(KEYINPUT15), .C1(new_n273), .C2(new_n266), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n268), .B1(new_n288), .B2(new_n284), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G85gat), .A2(G92gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT7), .ZN(new_n292));
  NAND2_X1  g091(.A1(G99gat), .A2(G106gat), .ZN(new_n293));
  INV_X1    g092(.A(G85gat), .ZN(new_n294));
  INV_X1    g093(.A(G92gat), .ZN(new_n295));
  AOI22_X1  g094(.A1(KEYINPUT8), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n296), .A2(KEYINPUT102), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(KEYINPUT102), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n292), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G99gat), .B(G106gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n300), .B(new_n292), .C1(new_n297), .C2(new_n298), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n263), .B1(new_n290), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT103), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT15), .ZN(new_n309));
  INV_X1    g108(.A(new_n272), .ZN(new_n310));
  NOR2_X1   g109(.A1(KEYINPUT91), .A2(G50gat), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n310), .A2(new_n311), .A3(G43gat), .ZN(new_n312));
  OAI211_X1 g111(.A(KEYINPUT92), .B(new_n309), .C1(new_n312), .C2(new_n265), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n285), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n268), .A2(new_n314), .B1(new_n275), .B2(new_n285), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT93), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT17), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND4_X1   g116(.A1(new_n316), .A2(new_n286), .A3(new_n289), .A4(KEYINPUT17), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n304), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n306), .A2(new_n308), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n308), .B1(new_n306), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT104), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT103), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n305), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n319), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n307), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT104), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(new_n320), .ZN(new_n329));
  XNOR2_X1  g128(.A(G190gat), .B(G218gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G134gat), .B(G162gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  NAND3_X1  g131(.A1(new_n323), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n332), .B1(new_n323), .B2(new_n329), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n262), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT105), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n323), .A2(new_n329), .ZN(new_n338));
  INV_X1    g137(.A(new_n332), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n333), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT105), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(new_n262), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT10), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n304), .A2(new_n219), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n345), .B2(KEYINPUT106), .ZN(new_n346));
  NAND2_X1  g145(.A1(G230gat), .A2(G233gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n304), .A2(new_n219), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT106), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n349), .B(KEYINPUT10), .C1(new_n304), .C2(new_n219), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n346), .A2(new_n347), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n209), .A2(new_n218), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n352), .A2(new_n215), .A3(new_n303), .A4(new_n302), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n347), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G120gat), .B(G148gat), .ZN(new_n357));
  INV_X1    g156(.A(G176gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G204gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n351), .A2(new_n356), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT107), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT107), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n351), .A2(new_n365), .A3(new_n356), .A4(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n356), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n361), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n337), .A2(new_n343), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(new_n202), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(new_n295), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT74), .B(G204gat), .ZN(new_n378));
  INV_X1    g177(.A(G197gat), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT22), .ZN(new_n381));
  INV_X1    g180(.A(G218gat), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n251), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n379), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G211gat), .B(G218gat), .Z(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT75), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n385), .B(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT65), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT24), .ZN(new_n392));
  INV_X1    g191(.A(G190gat), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n243), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n243), .A2(new_n393), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT67), .B1(new_n397), .B2(KEYINPUT23), .ZN(new_n398));
  NAND2_X1  g197(.A1(G169gat), .A2(G176gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n397), .A2(KEYINPUT67), .A3(KEYINPUT23), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT66), .B(G169gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(KEYINPUT23), .A3(new_n358), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n396), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(KEYINPUT69), .B(G190gat), .Z(new_n408));
  XOR2_X1   g207(.A(KEYINPUT68), .B(G183gat), .Z(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT70), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT70), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT69), .B(G190gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT68), .B(G183gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n410), .A2(new_n414), .A3(new_n394), .A4(new_n390), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT25), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n397), .B2(KEYINPUT23), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n402), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n407), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n397), .A2(KEYINPUT26), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n399), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n397), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT71), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT27), .B(G183gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n408), .A2(KEYINPUT28), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(new_n413), .B2(KEYINPUT27), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n412), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n426), .B1(new_n429), .B2(KEYINPUT28), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n419), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT76), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT76), .A3(new_n431), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(G226gat), .A2(G233gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(KEYINPUT29), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n389), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n434), .A2(new_n435), .A3(new_n439), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n431), .A3(new_n437), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n442), .A2(new_n389), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n377), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n389), .A3(new_n443), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n436), .A2(new_n437), .B1(new_n432), .B2(new_n439), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n446), .B(new_n376), .C1(new_n447), .C2(new_n389), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n448), .A3(KEYINPUT30), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n450), .B(new_n377), .C1(new_n441), .C2(new_n444), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G141gat), .B(G148gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT78), .ZN(new_n455));
  NAND2_X1  g254(.A1(G155gat), .A2(G162gat), .ZN(new_n456));
  INV_X1    g255(.A(G155gat), .ZN(new_n457));
  INV_X1    g256(.A(G162gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n456), .B1(new_n459), .B2(KEYINPUT2), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT77), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n454), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G141gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(G148gat), .ZN(new_n465));
  INV_X1    g264(.A(G148gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(G141gat), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT77), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT2), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n463), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n459), .A2(new_n456), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT81), .B(KEYINPUT3), .Z(new_n473));
  NAND3_X1  g272(.A1(new_n461), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT82), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n460), .A2(new_n455), .B1(new_n470), .B2(new_n471), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n473), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n476), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT79), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT3), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n476), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT80), .ZN(new_n485));
  XNOR2_X1  g284(.A(G113gat), .B(G120gat), .ZN(new_n486));
  OAI21_X1  g285(.A(G127gat), .B1(new_n486), .B2(KEYINPUT1), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT1), .ZN(new_n488));
  INV_X1    g287(.A(G127gat), .ZN(new_n489));
  INV_X1    g288(.A(G113gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(G120gat), .ZN(new_n491));
  INV_X1    g290(.A(G120gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(G113gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n488), .B(new_n489), .C1(new_n491), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n487), .A2(G134gat), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(G134gat), .B1(new_n487), .B2(new_n494), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n485), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n497), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(KEYINPUT80), .A3(new_n495), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n479), .A2(new_n481), .A3(new_n484), .A4(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n496), .A2(new_n497), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n476), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT4), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n506), .A3(new_n476), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G225gat), .A2(G233gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT83), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n505), .A2(new_n515), .A3(new_n507), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n504), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n502), .A2(new_n511), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n480), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n504), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n521), .B2(new_n512), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT84), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n518), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n523), .B1(new_n518), .B2(new_n522), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n514), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT0), .B(G57gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G85gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(G1gat), .B(G29gat), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n529), .B(new_n530), .Z(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n527), .A2(KEYINPUT6), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n522), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT84), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n535), .A2(new_n524), .B1(new_n510), .B2(new_n513), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n536), .A2(new_n531), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n531), .B(new_n514), .C1(new_n525), .C2(new_n526), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n533), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n453), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G22gat), .B(G50gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G78gat), .B(G106gat), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT31), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n477), .B1(new_n476), .B2(new_n473), .ZN(new_n549));
  AND4_X1   g348(.A1(new_n477), .A2(new_n461), .A3(new_n472), .A4(new_n473), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT29), .B1(new_n475), .B2(new_n478), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT87), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n555), .A3(new_n388), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n389), .A2(new_n548), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n476), .B1(new_n557), .B2(new_n483), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G228gat), .A2(G233gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n386), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n385), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n380), .A2(new_n386), .A3(new_n383), .A4(new_n384), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n548), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT85), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT85), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n565), .A2(new_n569), .A3(new_n548), .A4(new_n566), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n473), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n562), .B1(new_n571), .B2(new_n480), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT86), .B1(new_n554), .B2(new_n389), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n551), .A2(new_n574), .A3(new_n388), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n547), .B1(new_n563), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n561), .B1(new_n556), .B2(new_n559), .ZN(new_n578));
  INV_X1    g377(.A(new_n576), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n578), .A2(new_n579), .A3(new_n546), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n544), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n547), .A3(new_n576), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n546), .B1(new_n578), .B2(new_n579), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n543), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT73), .B(G71gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G99gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(G15gat), .B(G43gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G227gat), .ZN(new_n592));
  INV_X1    g391(.A(G233gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n419), .A2(new_n503), .A3(new_n431), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n503), .B1(new_n419), .B2(new_n431), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT33), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n591), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n594), .ZN(new_n601));
  INV_X1    g400(.A(new_n503), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n432), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n603), .B2(new_n595), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT32), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT72), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT72), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n598), .A2(new_n607), .A3(KEYINPUT32), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n600), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT34), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n598), .B(KEYINPUT32), .C1(new_n599), .C2(new_n591), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n609), .B2(new_n611), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n596), .A2(new_n597), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n601), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n609), .A2(new_n611), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT34), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n587), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n615), .B1(new_n612), .B2(new_n613), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n617), .A3(new_n620), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT36), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n542), .A2(new_n586), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n520), .A2(new_n511), .A3(new_n504), .ZN(new_n627));
  OAI211_X1 g426(.A(KEYINPUT39), .B(new_n627), .C1(new_n510), .C2(new_n511), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n531), .B(KEYINPUT88), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n511), .B1(new_n502), .B2(new_n508), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(KEYINPUT40), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n628), .A2(new_n633), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n527), .A2(new_n630), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n452), .A2(KEYINPUT89), .A3(new_n634), .A4(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n445), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n441), .B2(new_n444), .ZN(new_n641));
  OAI211_X1 g440(.A(KEYINPUT37), .B(new_n446), .C1(new_n447), .C2(new_n389), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n642), .A3(new_n376), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n639), .B1(new_n643), .B2(KEYINPUT38), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n538), .B(new_n539), .C1(new_n536), .C2(new_n629), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n447), .A2(new_n389), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n442), .A2(new_n443), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n646), .B(KEYINPUT37), .C1(new_n647), .C2(new_n389), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n648), .A2(new_n641), .A3(new_n649), .A4(new_n376), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n644), .A2(new_n645), .A3(new_n533), .A4(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT89), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n449), .A2(new_n451), .A3(new_n634), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n636), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n536), .B2(new_n629), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n652), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n638), .A2(new_n651), .A3(new_n656), .A4(new_n585), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n585), .A2(new_n624), .A3(new_n623), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT35), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n645), .A2(new_n533), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n453), .A4(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n585), .A2(new_n624), .A3(new_n623), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT35), .B1(new_n542), .B2(new_n662), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n626), .A2(new_n657), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n241), .B1(new_n317), .B2(new_n318), .ZN(new_n665));
  NAND2_X1  g464(.A1(G229gat), .A2(G233gat), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n315), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n666), .B(KEYINPUT13), .Z(new_n673));
  NOR2_X1   g472(.A1(new_n315), .A2(new_n667), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n668), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT97), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT97), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n677), .B(new_n673), .C1(new_n668), .C2(new_n674), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n665), .A2(KEYINPUT18), .A3(new_n666), .A4(new_n669), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n672), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT11), .B(G169gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G197gat), .ZN(new_n683));
  XOR2_X1   g482(.A(G113gat), .B(G141gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT12), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n672), .A2(new_n679), .A3(new_n686), .A4(new_n680), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n688), .B2(new_n690), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n664), .A2(KEYINPUT99), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT99), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n661), .A2(new_n663), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n542), .A2(new_n586), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n622), .A2(new_n625), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n657), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n696), .B1(new_n701), .B2(new_n693), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n373), .B1(new_n695), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT99), .B1(new_n664), .B2(new_n694), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n701), .A2(new_n696), .A3(new_n693), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(KEYINPUT108), .A3(new_n373), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n541), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g512(.A(KEYINPUT16), .B(G8gat), .Z(new_n714));
  NAND4_X1  g513(.A1(new_n710), .A2(KEYINPUT42), .A3(new_n452), .A4(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT108), .B1(new_n708), .B2(new_n373), .ZN(new_n717));
  AOI211_X1 g516(.A(new_n704), .B(new_n372), .C1(new_n706), .C2(new_n707), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n452), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n716), .B1(new_n719), .B2(G8gat), .ZN(new_n720));
  INV_X1    g519(.A(new_n714), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n715), .B1(new_n720), .B2(new_n722), .ZN(G1325gat));
  NOR2_X1   g522(.A1(new_n616), .A2(new_n621), .ZN(new_n724));
  AOI21_X1  g523(.A(G15gat), .B1(new_n710), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n699), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n710), .A2(G15gat), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(G1326gat));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n586), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT43), .B(G22gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1327gat));
  INV_X1    g530(.A(new_n341), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n262), .A2(new_n370), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n708), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(G29gat), .A3(new_n541), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT45), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n664), .B2(new_n341), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n341), .B1(new_n697), .B2(new_n700), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT44), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n688), .A2(new_n690), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n739), .A2(new_n741), .A3(new_n742), .A4(new_n733), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n743), .A2(new_n541), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n737), .B1(new_n744), .B2(G29gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n736), .B1(new_n745), .B2(new_n735), .ZN(G1328gat));
  AND2_X1   g545(.A1(new_n708), .A2(new_n733), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n277), .A2(new_n279), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n453), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n747), .A2(new_n748), .A3(new_n732), .A4(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n751), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT46), .B1(new_n734), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n750), .B1(new_n743), .B2(new_n453), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n752), .A2(new_n754), .A3(KEYINPUT109), .A4(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1329gat));
  OR3_X1    g559(.A1(new_n743), .A2(new_n264), .A3(new_n699), .ZN(new_n761));
  INV_X1    g560(.A(new_n724), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n264), .B1(new_n734), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT47), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1330gat));
  NOR2_X1   g567(.A1(new_n310), .A2(new_n311), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n747), .A2(new_n586), .A3(new_n770), .A4(new_n732), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n743), .B2(new_n585), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1331gat));
  NAND2_X1  g575(.A1(new_n337), .A2(new_n343), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n664), .A2(new_n777), .A3(new_n371), .ZN(new_n778));
  INV_X1    g577(.A(new_n742), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n711), .A2(KEYINPUT110), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n711), .A2(KEYINPUT110), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(new_n204), .ZN(G1332gat));
  NOR2_X1   g586(.A1(new_n780), .A2(new_n453), .ZN(new_n788));
  NOR2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  AND2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n788), .B2(new_n789), .ZN(G1333gat));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793));
  INV_X1    g592(.A(G71gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n780), .B2(new_n762), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n778), .A2(G71gat), .A3(new_n726), .A4(new_n779), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n796), .B1(new_n795), .B2(new_n797), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n793), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n800), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(KEYINPUT50), .A3(new_n798), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1334gat));
  NOR2_X1   g603(.A1(new_n780), .A2(new_n585), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(G78gat), .Z(G1335gat));
  AOI21_X1  g605(.A(KEYINPUT44), .B1(new_n701), .B2(new_n732), .ZN(new_n807));
  AOI211_X1 g606(.A(new_n738), .B(new_n341), .C1(new_n697), .C2(new_n700), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n262), .A2(new_n742), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n370), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT112), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n739), .A2(new_n741), .A3(new_n812), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n294), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n740), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT51), .B1(new_n740), .B2(new_n810), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n711), .A3(new_n370), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n819), .A2(new_n711), .B1(new_n294), .B2(new_n825), .ZN(G1336gat));
  OAI21_X1  g625(.A(G92gat), .B1(new_n815), .B2(new_n453), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n452), .A2(new_n295), .A3(new_n370), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT113), .Z(new_n830));
  OAI211_X1 g629(.A(new_n827), .B(new_n828), .C1(new_n823), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n823), .A2(new_n830), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n452), .B1(new_n813), .B2(new_n817), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(G92gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n831), .B1(new_n834), .B2(new_n828), .ZN(G1337gat));
  INV_X1    g634(.A(G99gat), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n814), .B2(new_n818), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n824), .A2(new_n724), .A3(new_n370), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n837), .A2(new_n726), .B1(new_n836), .B2(new_n838), .ZN(G1338gat));
  XNOR2_X1  g638(.A(KEYINPUT114), .B(G106gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n840), .B1(new_n815), .B2(new_n585), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842));
  INV_X1    g641(.A(G106gat), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n843), .B(new_n370), .C1(new_n821), .C2(new_n822), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n841), .B(new_n842), .C1(new_n844), .C2(new_n585), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n585), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n586), .B1(new_n813), .B2(new_n817), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n840), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n845), .B1(new_n848), .B2(new_n842), .ZN(G1339gat));
  AND4_X1   g648(.A1(new_n779), .A2(new_n337), .A3(new_n343), .A4(new_n371), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n350), .A2(new_n348), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT10), .B1(new_n353), .B2(new_n349), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n355), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n855), .A2(new_n351), .A3(KEYINPUT54), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n361), .B1(new_n351), .B2(KEYINPUT54), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n351), .A2(KEYINPUT54), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n855), .A2(new_n351), .A3(KEYINPUT54), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT55), .A4(new_n361), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n367), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n666), .B1(new_n665), .B2(new_n669), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n668), .A2(new_n674), .A3(new_n673), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n685), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n690), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n732), .A2(new_n863), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n370), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n779), .B2(new_n862), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n341), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n262), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n851), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n658), .A3(new_n784), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n875), .A2(KEYINPUT115), .A3(new_n658), .A4(new_n784), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n453), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n490), .A3(new_n742), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n662), .A2(new_n541), .A3(new_n452), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G113gat), .B1(new_n886), .B2(new_n694), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(G1340gat));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n492), .A3(new_n370), .ZN(new_n889));
  OAI21_X1  g688(.A(G120gat), .B1(new_n886), .B2(new_n371), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1341gat));
  NAND4_X1  g690(.A1(new_n878), .A2(new_n453), .A3(new_n262), .A4(new_n879), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n489), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n885), .A2(G127gat), .A3(new_n262), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT116), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n896), .A2(new_n898), .ZN(G1342gat));
  OR2_X1    g698(.A1(new_n341), .A2(G134gat), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n881), .A2(KEYINPUT56), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G134gat), .B1(new_n886), .B2(new_n341), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT56), .B1(new_n881), .B2(new_n900), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G1343gat));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n585), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n691), .A2(new_n692), .A3(new_n862), .ZN(new_n907));
  INV_X1    g706(.A(new_n870), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT118), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n692), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n863), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n870), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n909), .A2(new_n341), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n262), .B1(new_n915), .B2(new_n869), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n906), .B1(new_n916), .B2(new_n850), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n586), .B1(new_n850), .B2(new_n873), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n905), .ZN(new_n921));
  OAI211_X1 g720(.A(KEYINPUT119), .B(new_n906), .C1(new_n916), .C2(new_n850), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n726), .A2(new_n541), .A3(new_n452), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n464), .B1(new_n925), .B2(new_n742), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n785), .B1(new_n874), .B2(new_n851), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n726), .A2(new_n585), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n453), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n693), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(G141gat), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT58), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n923), .A2(new_n693), .A3(new_n924), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT58), .B1(new_n934), .B2(G141gat), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT120), .B1(new_n931), .B2(G141gat), .ZN(new_n936));
  OR4_X1    g735(.A1(KEYINPUT120), .A2(new_n929), .A3(G141gat), .A4(new_n694), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n933), .A2(new_n938), .ZN(G1344gat));
  NOR2_X1   g738(.A1(new_n372), .A2(new_n693), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n905), .B(new_n586), .C1(new_n916), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n920), .A2(KEYINPUT57), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n941), .A2(new_n942), .A3(new_n924), .A4(new_n370), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G148gat), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n943), .A2(new_n944), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT59), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n923), .A2(new_n370), .A3(new_n924), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n466), .A2(KEYINPUT59), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n948), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n930), .A2(new_n466), .A3(new_n370), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1345gat));
  NAND3_X1  g755(.A1(new_n925), .A2(G155gat), .A3(new_n262), .ZN(new_n957));
  INV_X1    g756(.A(new_n262), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n457), .B1(new_n929), .B2(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n957), .A2(new_n959), .ZN(G1346gat));
  NAND3_X1  g759(.A1(new_n925), .A2(G162gat), .A3(new_n732), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n458), .B1(new_n929), .B2(new_n341), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(G1347gat));
  AOI21_X1  g762(.A(new_n711), .B1(new_n851), .B2(new_n874), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n662), .A2(new_n453), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(new_n403), .A3(new_n742), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n966), .A2(KEYINPUT123), .A3(new_n403), .A4(new_n742), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n452), .B(new_n724), .C1(new_n782), .C2(new_n783), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n972), .A2(KEYINPUT124), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n586), .B1(new_n972), .B2(KEYINPUT124), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n973), .A2(new_n875), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(G169gat), .B1(new_n975), .B2(new_n694), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n971), .A2(KEYINPUT125), .A3(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1348gat));
  NOR3_X1   g780(.A1(new_n975), .A2(new_n358), .A3(new_n371), .ZN(new_n982));
  AOI21_X1  g781(.A(G176gat), .B1(new_n966), .B2(new_n370), .ZN(new_n983));
  OR2_X1    g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(G1349gat));
  INV_X1    g784(.A(new_n975), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n986), .A2(KEYINPUT126), .A3(new_n262), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n988), .B1(new_n975), .B2(new_n958), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n987), .A2(new_n413), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n966), .A2(new_n425), .A3(new_n262), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(KEYINPUT60), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT60), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n990), .A2(new_n994), .A3(new_n991), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(new_n995), .ZN(G1350gat));
  OAI21_X1  g795(.A(G190gat), .B1(new_n975), .B2(new_n341), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT61), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n966), .A2(new_n408), .A3(new_n732), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1351gat));
  NAND3_X1  g799(.A1(new_n964), .A2(new_n452), .A3(new_n928), .ZN(new_n1001));
  INV_X1    g800(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n1002), .A2(new_n379), .A3(new_n742), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n941), .A2(new_n942), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n785), .A2(new_n452), .A3(new_n699), .ZN(new_n1005));
  NOR3_X1   g804(.A1(new_n1004), .A2(new_n694), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1003), .B1(new_n1006), .B2(new_n379), .ZN(G1352gat));
  NAND2_X1  g806(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n1002), .A2(new_n360), .A3(new_n370), .A4(new_n1008), .ZN(new_n1009));
  NOR2_X1   g808(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NOR3_X1   g810(.A1(new_n1004), .A2(new_n371), .A3(new_n1005), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1011), .B1(new_n360), .B2(new_n1012), .ZN(G1353gat));
  NAND3_X1  g812(.A1(new_n1002), .A2(new_n251), .A3(new_n262), .ZN(new_n1014));
  OR3_X1    g813(.A1(new_n1004), .A2(new_n958), .A3(new_n1005), .ZN(new_n1015));
  AND3_X1   g814(.A1(new_n1015), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1016));
  AOI21_X1  g815(.A(KEYINPUT63), .B1(new_n1015), .B2(G211gat), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(G1354gat));
  NAND3_X1  g817(.A1(new_n1002), .A2(new_n382), .A3(new_n732), .ZN(new_n1019));
  NOR3_X1   g818(.A1(new_n1004), .A2(new_n341), .A3(new_n1005), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1019), .B1(new_n1020), .B2(new_n382), .ZN(G1355gat));
endmodule


