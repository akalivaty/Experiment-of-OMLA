//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT72), .B(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G210), .A3(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(G101), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT28), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G137), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n198), .B1(new_n196), .B2(G137), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G134), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT67), .B1(new_n203), .B2(new_n198), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n205), .B1(new_n203), .B2(KEYINPUT67), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n197), .B(new_n201), .C1(new_n204), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G131), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n196), .A2(G137), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT11), .B1(new_n209), .B2(new_n200), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n199), .A2(new_n200), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT68), .B(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n212), .A2(new_n197), .A3(new_n201), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT0), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT64), .B(G146), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n218), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g042(.A(G143), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n229), .A2(new_n230), .A3(new_n218), .A4(new_n221), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n220), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n226), .A2(G146), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n223), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n216), .A2(G143), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n221), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n225), .A2(new_n231), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n215), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n197), .A2(new_n203), .A3(KEYINPUT69), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n240), .B(G131), .C1(KEYINPUT69), .C2(new_n203), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n222), .B2(new_n223), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n243), .A2(G128), .B1(new_n236), .B2(new_n235), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n223), .B1(new_n233), .B2(new_n234), .ZN(new_n245));
  NOR4_X1   g059(.A1(new_n245), .A2(new_n242), .A3(new_n220), .A4(new_n217), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n214), .B(new_n241), .C1(new_n244), .C2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n239), .A2(KEYINPUT73), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n249));
  INV_X1    g063(.A(G116), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(G119), .ZN(new_n251));
  INV_X1    g065(.A(G119), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT71), .A3(G116), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n251), .B(new_n253), .C1(G116), .C2(new_n252), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n248), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT73), .B1(new_n239), .B2(new_n247), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n195), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n239), .A2(new_n247), .A3(new_n257), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n257), .B1(new_n239), .B2(new_n247), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT28), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n194), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n239), .A2(new_n266), .A3(new_n247), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n239), .B2(new_n247), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n256), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n269), .A2(new_n261), .A3(new_n194), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n187), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT74), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n273), .B(new_n187), .C1(new_n265), .C2(new_n270), .ZN(new_n274));
  INV_X1    g088(.A(new_n260), .ZN(new_n275));
  INV_X1    g089(.A(new_n264), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n194), .A2(new_n187), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n272), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G472), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n269), .A2(new_n261), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT31), .B1(new_n282), .B2(new_n194), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n269), .A2(new_n284), .A3(new_n261), .A4(new_n193), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n283), .B(new_n285), .C1(new_n277), .C2(new_n193), .ZN(new_n286));
  NOR2_X1   g100(.A1(G472), .A2(G902), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n286), .A2(KEYINPUT75), .A3(KEYINPUT32), .A4(new_n287), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n287), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n281), .A2(new_n290), .A3(new_n291), .A4(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT83), .ZN(new_n296));
  INV_X1    g110(.A(G140), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G125), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT78), .B1(new_n298), .B2(KEYINPUT16), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n300));
  INV_X1    g114(.A(G125), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(G140), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT76), .B(G140), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(new_n301), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(G140), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n297), .A2(KEYINPUT76), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n300), .B(G125), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n299), .B1(new_n309), .B2(KEYINPUT16), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT16), .ZN(new_n311));
  AOI211_X1 g125(.A(KEYINPUT78), .B(new_n311), .C1(new_n304), .C2(new_n308), .ZN(new_n312));
  OAI21_X1  g126(.A(G146), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n301), .A2(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT77), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n297), .A2(KEYINPUT76), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n305), .A2(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n316), .B1(new_n319), .B2(G125), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n303), .A2(KEYINPUT77), .A3(new_n301), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n314), .B(KEYINPUT16), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n311), .B1(new_n304), .B2(new_n308), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n322), .B(new_n216), .C1(new_n323), .C2(new_n299), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n313), .A2(KEYINPUT79), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n252), .A2(G128), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n252), .A2(G128), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT24), .B(G110), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n332), .B(G146), .C1(new_n310), .C2(new_n312), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(KEYINPUT23), .ZN(new_n334));
  MUX2_X1   g148(.A(new_n334), .B(KEYINPUT23), .S(new_n328), .Z(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G110), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n325), .A2(new_n331), .A3(new_n333), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n315), .A2(new_n298), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(new_n222), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n329), .A2(new_n330), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n335), .B2(G110), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n313), .B(new_n343), .C1(new_n342), .C2(new_n341), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n337), .A2(KEYINPUT81), .A3(new_n344), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT82), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT22), .B(G137), .Z(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n296), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n337), .A2(KEYINPUT81), .A3(new_n344), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT81), .B1(new_n337), .B2(new_n344), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n296), .B(new_n353), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n360));
  INV_X1    g174(.A(G902), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n345), .A2(new_n353), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G217), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(G234), .B2(new_n361), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT83), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n367), .A2(new_n361), .A3(new_n362), .A4(new_n357), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT25), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n365), .A2(G902), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n367), .A2(new_n362), .A3(new_n357), .A4(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n295), .A2(new_n370), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT85), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n295), .A2(new_n370), .A3(new_n377), .A4(new_n374), .ZN(new_n378));
  NOR2_X1   g192(.A1(G475), .A2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n325), .A2(new_n333), .ZN(new_n381));
  AND2_X1   g195(.A1(KEYINPUT72), .A2(G237), .ZN(new_n382));
  NOR2_X1   g196(.A1(KEYINPUT72), .A2(G237), .ZN(new_n383));
  OAI211_X1 g197(.A(G214), .B(new_n189), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n223), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n188), .A2(G143), .A3(G214), .A4(new_n189), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n213), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n387), .A2(KEYINPUT17), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n385), .A2(new_n386), .A3(new_n213), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(new_n387), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT17), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT97), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT97), .ZN(new_n394));
  NOR4_X1   g208(.A1(new_n390), .A2(new_n387), .A3(new_n394), .A4(KEYINPUT17), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n381), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G113), .B(G122), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT95), .B(G104), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n385), .A2(new_n386), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n304), .A2(G146), .A3(new_n308), .ZN(new_n404));
  INV_X1    g218(.A(new_n339), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT93), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT93), .B1(new_n404), .B2(new_n405), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n397), .A2(new_n400), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n391), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT19), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n414));
  OAI22_X1  g228(.A1(new_n309), .A2(new_n413), .B1(new_n338), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n313), .B(new_n412), .C1(new_n222), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n410), .ZN(new_n417));
  INV_X1    g231(.A(new_n400), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT96), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT96), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n421), .A3(new_n418), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n411), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT98), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT98), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n411), .A2(new_n420), .A3(new_n425), .A4(new_n422), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n380), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n397), .A2(new_n410), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n418), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n411), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n361), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n427), .A2(KEYINPUT20), .B1(G475), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G128), .B(G143), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n196), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n250), .A2(KEYINPUT14), .A3(G122), .ZN(new_n435));
  XNOR2_X1  g249(.A(G116), .B(G122), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(G107), .B(new_n435), .C1(new_n437), .C2(KEYINPUT14), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n434), .B(new_n438), .C1(G107), .C2(new_n437), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(KEYINPUT13), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n223), .A2(G128), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n440), .B(G134), .C1(KEYINPUT13), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G107), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n436), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n433), .A2(new_n196), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT9), .B(G234), .Z(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(G217), .A3(new_n189), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n447), .B(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n361), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n451), .A2(KEYINPUT99), .ZN(new_n452));
  INV_X1    g266(.A(G478), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(KEYINPUT15), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n451), .B(KEYINPUT99), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n189), .A2(G952), .ZN(new_n458));
  NAND2_X1  g272(.A1(G234), .A2(G237), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(G898), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT100), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n459), .A2(G902), .A3(G953), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n423), .A2(new_n379), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n432), .A2(new_n457), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G104), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT87), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G104), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n474), .A3(new_n443), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n474), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G107), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n443), .A3(G104), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT88), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n482), .A2(new_n479), .A3(new_n443), .A4(G104), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n476), .A2(new_n478), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G101), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n481), .A2(new_n483), .ZN(new_n486));
  INV_X1    g300(.A(G101), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n476), .A4(new_n478), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(KEYINPUT4), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n484), .A2(new_n490), .A3(G101), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n256), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n475), .B1(G104), .B2(new_n443), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G101), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT5), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n252), .A3(G116), .ZN(new_n497));
  OAI211_X1 g311(.A(G113), .B(new_n497), .C1(new_n254), .C2(new_n496), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n255), .B2(new_n254), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g315(.A(G110), .B(G122), .Z(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n502), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n492), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(KEYINPUT6), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n244), .A2(new_n246), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n301), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n301), .B2(new_n238), .ZN(new_n509));
  INV_X1    g323(.A(G224), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(G953), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n509), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n501), .A2(new_n513), .A3(new_n502), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n506), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n516));
  OR3_X1    g330(.A1(new_n509), .A2(new_n516), .A3(new_n511), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n509), .B1(new_n516), .B2(new_n511), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n495), .B(new_n499), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n502), .B(KEYINPUT8), .Z(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(new_n518), .A3(new_n521), .A4(new_n505), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n515), .A2(new_n361), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(G210), .B1(G237), .B2(G902), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT91), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n525), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n515), .A2(new_n361), .A3(new_n527), .A4(new_n522), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G214), .B1(G237), .B2(G902), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n530), .B(KEYINPUT90), .Z(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT92), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n534));
  AOI211_X1 g348(.A(new_n534), .B(new_n531), .C1(new_n526), .C2(new_n528), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT70), .B(KEYINPUT1), .Z(new_n537));
  NAND4_X1  g351(.A1(new_n229), .A2(G128), .A3(new_n218), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G128), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n245), .B2(new_n217), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n488), .A2(new_n542), .A3(new_n494), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT89), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n488), .A2(new_n542), .A3(new_n545), .A4(new_n494), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n495), .A2(new_n507), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(KEYINPUT12), .A3(new_n215), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n544), .A2(new_n546), .B1(new_n507), .B2(new_n495), .ZN(new_n552));
  INV_X1    g366(.A(new_n215), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT10), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n495), .A2(new_n507), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n547), .B2(new_n556), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n489), .A2(new_n238), .A3(new_n491), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(new_n553), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(G110), .B(G140), .ZN(new_n562));
  INV_X1    g376(.A(G227), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(G953), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n562), .B(new_n564), .Z(new_n565));
  NAND3_X1  g379(.A1(new_n555), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n565), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n553), .B1(new_n558), .B2(new_n560), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT10), .B1(new_n544), .B2(new_n546), .ZN(new_n569));
  NOR4_X1   g383(.A1(new_n569), .A2(new_n559), .A3(new_n215), .A4(new_n557), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n567), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G469), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(new_n361), .ZN(new_n574));
  NAND2_X1  g388(.A1(G469), .A2(G902), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n570), .B1(new_n550), .B2(new_n554), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n565), .B(KEYINPUT86), .Z(new_n577));
  NAND2_X1  g391(.A1(new_n561), .A2(new_n565), .ZN(new_n578));
  OAI22_X1  g392(.A1(new_n576), .A2(new_n577), .B1(new_n568), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n574), .B(new_n575), .C1(new_n573), .C2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n448), .ZN(new_n581));
  OAI21_X1  g395(.A(G221), .B1(new_n581), .B2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n470), .A2(new_n536), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n376), .A2(new_n378), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  AND2_X1   g400(.A1(new_n580), .A2(new_n582), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n286), .A2(new_n361), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G472), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n589), .A2(new_n288), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n587), .A2(new_n370), .A3(new_n374), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI211_X1 g406(.A(KEYINPUT96), .B(new_n400), .C1(new_n416), .C2(new_n410), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n388), .B1(new_n325), .B2(new_n333), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n408), .A2(new_n409), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n594), .A2(new_n396), .B1(new_n595), .B2(new_n403), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n593), .B1(new_n596), .B2(new_n400), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n425), .B1(new_n597), .B2(new_n420), .ZN(new_n598));
  INV_X1    g412(.A(new_n426), .ZN(new_n599));
  OAI211_X1 g413(.A(KEYINPUT20), .B(new_n379), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n431), .A2(G475), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n469), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT102), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(KEYINPUT102), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n450), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n450), .B2(new_n605), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(G478), .A3(new_n361), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n451), .A2(new_n453), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n602), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n465), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n524), .A2(KEYINPUT101), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n523), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n515), .A2(new_n361), .A3(new_n522), .A4(new_n614), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n524), .A2(KEYINPUT101), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n531), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n592), .A2(new_n613), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  OR2_X1    g438(.A1(new_n427), .A2(KEYINPUT20), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n432), .ZN(new_n626));
  INV_X1    g440(.A(new_n621), .ZN(new_n627));
  NOR4_X1   g441(.A1(new_n626), .A2(new_n627), .A3(new_n457), .A4(new_n465), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n592), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n349), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n371), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n370), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n584), .A2(new_n590), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  AND2_X1   g452(.A1(new_n295), .A2(new_n587), .ZN(new_n639));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n460), .B1(new_n464), .B2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n626), .A2(new_n457), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n639), .A2(new_n642), .A3(new_n621), .A4(new_n635), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  AND2_X1   g458(.A1(new_n294), .A2(new_n291), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n282), .A2(new_n193), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n262), .A2(new_n263), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n646), .B(new_n361), .C1(new_n647), .C2(new_n193), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G472), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n645), .A2(new_n290), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n457), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n529), .B(KEYINPUT38), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n650), .A2(new_n651), .A3(new_n602), .A4(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n653), .A2(new_n531), .A3(new_n635), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT103), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n641), .B(KEYINPUT39), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n583), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT40), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  NOR2_X1   g474(.A1(new_n612), .A2(new_n641), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n639), .A2(new_n621), .A3(new_n635), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G146), .ZN(G48));
  AOI21_X1  g477(.A(new_n573), .B1(new_n572), .B2(new_n361), .ZN(new_n664));
  AOI211_X1 g478(.A(G469), .B(G902), .C1(new_n566), .C2(new_n571), .ZN(new_n665));
  INV_X1    g479(.A(new_n582), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n621), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n281), .A2(new_n290), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n668), .B1(new_n669), .B2(new_n645), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n370), .A2(new_n374), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n671), .A3(new_n613), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NAND3_X1  g488(.A1(new_n628), .A2(new_n671), .A3(new_n670), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G116), .ZN(G18));
  NAND4_X1  g490(.A1(new_n600), .A2(new_n466), .A3(new_n469), .A4(new_n601), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n651), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n664), .A2(new_n665), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n621), .A2(new_n582), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n635), .A2(new_n295), .A3(new_n678), .A4(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n670), .A2(KEYINPUT104), .A3(new_n678), .A4(new_n635), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G119), .ZN(G21));
  NAND2_X1  g500(.A1(new_n602), .A2(new_n651), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n668), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT105), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n260), .B2(new_n264), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n689), .A2(new_n193), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n283), .A2(new_n285), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n287), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n589), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n671), .A2(new_n688), .A3(new_n466), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  AOI21_X1  g512(.A(new_n695), .B1(new_n370), .B2(new_n634), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n661), .A3(new_n680), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G125), .ZN(G27));
  INV_X1    g515(.A(new_n641), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n529), .A2(new_n531), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n602), .A2(new_n611), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n575), .B(KEYINPUT106), .Z(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n574), .B(new_n706), .C1(new_n573), .C2(new_n579), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n582), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n281), .A2(new_n290), .A3(new_n292), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n370), .A3(new_n374), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT42), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n375), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n612), .A2(KEYINPUT42), .A3(new_n641), .ZN(new_n714));
  INV_X1    g528(.A(new_n708), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n713), .A2(new_n714), .A3(new_n715), .A4(new_n703), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n717), .B(G131), .Z(G33));
  NAND4_X1  g532(.A1(new_n713), .A2(new_n642), .A3(new_n715), .A4(new_n703), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G134), .ZN(G36));
  AOI21_X1  g534(.A(new_n602), .B1(new_n610), .B2(new_n609), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT43), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n590), .B1(new_n370), .B2(new_n634), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(KEYINPUT107), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n579), .B(KEYINPUT45), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(KEYINPUT46), .A3(new_n706), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n574), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT46), .B1(new_n729), .B2(new_n706), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n582), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n733), .A2(new_n656), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n725), .B2(new_n724), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n727), .A2(new_n703), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G137), .ZN(G39));
  XOR2_X1   g551(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n738));
  NOR2_X1   g552(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n739));
  MUX2_X1   g553(.A(new_n738), .B(new_n739), .S(new_n733), .Z(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  OR4_X1    g555(.A1(new_n295), .A2(new_n741), .A3(new_n671), .A4(new_n704), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G140), .ZN(G42));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n671), .A2(new_n696), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n722), .A2(new_n460), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT114), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n722), .A2(new_n748), .A3(new_n460), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n745), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n703), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n679), .A2(new_n666), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n741), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n744), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n671), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n650), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n667), .A2(new_n703), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(KEYINPUT116), .Z(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n460), .A3(new_n759), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n760), .A2(new_n602), .A3(new_n611), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n747), .A2(new_n749), .ZN(new_n762));
  INV_X1    g576(.A(new_n745), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n531), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n652), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(KEYINPUT50), .A3(new_n766), .A4(new_n667), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n750), .A2(new_n531), .A3(new_n766), .A4(new_n667), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n761), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n762), .A2(KEYINPUT117), .A3(new_n759), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT117), .B1(new_n762), .B2(new_n759), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n699), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n771), .A2(KEYINPUT119), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT119), .B1(new_n771), .B2(new_n775), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n755), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n741), .B1(new_n779), .B2(new_n753), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT115), .B1(new_n679), .B2(new_n666), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n752), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n771), .A2(new_n775), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n744), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(KEYINPUT118), .A3(new_n744), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n458), .A2(new_n778), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n750), .A2(new_n680), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n760), .A2(new_n612), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n712), .A2(new_n716), .A3(new_n719), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n704), .A2(new_n708), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n793), .A2(KEYINPUT111), .A3(new_n699), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT111), .B1(new_n793), .B2(new_n699), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n639), .A2(new_n635), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n703), .A2(new_n457), .A3(new_n702), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n797), .A2(new_n626), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n792), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n587), .A2(new_n370), .A3(new_n374), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n533), .A2(new_n535), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n613), .A4(new_n590), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n585), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT109), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n585), .A2(new_n806), .A3(new_n803), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n672), .A2(new_n685), .A3(new_n675), .A4(new_n697), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n602), .A2(new_n457), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n802), .A2(new_n466), .A3(new_n810), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(new_n591), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n636), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT110), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n636), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n800), .A2(new_n808), .A3(new_n809), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT112), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n635), .A2(new_n641), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n715), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n687), .A2(new_n627), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n650), .B(new_n824), .C1(new_n820), .C2(new_n821), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n643), .A2(new_n662), .A3(new_n700), .ZN(new_n827));
  OR3_X1    g641(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT52), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT52), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n805), .A2(new_n807), .B1(new_n814), .B2(new_n816), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n800), .A4(new_n809), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n819), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n819), .A2(new_n830), .A3(KEYINPUT53), .A4(new_n833), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n791), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n828), .A2(KEYINPUT53), .A3(new_n829), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n818), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n834), .B2(new_n835), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n838), .B1(new_n791), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n788), .A2(new_n789), .A3(new_n790), .A4(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n671), .B(new_n710), .C1(new_n773), .C2(new_n774), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n844), .B(KEYINPUT48), .Z(new_n845));
  OAI22_X1  g659(.A1(new_n843), .A2(new_n845), .B1(G952), .B2(G953), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT49), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n432), .B(new_n469), .C1(new_n847), .C2(new_n679), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n766), .A2(new_n532), .A3(new_n582), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n848), .B(new_n849), .C1(new_n847), .C2(new_n679), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n611), .A3(new_n757), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n846), .A2(new_n851), .ZN(G75));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n853));
  INV_X1    g667(.A(new_n841), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(G902), .ZN(new_n855));
  INV_X1    g669(.A(G210), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n506), .A2(new_n514), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(new_n512), .Z(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT55), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n857), .B(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n189), .A2(G952), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(G51));
  XNOR2_X1  g677(.A(new_n841), .B(new_n791), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n706), .A2(KEYINPUT57), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n706), .A2(KEYINPUT57), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n572), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n855), .A2(new_n729), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n862), .B1(new_n868), .B2(new_n869), .ZN(G54));
  AND4_X1   g684(.A1(KEYINPUT58), .A2(new_n854), .A3(G475), .A4(G902), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n424), .A2(new_n426), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT120), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n874), .A2(new_n862), .A3(new_n875), .ZN(G60));
  INV_X1    g690(.A(new_n608), .ZN(new_n877));
  NAND2_X1  g691(.A1(G478), .A2(G902), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT59), .Z(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n842), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n879), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n864), .A2(new_n608), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n862), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(G63));
  NAND2_X1  g698(.A1(new_n359), .A2(new_n362), .ZN(new_n885));
  NAND2_X1  g699(.A1(G217), .A2(G902), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT60), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n841), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n883), .A2(KEYINPUT61), .ZN(new_n890));
  INV_X1    g704(.A(new_n840), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n887), .B1(new_n836), .B2(new_n891), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n633), .B(KEYINPUT121), .Z(new_n893));
  AOI21_X1  g707(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n885), .C1(new_n841), .C2(new_n887), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n889), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n889), .A2(new_n894), .A3(KEYINPUT124), .A4(new_n896), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n888), .A2(new_n883), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n892), .A2(new_n893), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n888), .A2(KEYINPUT122), .A3(new_n883), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n901), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n901), .A2(new_n909), .A3(KEYINPUT125), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(G66));
  OAI21_X1  g728(.A(G953), .B1(new_n463), .B2(new_n510), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n831), .A2(new_n809), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n858), .B1(G898), .B2(new_n189), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G69));
  INV_X1    g733(.A(new_n827), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n659), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT62), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n657), .A2(new_n531), .A3(new_n529), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n612), .B1(new_n457), .B2(new_n602), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n923), .A2(new_n376), .A3(new_n378), .A4(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n742), .A2(new_n736), .A3(new_n925), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n189), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n267), .A2(new_n268), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n415), .B(KEYINPUT126), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(G900), .B2(new_n189), .ZN(new_n933));
  INV_X1    g747(.A(new_n792), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n742), .A2(new_n736), .A3(new_n920), .A4(new_n934), .ZN(new_n935));
  NOR4_X1   g749(.A1(new_n734), .A2(new_n627), .A3(new_n687), .A4(new_n711), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT127), .Z(new_n937));
  OR2_X1    g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n933), .B1(new_n938), .B2(new_n189), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n932), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(G953), .B1(new_n563), .B2(new_n640), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n940), .B(new_n941), .Z(G72));
  NAND2_X1  g756(.A1(G472), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT63), .Z(new_n944));
  INV_X1    g758(.A(new_n270), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(new_n646), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n927), .A2(new_n646), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n938), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n916), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n883), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n945), .A2(new_n646), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n836), .B2(new_n837), .ZN(new_n952));
  AOI211_X1 g766(.A(new_n946), .B(new_n950), .C1(new_n944), .C2(new_n952), .ZN(G57));
endmodule


