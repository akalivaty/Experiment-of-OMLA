//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT64), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT3), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n473), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n472), .A2(new_n476), .A3(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n471), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n470), .A2(new_n475), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n475), .A2(G138), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n473), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n468), .A2(new_n469), .A3(new_n488), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n491), .A2(KEYINPUT65), .A3(KEYINPUT4), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n468), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n496), .A2(new_n500), .ZN(G164));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT66), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n504), .A2(new_n505), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(G50), .A2(new_n516), .B1(new_n520), .B2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n514), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n510), .A2(KEYINPUT67), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n525), .A2(new_n526), .A3(G63), .A4(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT68), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n513), .A2(G89), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT69), .B(G51), .Z(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n516), .A2(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT70), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n528), .A2(new_n537), .A3(new_n529), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(G168));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n525), .A2(new_n526), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n516), .A2(G52), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n512), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n541), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n513), .A2(G81), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n552), .B(new_n553), .C1(new_n554), .C2(new_n515), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT71), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  AND3_X1   g137(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT66), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT66), .B1(new_n509), .B2(new_n510), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT72), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n508), .A2(new_n566), .A3(new_n511), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G91), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OR3_X1    g145(.A1(new_n515), .A2(KEYINPUT9), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT9), .B1(new_n515), .B2(new_n570), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT73), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n518), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n571), .A2(new_n572), .B1(new_n576), .B2(G651), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n569), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n541), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G49), .B2(new_n516), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n565), .A2(G87), .A3(new_n567), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G288));
  AOI22_X1  g160(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G651), .ZN(new_n587));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n586), .A2(new_n587), .B1(new_n588), .B2(new_n515), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n565), .A2(G86), .A3(new_n567), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT74), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n565), .A2(new_n592), .A3(G86), .A4(new_n567), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n589), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n541), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT75), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n513), .A2(G85), .B1(G47), .B2(new_n516), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n599), .A2(new_n600), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT76), .B(G66), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n510), .A2(new_n608), .B1(G79), .B2(G543), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G54), .B2(new_n516), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n568), .A2(G92), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n568), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n607), .B1(new_n617), .B2(G868), .ZN(G284));
  XNOR2_X1  g193(.A(G284), .B(KEYINPUT77), .ZN(G321));
  NOR2_X1   g194(.A1(G299), .A2(G868), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G168), .B2(G868), .ZN(G297));
  XOR2_X1   g196(.A(G297), .B(KEYINPUT78), .Z(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n556), .ZN(G323));
  XOR2_X1   g202(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n628));
  XNOR2_X1  g203(.A(G323), .B(new_n628), .ZN(G282));
  NAND2_X1  g204(.A1(new_n477), .A2(new_n473), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT13), .Z(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n471), .A2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n481), .A2(G123), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n632), .A2(G2100), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT82), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  OAI21_X1  g232(.A(G14), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n657), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT84), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n655), .A2(new_n661), .A3(new_n657), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n658), .B1(new_n660), .B2(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT85), .ZN(new_n666));
  NOR2_X1   g241(.A1(G2072), .A2(G2078), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n444), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n664), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n668), .B(KEYINPUT17), .Z(new_n671));
  OAI21_X1  g246(.A(new_n670), .B1(new_n671), .B2(new_n666), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n665), .A3(new_n664), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n666), .A3(new_n664), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n684), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n681), .A2(KEYINPUT20), .A3(new_n684), .ZN(new_n690));
  OAI221_X1 g265(.A(new_n686), .B1(new_n681), .B2(new_n685), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT87), .ZN(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n692), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT88), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  INV_X1    g275(.A(G34), .ZN(new_n701));
  AOI21_X1  g276(.A(G29), .B1(new_n701), .B2(KEYINPUT24), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(KEYINPUT24), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G160), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G2084), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n638), .A2(new_n705), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n706), .A2(new_n707), .B1(KEYINPUT97), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n471), .A2(G141), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n481), .A2(G129), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT26), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  AOI22_X1  g290(.A1(G105), .A2(new_n477), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n710), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G32), .B(new_n717), .S(G29), .Z(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n708), .A2(KEYINPUT97), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT31), .B(G11), .Z(new_n723));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n705), .B1(new_n724), .B2(G28), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT98), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n726), .A2(KEYINPUT98), .B1(new_n724), .B2(G28), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n709), .A2(new_n721), .A3(new_n722), .A4(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G5), .A2(G16), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G171), .B2(G16), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1961), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n705), .A2(G27), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G164), .B2(new_n705), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2078), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n730), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n706), .A2(new_n707), .B1(new_n718), .B2(new_n720), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT96), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n705), .A2(G33), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  AOI22_X1  g318(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  INV_X1    g319(.A(new_n471), .ZN(new_n745));
  INV_X1    g320(.A(G139), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n743), .B1(new_n475), .B2(new_n744), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2072), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n739), .A2(new_n740), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n748), .B(new_n442), .ZN(new_n751));
  OAI21_X1  g326(.A(KEYINPUT96), .B1(new_n751), .B2(new_n738), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n536), .B2(new_n538), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G21), .ZN(new_n756));
  OR3_X1    g331(.A1(new_n755), .A2(G1966), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(G1966), .B1(new_n755), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n737), .A2(new_n753), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT99), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n737), .A2(new_n753), .A3(new_n759), .A4(KEYINPUT99), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT89), .B(G16), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G20), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT23), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1956), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n705), .A2(G35), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n705), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT29), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G2090), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n774), .A2(KEYINPUT100), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n705), .A2(G26), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT28), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n471), .A2(G140), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n481), .A2(G128), .ZN(new_n779));
  INV_X1    g354(.A(G104), .ZN(new_n780));
  AND3_X1   g355(.A1(new_n780), .A2(new_n475), .A3(KEYINPUT95), .ZN(new_n781));
  AOI21_X1  g356(.A(KEYINPUT95), .B1(new_n780), .B2(new_n475), .ZN(new_n782));
  OAI221_X1 g357(.A(G2104), .B1(G116), .B2(new_n475), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n778), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(G29), .ZN(new_n785));
  INV_X1    g360(.A(G2067), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n765), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(G19), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n556), .B2(new_n788), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT94), .B(G1341), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n792), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n787), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(G4), .A2(G16), .ZN(new_n796));
  INV_X1    g371(.A(new_n617), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n754), .ZN(new_n798));
  INV_X1    g373(.A(G1348), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n772), .A2(G2090), .ZN(new_n801));
  OAI211_X1 g376(.A(G1348), .B(new_n796), .C1(new_n797), .C2(new_n754), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n795), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n774), .A2(KEYINPUT100), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n775), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n764), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT101), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT101), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n764), .A2(new_n808), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n811));
  NAND2_X1  g386(.A1(G288), .A2(KEYINPUT90), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n584), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G16), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G16), .B2(G23), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT33), .B(G1976), .Z(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n594), .A2(new_n754), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G6), .B2(new_n754), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT32), .B(G1981), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n823), .A2(new_n825), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n788), .A2(G22), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G166), .B2(new_n788), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT91), .B(G1971), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n817), .B(new_n819), .C1(G16), .C2(G23), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n827), .A2(new_n828), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n834), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n821), .A2(new_n835), .A3(new_n826), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT92), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n836), .A2(new_n839), .A3(KEYINPUT34), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n765), .A2(G24), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n605), .B2(new_n765), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n842), .A2(G1986), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(G1986), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n471), .A2(G131), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n481), .A2(G119), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n475), .A2(G107), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n845), .B(new_n846), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  MUX2_X1   g424(.A(G25), .B(new_n849), .S(G29), .Z(new_n850));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G1991), .Z(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  NOR4_X1   g428(.A1(new_n843), .A2(new_n844), .A3(new_n853), .A4(KEYINPUT93), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n840), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT34), .B1(new_n836), .B2(new_n839), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n811), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n856), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n858), .A2(KEYINPUT36), .A3(new_n840), .A4(new_n854), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n810), .A2(new_n857), .A3(new_n859), .ZN(G311));
  NAND3_X1  g435(.A1(new_n810), .A2(new_n857), .A3(new_n859), .ZN(G150));
  NAND2_X1  g436(.A1(G80), .A2(G543), .ZN(new_n862));
  INV_X1    g437(.A(G67), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n541), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n864), .A2(KEYINPUT102), .A3(G651), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(G651), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n513), .A2(G93), .B1(G55), .B2(new_n516), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n555), .A2(new_n865), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(new_n869), .ZN(new_n874));
  INV_X1    g449(.A(new_n865), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n873), .B1(new_n876), .B2(new_n555), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n556), .B(KEYINPUT103), .C1(new_n874), .C2(new_n875), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(KEYINPUT38), .B1(new_n797), .B2(new_n623), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n617), .A2(new_n882), .A3(G559), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n872), .A2(new_n879), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G860), .B1(new_n888), .B2(KEYINPUT39), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n884), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n891), .A2(KEYINPUT105), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(KEYINPUT105), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(G860), .B1(new_n874), .B2(new_n875), .ZN(new_n895));
  XOR2_X1   g470(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(KEYINPUT107), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(G145));
  AND3_X1   g477(.A1(new_n491), .A2(KEYINPUT65), .A3(KEYINPUT4), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT65), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n489), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n497), .A2(new_n906), .A3(new_n499), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n497), .B2(new_n499), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(new_n784), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(new_n717), .Z(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n747), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n911), .B(new_n717), .ZN(new_n914));
  INV_X1    g489(.A(new_n747), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n471), .A2(G142), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n481), .A2(G130), .ZN(new_n919));
  OR2_X1    g494(.A1(G106), .A2(G2105), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n920), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n849), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n849), .A2(new_n923), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n631), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n631), .B1(new_n924), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n925), .ZN(new_n930));
  INV_X1    g505(.A(new_n631), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n922), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n926), .A3(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n929), .A2(KEYINPUT110), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT110), .B1(new_n929), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n917), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(G160), .B(new_n638), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(G162), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n927), .A2(new_n922), .A3(new_n928), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n933), .B1(new_n932), .B2(new_n926), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n938), .B(new_n941), .C1(new_n944), .C2(new_n917), .ZN(new_n945));
  INV_X1    g520(.A(G37), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n913), .B(new_n916), .C1(new_n935), .C2(new_n936), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n938), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n945), .B(new_n946), .C1(new_n948), .C2(new_n941), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g525(.A1(G290), .A2(new_n594), .ZN(new_n951));
  NAND2_X1  g526(.A1(G305), .A2(new_n605), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n816), .A2(G303), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n815), .A2(G166), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n951), .A2(new_n954), .A3(new_n955), .A4(new_n952), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT113), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n957), .A2(KEYINPUT112), .A3(new_n959), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT112), .B1(new_n957), .B2(new_n959), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT42), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n625), .A2(KEYINPUT111), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n617), .B2(new_n623), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n880), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n886), .B1(new_n966), .B2(new_n968), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n797), .A2(G299), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n617), .A2(new_n569), .A3(new_n577), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT41), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(KEYINPUT41), .A3(new_n974), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n975), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(new_n972), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n965), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n965), .A2(new_n982), .ZN(new_n984));
  OAI21_X1  g559(.A(G868), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(G868), .B2(new_n876), .ZN(G295));
  OAI21_X1  g561(.A(new_n985), .B1(G868), .B2(new_n876), .ZN(G331));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g564(.A1(G286), .A2(G301), .ZN(new_n990));
  AOI21_X1  g565(.A(G301), .B1(new_n536), .B2(new_n538), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n886), .A2(new_n993), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n879), .A2(new_n872), .B1(new_n990), .B2(new_n992), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n981), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n886), .A2(new_n993), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n872), .A2(new_n990), .A3(new_n879), .A4(new_n992), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(new_n977), .A3(new_n998), .A4(new_n978), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n962), .A2(new_n963), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n996), .B(new_n999), .C1(new_n962), .C2(new_n963), .ZN(new_n1003));
  AND4_X1   g578(.A1(new_n989), .A2(new_n1002), .A3(new_n946), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G37), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n989), .B1(new_n1005), .B2(new_n1003), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n988), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1002), .A2(new_n946), .A3(new_n1003), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT43), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1005), .A2(new_n989), .A3(new_n1003), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(KEYINPUT44), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1011), .ZN(G397));
  AOI21_X1  g587(.A(G1384), .B1(new_n905), .B2(new_n909), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n472), .A2(new_n476), .A3(G40), .A4(new_n478), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1013), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n784), .B(new_n786), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n717), .B(G1996), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n849), .B(new_n852), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT115), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1015), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1986), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n605), .B(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1026), .B1(new_n1015), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1014), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1013), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G288), .A2(G1976), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT118), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n508), .A2(G86), .A3(new_n511), .ZN(new_n1035));
  OAI21_X1  g610(.A(G1981), .B1(new_n1035), .B2(new_n589), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT116), .B(G1981), .C1(new_n1035), .C2(new_n589), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1981), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n594), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT49), .B1(new_n1042), .B2(KEYINPUT117), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT49), .ZN(new_n1045));
  AOI211_X1 g620(.A(G1981), .B(new_n589), .C1(new_n591), .C2(new_n593), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1044), .B(new_n1045), .C1(new_n1046), .C2(new_n1040), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1034), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1032), .B1(new_n1048), .B2(new_n1046), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G1384), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n500), .A2(KEYINPUT108), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n497), .A2(new_n906), .A3(new_n499), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n496), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n500), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1384), .B1(new_n905), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1055), .B(new_n1031), .C1(new_n1057), .C2(KEYINPUT45), .ZN(new_n1058));
  INV_X1    g633(.A(G1971), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n1061));
  INV_X1    g636(.A(G1384), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1061), .B(new_n1062), .C1(new_n496), .C2(new_n1054), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(new_n1031), .C1(new_n1061), .C2(new_n1057), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1060), .B1(G2090), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G303), .A2(G8), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT55), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(G8), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1043), .A2(new_n1032), .A3(new_n1047), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n812), .A2(G1976), .A3(new_n814), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(new_n1032), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1072), .A2(new_n1032), .ZN(new_n1074));
  INV_X1    g649(.A(G1976), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(G288), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1073), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1070), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1049), .B1(new_n1069), .B2(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1070), .A2(new_n1077), .ZN(new_n1080));
  NOR2_X1   g655(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n496), .B2(new_n500), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(new_n1031), .C1(new_n1013), .C2(new_n1061), .ZN(new_n1083));
  AOI21_X1  g658(.A(G2090), .B1(new_n1083), .B2(KEYINPUT119), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1062), .B1(new_n496), .B2(new_n1054), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT50), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n905), .A2(new_n1056), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1014), .B1(new_n1087), .B2(new_n1081), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1084), .A2(new_n1090), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1067), .B1(new_n1091), .B2(new_n1030), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G168), .A2(G8), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1087), .A2(new_n1051), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(new_n1031), .C1(KEYINPUT45), .C2(new_n1013), .ZN(new_n1095));
  INV_X1    g670(.A(G1966), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1014), .B1(new_n1013), .B2(new_n1061), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(KEYINPUT120), .A4(new_n707), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1064), .B2(G2084), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1093), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1080), .A2(new_n1092), .A3(new_n1069), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT63), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1065), .A2(G8), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1108), .B2(new_n1067), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1080), .A2(new_n1109), .A3(new_n1069), .A4(new_n1104), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1079), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1080), .A2(new_n1092), .A3(new_n1069), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1058), .B2(G2078), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1014), .B1(new_n1085), .B2(new_n1050), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1115), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1094), .ZN(new_n1116));
  INV_X1    g691(.A(G1961), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1064), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT54), .B1(new_n1119), .B2(G171), .ZN(new_n1120));
  AOI211_X1 g695(.A(new_n1113), .B(G2078), .C1(new_n910), .C2(new_n1051), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1117), .A2(new_n1064), .B1(new_n1121), .B2(new_n1115), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(KEYINPUT124), .A3(new_n1114), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1115), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1114), .A2(new_n1118), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n1126));
  AOI21_X1  g701(.A(G301), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1120), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1112), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1103), .A2(G168), .A3(new_n1097), .A4(new_n1100), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(G8), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1131), .A2(KEYINPUT51), .ZN(new_n1132));
  AOI21_X1  g707(.A(G168), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT51), .B1(new_n1133), .B2(new_n1131), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n1136));
  XNOR2_X1  g711(.A(G299), .B(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1050), .B1(G164), .B2(G1384), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT56), .B(G2072), .Z(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1138), .A2(new_n1031), .A3(new_n1055), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1956), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1083), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1137), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n910), .A2(new_n1031), .A3(new_n1062), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT121), .B1(new_n1145), .B2(G2067), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1013), .A2(new_n1147), .A3(new_n786), .A4(new_n1031), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(G1348), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n797), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(G299), .B(KEYINPUT57), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1058), .A2(new_n1139), .ZN(new_n1155));
  AOI21_X1  g730(.A(G1956), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1144), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT58), .B(G1341), .Z(new_n1160));
  NAND2_X1  g735(.A1(new_n1145), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1014), .A2(G1996), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1055), .B(new_n1162), .C1(new_n1057), .C2(KEYINPUT45), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n555), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1157), .A2(new_n1144), .A3(KEYINPUT61), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n617), .A2(KEYINPUT60), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n617), .A2(KEYINPUT60), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1150), .A2(new_n1152), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(KEYINPUT60), .B(new_n617), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1166), .A2(new_n1167), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT61), .B1(new_n1157), .B2(new_n1144), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1159), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1129), .A2(new_n1135), .A3(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1114), .A2(new_n1118), .A3(G301), .A4(new_n1124), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1119), .A2(G171), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1122), .A2(KEYINPUT122), .A3(G301), .A4(new_n1114), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(KEYINPUT123), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1181), .A2(new_n1185), .A3(new_n1182), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1111), .B1(new_n1175), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1112), .A2(new_n1179), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1189), .B1(new_n1135), .B2(KEYINPUT62), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1029), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n784), .A2(G2067), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n849), .A2(new_n852), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1195), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g776(.A(KEYINPUT125), .B(new_n1195), .C1(new_n1196), .C2(new_n1198), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1201), .A2(new_n1015), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(G1996), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1015), .A2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT46), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1015), .B1(new_n1017), .B2(new_n717), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT47), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1015), .A2(new_n1027), .A3(new_n605), .ZN(new_n1210));
  XOR2_X1   g785(.A(new_n1210), .B(KEYINPUT48), .Z(new_n1211));
  OR2_X1    g786(.A1(new_n1026), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1203), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1213), .A2(KEYINPUT126), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1203), .A2(new_n1209), .A3(new_n1215), .A4(new_n1212), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1194), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g793(.A1(G227), .A2(new_n462), .ZN(new_n1220));
  INV_X1    g794(.A(new_n1220), .ZN(new_n1221));
  OAI21_X1  g795(.A(KEYINPUT127), .B1(G401), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n1222), .A2(new_n699), .ZN(new_n1223));
  NOR3_X1   g797(.A1(G401), .A2(KEYINPUT127), .A3(new_n1221), .ZN(new_n1224));
  NOR2_X1   g798(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g799(.A(new_n949), .B(new_n1225), .C1(new_n1004), .C2(new_n1006), .ZN(G225));
  INV_X1    g800(.A(G225), .ZN(G308));
endmodule


