//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160,
    new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT64), .Z(G173));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(KEYINPUT67), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(KEYINPUT67), .B2(new_n461), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT69), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n467), .A2(G137), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n466), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT68), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n466), .A2(new_n475), .A3(new_n479), .A4(G125), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n478), .A2(new_n480), .B1(G113), .B2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n473), .B1(new_n481), .B2(new_n468), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(G160));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n467), .A2(new_n469), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n468), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(G2105), .ZN(new_n490));
  OAI221_X1 g065(.A(new_n485), .B1(new_n487), .B2(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  AND2_X1   g067(.A1(new_n468), .A2(G138), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n474), .B2(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n474), .A2(G2104), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n469), .B(new_n493), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n467), .A2(KEYINPUT73), .A3(new_n469), .A4(new_n493), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(KEYINPUT4), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n476), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n502), .A2(KEYINPUT74), .A3(new_n503), .A4(new_n493), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n493), .A2(new_n503), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(new_n476), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n467), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n468), .A2(G114), .ZN(new_n511));
  OAI21_X1  g086(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT71), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(G102), .A2(G2105), .ZN(new_n514));
  INV_X1    g089(.A(G114), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G2105), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n514), .A2(new_n516), .A3(new_n517), .A4(G2104), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n510), .A2(new_n519), .A3(KEYINPUT72), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n509), .A2(new_n524), .ZN(G164));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT5), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n530), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT75), .B(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G50), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n530), .ZN(new_n535));
  INV_X1    g110(.A(G88), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT75), .ZN(new_n539));
  NAND2_X1  g114(.A1(KEYINPUT76), .A2(G651), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n539), .B(KEYINPUT6), .C1(KEYINPUT75), .C2(new_n540), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n540), .A2(KEYINPUT6), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n533), .B1(new_n537), .B2(new_n543), .ZN(G166));
  NAND2_X1  g119(.A1(new_n543), .A2(KEYINPUT77), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n541), .A2(new_n542), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n545), .A2(G543), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G51), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n543), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n535), .ZN(new_n552));
  NAND3_X1  g127(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT7), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(G286));
  INV_X1    g130(.A(G286), .ZN(G168));
  AOI22_X1  g131(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n532), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT78), .Z(new_n559));
  NAND2_X1  g134(.A1(new_n549), .A2(G52), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n546), .A2(new_n535), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G90), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(G301));
  INV_X1    g138(.A(G301), .ZN(G171));
  AOI22_X1  g139(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(new_n532), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(G81), .B2(new_n561), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n545), .A2(G43), .A3(G543), .A4(new_n548), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  NAND3_X1  g150(.A1(new_n549), .A2(KEYINPUT9), .A3(G53), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(G65), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(G65), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n530), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G78), .A2(G543), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT79), .Z(new_n582));
  AOI21_X1  g157(.A(new_n538), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(G91), .B2(new_n561), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT9), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n545), .A2(G543), .A3(new_n548), .ZN(new_n586));
  INV_X1    g161(.A(G53), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n576), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G299));
  INV_X1    g167(.A(G166), .ZN(G303));
  NAND2_X1  g168(.A1(new_n549), .A2(G49), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n561), .A2(G87), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  AOI22_X1  g172(.A1(new_n530), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n546), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n530), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n532), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(G305));
  XOR2_X1   g177(.A(KEYINPUT82), .B(G47), .Z(new_n603));
  NAND2_X1  g178(.A1(new_n549), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n532), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT83), .B(G85), .Z(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n561), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n561), .A2(G92), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G54), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n530), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n586), .A2(new_n613), .B1(new_n538), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT84), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n610), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n610), .B1(new_n618), .B2(G868), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  XOR2_X1   g196(.A(G299), .B(KEYINPUT85), .Z(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G297));
  XNOR2_X1  g198(.A(G297), .B(KEYINPUT86), .ZN(G280));
  NOR2_X1   g199(.A1(new_n617), .A2(G559), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(G860), .B2(new_n618), .ZN(G148));
  NAND2_X1  g201(.A1(new_n567), .A2(new_n568), .ZN(new_n627));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n625), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g206(.A(new_n490), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G123), .ZN(new_n633));
  INV_X1    g208(.A(new_n487), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G135), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n468), .A2(G111), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n633), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND3_X1  g214(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  NOR2_X1   g217(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n643));
  AND2_X1   g218(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n639), .B(new_n645), .C1(new_n643), .C2(new_n642), .ZN(G156));
  XOR2_X1   g221(.A(KEYINPUT88), .B(G2438), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT89), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT14), .ZN(new_n653));
  XOR2_X1   g228(.A(G2443), .B(G2446), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1341), .B(G1348), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(new_n659), .Z(new_n660));
  AND2_X1   g235(.A1(new_n660), .A2(G14), .ZN(G401));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(KEYINPUT90), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n668), .B2(new_n662), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n664), .B(KEYINPUT17), .Z(new_n670));
  OAI21_X1  g245(.A(new_n669), .B1(new_n662), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n662), .A3(new_n665), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(new_n677), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n686), .B(new_n687), .C1(new_n685), .C2(new_n684), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  INV_X1    g266(.A(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n690), .B(new_n694), .ZN(G229));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G35), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G162), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G2090), .ZN(new_n700));
  NAND2_X1  g275(.A1(G168), .A2(G16), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G16), .B2(G21), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT101), .B(G1966), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT102), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G5), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G171), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1961), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT28), .ZN(new_n711));
  INV_X1    g286(.A(G26), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G29), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n632), .A2(G128), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n634), .A2(G140), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n468), .A2(G116), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n714), .B1(new_n719), .B2(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n713), .B1(new_n720), .B2(new_n711), .ZN(new_n721));
  INV_X1    g296(.A(G11), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n721), .A2(G2067), .B1(KEYINPUT31), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n696), .A2(G27), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G164), .B2(new_n696), .ZN(new_n725));
  OR2_X1    g300(.A1(KEYINPUT24), .A2(G34), .ZN(new_n726));
  NAND2_X1  g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n726), .A2(new_n696), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G160), .B2(new_n696), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n723), .B1(G2078), .B2(new_n725), .C1(G2084), .C2(new_n729), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n706), .A2(new_n710), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n702), .A2(new_n704), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT30), .B(G28), .Z(new_n733));
  MUX2_X1   g308(.A(new_n733), .B(new_n638), .S(G29), .Z(new_n734));
  NOR2_X1   g309(.A1(G29), .A2(G32), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n634), .A2(G141), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n632), .A2(G129), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT99), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT26), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT100), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n735), .B1(new_n743), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n732), .B(new_n734), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n722), .A2(KEYINPUT31), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT98), .B1(G29), .B2(G33), .ZN(new_n751));
  OR3_X1    g326(.A1(KEYINPUT98), .A2(G29), .A3(G33), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  AOI22_X1  g329(.A1(new_n502), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  INV_X1    g330(.A(G139), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n754), .B1(new_n755), .B2(new_n468), .C1(new_n487), .C2(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n751), .B(new_n752), .C1(new_n757), .C2(new_n696), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2072), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n731), .A2(new_n749), .A3(new_n750), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G4), .A2(G16), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n618), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT97), .B(G1348), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n707), .A2(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n569), .B2(new_n707), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1341), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n699), .A2(G2090), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n767), .B(new_n768), .C1(G2084), .C2(new_n729), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n764), .B(new_n769), .C1(G2067), .C2(new_n721), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(G25), .A2(G29), .ZN(new_n772));
  INV_X1    g347(.A(G131), .ZN(new_n773));
  OR3_X1    g348(.A1(new_n487), .A2(KEYINPUT91), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n632), .A2(G119), .ZN(new_n775));
  OR2_X1    g350(.A1(G95), .A2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n777));
  OAI21_X1  g352(.A(KEYINPUT91), .B1(new_n487), .B2(new_n773), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n774), .A2(new_n775), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT92), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n772), .B1(new_n780), .B2(new_n696), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n781), .A2(KEYINPUT93), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(KEYINPUT93), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT35), .B(G1991), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n784), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G24), .ZN(new_n788));
  INV_X1    g363(.A(G290), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G16), .ZN(new_n790));
  INV_X1    g365(.A(G1986), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT36), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n707), .A2(G23), .ZN(new_n795));
  INV_X1    g370(.A(G288), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(new_n707), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT33), .B(G1976), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT96), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n797), .B(new_n799), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n707), .A2(G6), .ZN(new_n801));
  INV_X1    g376(.A(G305), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n707), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT95), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT32), .B(G1981), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n707), .A2(G22), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n707), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1971), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n800), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT94), .B(KEYINPUT34), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n793), .A2(new_n794), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n794), .B1(new_n793), .B2(new_n812), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n700), .B(new_n771), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n707), .A2(G20), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT103), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT23), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G299), .B2(G16), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT104), .B(G1956), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n725), .A2(G2078), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n815), .A2(new_n821), .A3(new_n823), .ZN(G311));
  INV_X1    g399(.A(new_n771), .ZN(new_n825));
  INV_X1    g400(.A(new_n814), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n793), .A2(new_n794), .A3(new_n812), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n821), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n828), .A2(new_n829), .A3(new_n822), .A4(new_n700), .ZN(G150));
  XNOR2_X1  g405(.A(KEYINPUT105), .B(G55), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n549), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n532), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  INV_X1    g409(.A(G67), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n535), .B2(new_n835), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n833), .A2(new_n836), .B1(new_n561), .B2(G93), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT37), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n618), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT39), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n841), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n838), .A2(new_n569), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n627), .A2(new_n832), .A3(new_n837), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n844), .B(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n840), .B1(new_n849), .B2(G860), .ZN(G145));
  XNOR2_X1  g425(.A(G160), .B(new_n638), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G162), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n780), .B(new_n743), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n501), .A2(new_n508), .ZN(new_n855));
  INV_X1    g430(.A(new_n520), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n641), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n757), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n634), .A2(G142), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n468), .A2(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G130), .B2(new_n632), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n719), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n859), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n854), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n854), .A2(new_n867), .ZN(new_n869));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g447(.A(new_n625), .B(new_n848), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n590), .A2(new_n591), .A3(new_n616), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n616), .B1(new_n590), .B2(new_n591), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n874), .B2(new_n875), .ZN(new_n879));
  INV_X1    g454(.A(new_n616), .ZN(new_n880));
  NAND2_X1  g455(.A1(G299), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n590), .A2(new_n591), .A3(new_n616), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n877), .B1(new_n873), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  XNOR2_X1  g463(.A(G288), .B(G290), .ZN(new_n889));
  XOR2_X1   g464(.A(G166), .B(G305), .Z(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n887), .B2(new_n888), .ZN(new_n894));
  OAI21_X1  g469(.A(G868), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n838), .A2(new_n628), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(G295));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n896), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n845), .A2(new_n846), .A3(G286), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G286), .B1(new_n845), .B2(new_n846), .ZN(new_n902));
  OAI21_X1  g477(.A(G301), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(G171), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n881), .A2(new_n882), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n876), .A2(KEYINPUT107), .A3(new_n905), .A4(new_n903), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n879), .A3(new_n883), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n891), .A4(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n908), .A2(new_n912), .A3(new_n891), .A4(new_n909), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT108), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n908), .A2(new_n912), .A3(new_n909), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n892), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n913), .A2(new_n870), .A3(new_n915), .A4(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n876), .A2(new_n905), .A3(new_n903), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n912), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n923), .B(new_n892), .C1(new_n921), .C2(new_n922), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n913), .A2(new_n924), .A3(new_n870), .A4(new_n915), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n925), .A2(new_n919), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT44), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n914), .B(new_n911), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n928), .A2(new_n919), .A3(new_n870), .A4(new_n924), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n927), .B1(KEYINPUT44), .B2(new_n931), .ZN(G397));
  NOR2_X1   g507(.A1(G290), .A2(G1986), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT112), .ZN(new_n934));
  AOI21_X1  g509(.A(G1384), .B1(new_n855), .B2(new_n856), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT110), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n520), .B1(new_n501), .B2(new_n508), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n939), .B2(G1384), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT111), .B(G40), .Z(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n473), .B(new_n943), .C1(new_n481), .C2(new_n468), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n934), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT127), .ZN(new_n948));
  XOR2_X1   g523(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n949));
  XNOR2_X1  g524(.A(new_n948), .B(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n719), .A2(G2067), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n719), .A2(G2067), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(KEYINPUT113), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(KEYINPUT113), .ZN(new_n955));
  INV_X1    g530(.A(G1996), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n743), .B(new_n956), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n954), .A2(new_n955), .B1(new_n945), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n780), .B(new_n786), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n946), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n780), .A2(new_n785), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n952), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n950), .A2(new_n960), .B1(new_n962), .B2(new_n946), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n953), .B1(new_n743), .B2(new_n946), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT125), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n946), .A2(G1996), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT46), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT118), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  NOR2_X1   g547(.A1(G166), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT55), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT116), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(KEYINPUT116), .A3(KEYINPUT55), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n976), .B(new_n977), .C1(KEYINPUT55), .C2(new_n973), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n857), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n478), .A2(new_n480), .ZN(new_n981));
  NAND2_X1  g556(.A1(G113), .A2(G2104), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n468), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n983), .A2(new_n472), .A3(new_n942), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n510), .A2(KEYINPUT72), .A3(new_n519), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT72), .B1(new_n510), .B2(new_n519), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n988), .B2(new_n855), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT114), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n979), .B1(new_n509), .B2(new_n524), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n937), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n944), .B1(new_n935), .B2(KEYINPUT45), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G1971), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n999));
  AOI21_X1  g574(.A(new_n944), .B1(new_n935), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(G2090), .ZN(new_n1002));
  OAI211_X1 g577(.A(G8), .B(new_n978), .C1(new_n997), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1976), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(G288), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n972), .B1(new_n935), .B2(new_n984), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1005), .B(new_n1006), .C1(new_n1004), .C2(G288), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1004), .B2(G288), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT52), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n802), .A2(new_n692), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G305), .A2(G1981), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(KEYINPUT49), .A3(new_n1011), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n1006), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1007), .A2(new_n1009), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1971), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n995), .B1(new_n993), .B2(new_n994), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n935), .A2(new_n984), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n984), .A2(new_n999), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(KEYINPUT117), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G2090), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n989), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(new_n984), .C1(new_n935), .C2(new_n999), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n972), .B1(new_n1022), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1003), .B(new_n1018), .C1(new_n1032), .C2(new_n978), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n984), .B1(new_n935), .B2(KEYINPUT45), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n937), .B(G1384), .C1(new_n988), .C2(new_n855), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n704), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G2084), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n998), .A2(new_n1000), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n972), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G168), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n971), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT63), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1002), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n972), .B1(new_n1022), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1017), .B1(new_n1044), .B2(new_n978), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1031), .ZN(new_n1046));
  OAI21_X1  g621(.A(G8), .B1(new_n997), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n978), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1040), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1045), .A2(KEYINPUT118), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1041), .A2(new_n1042), .A3(new_n1051), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1044), .A2(new_n978), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1053), .A2(new_n1045), .A3(KEYINPUT63), .A4(new_n1050), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1016), .A2(new_n1004), .A3(new_n796), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1010), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1006), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1003), .B2(new_n1017), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1036), .A2(new_n1038), .A3(G168), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G8), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT51), .B1(new_n1039), .B2(KEYINPUT121), .ZN(new_n1063));
  AOI21_X1  g638(.A(G168), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1061), .B(KEYINPUT51), .C1(KEYINPUT121), .C2(new_n1039), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G2078), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n991), .A2(new_n1069), .A3(new_n996), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1071), .A2(G2078), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G1961), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1001), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1072), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(G301), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1033), .B1(new_n1081), .B2(KEYINPUT62), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1059), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1348), .B1(new_n998), .B2(new_n1000), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1023), .A2(G2067), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n857), .A2(new_n979), .A3(new_n999), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n984), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n989), .A2(new_n1027), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1086), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT120), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1087), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1025), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1096));
  INV_X1    g671(.A(G1956), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1099), .A2(KEYINPUT57), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n576), .A2(new_n584), .A3(new_n588), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(KEYINPUT57), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1101), .B(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n985), .A2(new_n990), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1098), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1095), .A2(new_n616), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1098), .A2(new_n1106), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1103), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT60), .B1(new_n1087), .B2(new_n1094), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n616), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT60), .B(new_n880), .C1(new_n1087), .C2(new_n1094), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1114), .A2(new_n1115), .B1(new_n1116), .B2(new_n1095), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1098), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1103), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1111), .A2(KEYINPUT61), .A3(new_n1107), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1117), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1104), .A2(new_n956), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1023), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n627), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT59), .Z(new_n1129));
  AOI21_X1  g704(.A(new_n1112), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n481), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(G2105), .B1(new_n481), .B2(new_n1132), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n473), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(KEYINPUT45), .B2(new_n935), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n941), .A2(new_n1136), .A3(G40), .A4(new_n1074), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1137), .A2(new_n1077), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1072), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(G171), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1131), .B1(new_n1079), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1033), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1131), .B1(new_n1078), .B2(G301), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1072), .A2(new_n1138), .A3(KEYINPUT123), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(G171), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1141), .A2(new_n1142), .A3(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1055), .B(new_n1083), .C1(new_n1130), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n934), .B1(new_n791), .B2(new_n789), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n960), .B1(new_n945), .B2(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1151), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n970), .B1(new_n1154), .B2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g731(.A1(new_n929), .A2(new_n930), .ZN(new_n1158));
  AOI21_X1  g732(.A(G227), .B1(new_n660), .B2(G14), .ZN(new_n1159));
  AND2_X1   g733(.A1(new_n1159), .A2(new_n871), .ZN(new_n1160));
  INV_X1    g734(.A(G229), .ZN(new_n1161));
  NAND4_X1  g735(.A1(new_n1158), .A2(new_n1160), .A3(G319), .A4(new_n1161), .ZN(G225));
  INV_X1    g736(.A(G225), .ZN(G308));
endmodule


