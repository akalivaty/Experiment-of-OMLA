

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752;

  NOR2_X1 U381 ( .A1(n586), .A2(n585), .ZN(n587) );
  OR2_X1 U382 ( .A1(n673), .A2(G902), .ZN(n407) );
  INV_X1 U383 ( .A(G953), .ZN(n737) );
  XNOR2_X1 U384 ( .A(n506), .B(n505), .ZN(n700) );
  NOR2_X1 U385 ( .A1(n550), .A2(n524), .ZN(n687) );
  NAND2_X2 U386 ( .A1(n392), .A2(n366), .ZN(n391) );
  XNOR2_X2 U387 ( .A(n391), .B(n390), .ZN(n746) );
  NOR2_X1 U388 ( .A1(n611), .A2(n608), .ZN(n559) );
  NOR2_X2 U389 ( .A1(n623), .A2(n405), .ZN(n404) );
  XNOR2_X2 U390 ( .A(KEYINPUT3), .B(G119), .ZN(n447) );
  NOR2_X2 U391 ( .A1(n555), .A2(n750), .ZN(n413) );
  INV_X1 U392 ( .A(n687), .ZN(n399) );
  NAND2_X1 U393 ( .A1(n578), .A2(n611), .ZN(n585) );
  INV_X1 U394 ( .A(n633), .ZN(n625) );
  NAND2_X1 U395 ( .A1(n521), .A2(n579), .ZN(n522) );
  XNOR2_X1 U396 ( .A(n414), .B(n373), .ZN(n553) );
  NOR2_X1 U397 ( .A1(n615), .A2(n631), .ZN(n619) );
  XNOR2_X1 U398 ( .A(n520), .B(n378), .ZN(n521) );
  NAND2_X1 U399 ( .A1(n580), .A2(n559), .ZN(n520) );
  XNOR2_X1 U400 ( .A(n603), .B(n406), .ZN(n579) );
  OR2_X1 U401 ( .A1(n716), .A2(G902), .ZN(n410) );
  XNOR2_X1 U402 ( .A(n444), .B(n443), .ZN(n551) );
  XOR2_X1 U403 ( .A(n704), .B(KEYINPUT59), .Z(n707) );
  XNOR2_X1 U404 ( .A(n387), .B(n385), .ZN(n704) );
  XNOR2_X1 U405 ( .A(n466), .B(G125), .ZN(n456) );
  XNOR2_X1 U406 ( .A(n721), .B(KEYINPUT69), .ZN(n500) );
  XNOR2_X1 U407 ( .A(n380), .B(KEYINPUT67), .ZN(n468) );
  XNOR2_X1 U408 ( .A(KEYINPUT85), .B(KEYINPUT36), .ZN(n626) );
  INV_X1 U409 ( .A(KEYINPUT39), .ZN(n616) );
  XNOR2_X1 U410 ( .A(KEYINPUT66), .B(G131), .ZN(n380) );
  BUF_X1 U411 ( .A(n658), .Z(n360) );
  XNOR2_X1 U412 ( .A(n460), .B(n459), .ZN(n658) );
  XNOR2_X1 U413 ( .A(n465), .B(n464), .ZN(n653) );
  NOR2_X1 U414 ( .A1(n544), .A2(n525), .ZN(n465) );
  XNOR2_X2 U415 ( .A(n625), .B(n463), .ZN(n601) );
  BUF_X1 U416 ( .A(n664), .Z(n361) );
  BUF_X1 U417 ( .A(n580), .Z(n362) );
  XNOR2_X1 U418 ( .A(n606), .B(KEYINPUT1), .ZN(n580) );
  NOR2_X2 U419 ( .A1(n653), .A2(n598), .ZN(n600) );
  XNOR2_X1 U420 ( .A(n592), .B(n593), .ZN(n384) );
  NAND2_X1 U421 ( .A1(n692), .A2(n399), .ZN(n592) );
  NOR2_X1 U422 ( .A1(G953), .A2(G237), .ZN(n470) );
  XNOR2_X1 U423 ( .A(n456), .B(KEYINPUT10), .ZN(n477) );
  XNOR2_X1 U424 ( .A(n736), .B(n663), .ZN(n665) );
  XNOR2_X1 U425 ( .A(n442), .B(G475), .ZN(n443) );
  NOR2_X1 U426 ( .A1(n704), .A2(G902), .ZN(n444) );
  XNOR2_X1 U427 ( .A(n421), .B(n420), .ZN(n485) );
  INV_X1 U428 ( .A(KEYINPUT8), .ZN(n420) );
  NAND2_X1 U429 ( .A1(n737), .A2(G234), .ZN(n421) );
  XNOR2_X1 U430 ( .A(G119), .B(G128), .ZN(n482) );
  XOR2_X1 U431 ( .A(KEYINPUT24), .B(G110), .Z(n483) );
  XNOR2_X1 U432 ( .A(G113), .B(G143), .ZN(n440) );
  INV_X1 U433 ( .A(n477), .ZN(n479) );
  NAND2_X1 U434 ( .A1(n648), .A2(KEYINPUT2), .ZN(n662) );
  NAND2_X1 U435 ( .A1(G234), .A2(G237), .ZN(n431) );
  INV_X1 U436 ( .A(KEYINPUT102), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n437), .B(n436), .ZN(n550) );
  XNOR2_X1 U438 ( .A(n494), .B(n370), .ZN(n409) );
  XNOR2_X1 U439 ( .A(n676), .B(n675), .ZN(n419) );
  NAND2_X1 U440 ( .A1(n705), .A2(G472), .ZN(n676) );
  XOR2_X1 U441 ( .A(KEYINPUT87), .B(n657), .Z(n718) );
  AND2_X1 U442 ( .A1(n384), .A2(n594), .ZN(n595) );
  INV_X1 U443 ( .A(KEYINPUT104), .ZN(n401) );
  XNOR2_X1 U444 ( .A(G137), .B(G116), .ZN(n473) );
  XOR2_X1 U445 ( .A(G137), .B(G140), .Z(n501) );
  XOR2_X1 U446 ( .A(G902), .B(KEYINPUT15), .Z(n661) );
  XNOR2_X1 U447 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U448 ( .A(G134), .B(G122), .ZN(n434) );
  INV_X1 U449 ( .A(G107), .ZN(n408) );
  XOR2_X1 U450 ( .A(KEYINPUT77), .B(KEYINPUT90), .Z(n498) );
  NOR2_X1 U451 ( .A1(n696), .A2(n382), .ZN(n381) );
  XNOR2_X1 U452 ( .A(n403), .B(n402), .ZN(n383) );
  INV_X1 U453 ( .A(n695), .ZN(n382) );
  NOR2_X1 U454 ( .A1(KEYINPUT2), .A2(n727), .ZN(n570) );
  NOR2_X1 U455 ( .A1(n612), .A2(n611), .ZN(n613) );
  AND2_X1 U456 ( .A1(n584), .A2(n377), .ZN(n543) );
  AND2_X1 U457 ( .A1(n542), .A2(n576), .ZN(n377) );
  INV_X1 U458 ( .A(KEYINPUT6), .ZN(n406) );
  XNOR2_X1 U459 ( .A(n488), .B(n487), .ZN(n716) );
  XNOR2_X1 U460 ( .A(n486), .B(n364), .ZN(n487) );
  XNOR2_X1 U461 ( .A(n426), .B(n424), .ZN(n710) );
  XNOR2_X1 U462 ( .A(n425), .B(n446), .ZN(n424) );
  XNOR2_X1 U463 ( .A(n433), .B(n367), .ZN(n426) );
  XNOR2_X1 U464 ( .A(n435), .B(n434), .ZN(n425) );
  XNOR2_X1 U465 ( .A(n479), .B(n386), .ZN(n385) );
  XNOR2_X1 U466 ( .A(n365), .B(n441), .ZN(n387) );
  XNOR2_X1 U467 ( .A(n429), .B(n440), .ZN(n386) );
  XNOR2_X1 U468 ( .A(n660), .B(n659), .ZN(n670) );
  INV_X1 U469 ( .A(KEYINPUT35), .ZN(n390) );
  XNOR2_X1 U470 ( .A(n523), .B(KEYINPUT100), .ZN(n692) );
  INV_X1 U471 ( .A(n718), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U473 ( .A1(n650), .A2(n416), .ZN(n415) );
  AND2_X1 U474 ( .A1(n651), .A2(n363), .ZN(n416) );
  NOR2_X1 U475 ( .A1(n656), .A2(G953), .ZN(n363) );
  AND2_X1 U476 ( .A1(n485), .A2(G221), .ZN(n364) );
  XOR2_X1 U477 ( .A(n468), .B(n445), .Z(n365) );
  XOR2_X1 U478 ( .A(KEYINPUT78), .B(n632), .Z(n366) );
  XNOR2_X1 U479 ( .A(n432), .B(KEYINPUT98), .ZN(n367) );
  XNOR2_X1 U480 ( .A(KEYINPUT101), .B(n545), .ZN(n368) );
  AND2_X1 U481 ( .A1(n597), .A2(n596), .ZN(n369) );
  XOR2_X1 U482 ( .A(n490), .B(n489), .Z(n370) );
  INV_X1 U483 ( .A(G146), .ZN(n466) );
  XOR2_X1 U484 ( .A(n415), .B(KEYINPUT53), .Z(G75) );
  XNOR2_X1 U485 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n372) );
  XOR2_X1 U486 ( .A(n546), .B(KEYINPUT72), .Z(n373) );
  XOR2_X1 U487 ( .A(n569), .B(KEYINPUT45), .Z(n374) );
  XOR2_X1 U488 ( .A(KEYINPUT63), .B(KEYINPUT109), .Z(n375) );
  XNOR2_X1 U489 ( .A(n376), .B(n504), .ZN(n506) );
  XNOR2_X1 U490 ( .A(n503), .B(n502), .ZN(n376) );
  XNOR2_X1 U491 ( .A(n500), .B(n408), .ZN(n503) );
  XNOR2_X1 U492 ( .A(n549), .B(n372), .ZN(n392) );
  XNOR2_X2 U493 ( .A(n733), .B(G146), .ZN(n505) );
  XNOR2_X2 U494 ( .A(n389), .B(n469), .ZN(n733) );
  NOR2_X1 U495 ( .A1(n708), .A2(n718), .ZN(n709) );
  NOR2_X1 U496 ( .A1(n671), .A2(n718), .ZN(n379) );
  XNOR2_X2 U497 ( .A(n600), .B(n599), .ZN(n752) );
  NAND2_X2 U498 ( .A1(n383), .A2(n381), .ZN(n736) );
  NOR2_X4 U499 ( .A1(n668), .A2(n667), .ZN(n705) );
  NOR2_X1 U500 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U501 ( .A1(n746), .A2(n683), .ZN(n555) );
  XNOR2_X1 U502 ( .A(n379), .B(n672), .ZN(G51) );
  XNOR2_X2 U503 ( .A(n388), .B(G143), .ZN(n467) );
  XNOR2_X2 U504 ( .A(G128), .B(KEYINPUT4), .ZN(n388) );
  XNOR2_X2 U505 ( .A(n467), .B(G134), .ZN(n389) );
  INV_X1 U506 ( .A(n422), .ZN(n397) );
  NAND2_X1 U507 ( .A1(n393), .A2(n602), .ZN(n624) );
  NAND2_X1 U508 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U509 ( .A1(n396), .A2(n397), .ZN(n394) );
  AND2_X1 U510 ( .A1(n687), .A2(KEYINPUT104), .ZN(n396) );
  AND2_X1 U511 ( .A1(n400), .A2(n398), .ZN(n395) );
  NAND2_X1 U512 ( .A1(n399), .A2(n401), .ZN(n398) );
  NAND2_X1 U513 ( .A1(n422), .A2(n401), .ZN(n400) );
  INV_X1 U514 ( .A(KEYINPUT48), .ZN(n402) );
  NAND2_X1 U515 ( .A1(n404), .A2(n643), .ZN(n403) );
  NAND2_X1 U516 ( .A1(n369), .A2(n642), .ZN(n405) );
  XNOR2_X2 U517 ( .A(n407), .B(G472), .ZN(n603) );
  XNOR2_X1 U518 ( .A(n505), .B(n476), .ZN(n673) );
  XNOR2_X2 U519 ( .A(G110), .B(KEYINPUT88), .ZN(n721) );
  XNOR2_X2 U520 ( .A(n410), .B(n409), .ZN(n611) );
  NAND2_X1 U521 ( .A1(n419), .A2(n418), .ZN(n417) );
  XNOR2_X1 U522 ( .A(n417), .B(n375), .ZN(G57) );
  XNOR2_X2 U523 ( .A(n620), .B(KEYINPUT40), .ZN(n751) );
  XNOR2_X2 U524 ( .A(n411), .B(n374), .ZN(n664) );
  NAND2_X1 U525 ( .A1(n412), .A2(n430), .ZN(n411) );
  XNOR2_X1 U526 ( .A(n413), .B(KEYINPUT44), .ZN(n412) );
  XNOR2_X2 U527 ( .A(n462), .B(n428), .ZN(n633) );
  INV_X1 U528 ( .A(n557), .ZN(n561) );
  NAND2_X1 U529 ( .A1(n557), .A2(n368), .ZN(n414) );
  XNOR2_X2 U530 ( .A(n543), .B(KEYINPUT0), .ZN(n557) );
  NAND2_X1 U531 ( .A1(n423), .A2(n579), .ZN(n422) );
  INV_X1 U532 ( .A(n585), .ZN(n423) );
  NOR2_X2 U533 ( .A1(G902), .A2(n700), .ZN(n508) );
  XOR2_X1 U534 ( .A(n699), .B(n698), .Z(n427) );
  AND2_X1 U535 ( .A1(G210), .A2(n461), .ZN(n428) );
  AND2_X1 U536 ( .A1(G214), .A2(n470), .ZN(n429) );
  AND2_X1 U537 ( .A1(n568), .A2(n677), .ZN(n430) );
  XNOR2_X1 U538 ( .A(KEYINPUT46), .B(KEYINPUT64), .ZN(n621) );
  INV_X1 U539 ( .A(KEYINPUT17), .ZN(n452) );
  XNOR2_X1 U540 ( .A(n472), .B(n471), .ZN(n475) );
  XNOR2_X1 U541 ( .A(n455), .B(n454), .ZN(n458) );
  XNOR2_X1 U542 ( .A(n475), .B(n474), .ZN(n476) );
  INV_X1 U543 ( .A(KEYINPUT83), .ZN(n569) );
  INV_X1 U544 ( .A(G469), .ZN(n507) );
  XNOR2_X1 U545 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U546 ( .A(n700), .B(n427), .ZN(n701) );
  XOR2_X1 U547 ( .A(KEYINPUT14), .B(n431), .Z(n571) );
  XNOR2_X1 U548 ( .A(KEYINPUT99), .B(G478), .ZN(n437) );
  XNOR2_X1 U549 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n435) );
  XOR2_X1 U550 ( .A(G143), .B(G128), .Z(n432) );
  NAND2_X1 U551 ( .A1(G217), .A2(n485), .ZN(n433) );
  XOR2_X1 U552 ( .A(G116), .B(G107), .Z(n446) );
  NOR2_X1 U553 ( .A1(G902), .A2(n710), .ZN(n436) );
  XOR2_X1 U554 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n439) );
  XNOR2_X1 U555 ( .A(G140), .B(KEYINPUT95), .ZN(n438) );
  XOR2_X1 U556 ( .A(n439), .B(n438), .Z(n441) );
  XOR2_X1 U557 ( .A(G122), .B(G104), .Z(n445) );
  XNOR2_X1 U558 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n442) );
  NOR2_X1 U559 ( .A1(n550), .A2(n551), .ZN(n528) );
  INV_X1 U560 ( .A(n528), .ZN(n544) );
  OR2_X1 U561 ( .A1(G237), .A2(G902), .ZN(n461) );
  NAND2_X1 U562 ( .A1(G214), .A2(n461), .ZN(n602) );
  XOR2_X1 U563 ( .A(n446), .B(n445), .Z(n450) );
  XOR2_X2 U564 ( .A(G101), .B(G113), .Z(n448) );
  XNOR2_X2 U565 ( .A(n448), .B(n447), .ZN(n472) );
  XNOR2_X1 U566 ( .A(n472), .B(KEYINPUT16), .ZN(n449) );
  XNOR2_X1 U567 ( .A(n449), .B(n450), .ZN(n719) );
  XNOR2_X1 U568 ( .A(n719), .B(n467), .ZN(n460) );
  INV_X1 U569 ( .A(KEYINPUT18), .ZN(n451) );
  XNOR2_X1 U570 ( .A(n451), .B(n500), .ZN(n455) );
  NAND2_X1 U571 ( .A1(G224), .A2(n737), .ZN(n453) );
  XNOR2_X1 U572 ( .A(n456), .B(KEYINPUT89), .ZN(n457) );
  XNOR2_X1 U573 ( .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U574 ( .A(n661), .ZN(n491) );
  NAND2_X1 U575 ( .A1(n658), .A2(n491), .ZN(n462) );
  XNOR2_X1 U576 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n463) );
  NAND2_X1 U577 ( .A1(n602), .A2(n601), .ZN(n525) );
  XNOR2_X1 U578 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n464) );
  INV_X1 U579 ( .A(n468), .ZN(n469) );
  NAND2_X1 U580 ( .A1(n470), .A2(G210), .ZN(n471) );
  XOR2_X1 U581 ( .A(n473), .B(KEYINPUT5), .Z(n474) );
  INV_X1 U582 ( .A(n603), .ZN(n586) );
  NAND2_X1 U583 ( .A1(n477), .A2(n501), .ZN(n481) );
  INV_X1 U584 ( .A(n501), .ZN(n478) );
  NAND2_X1 U585 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U586 ( .A1(n481), .A2(n480), .ZN(n732) );
  XNOR2_X1 U587 ( .A(n732), .B(KEYINPUT91), .ZN(n488) );
  XNOR2_X1 U588 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U589 ( .A(n484), .B(KEYINPUT23), .Z(n486) );
  XNOR2_X1 U590 ( .A(KEYINPUT76), .B(KEYINPUT25), .ZN(n490) );
  INV_X1 U591 ( .A(KEYINPUT92), .ZN(n489) );
  XOR2_X1 U592 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n493) );
  NAND2_X1 U593 ( .A1(G234), .A2(n491), .ZN(n492) );
  XNOR2_X1 U594 ( .A(n493), .B(n492), .ZN(n495) );
  NAND2_X1 U595 ( .A1(n495), .A2(G217), .ZN(n494) );
  NAND2_X1 U596 ( .A1(n495), .A2(G221), .ZN(n496) );
  XNOR2_X1 U597 ( .A(n496), .B(KEYINPUT21), .ZN(n608) );
  NAND2_X1 U598 ( .A1(G227), .A2(n737), .ZN(n497) );
  XNOR2_X1 U599 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U600 ( .A(G101), .B(n499), .ZN(n504) );
  XNOR2_X1 U601 ( .A(n501), .B(G104), .ZN(n502) );
  XNOR2_X2 U602 ( .A(n508), .B(n507), .ZN(n606) );
  NOR2_X1 U603 ( .A1(n586), .A2(n520), .ZN(n556) );
  NOR2_X1 U604 ( .A1(n559), .A2(n362), .ZN(n510) );
  XNOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT113), .ZN(n509) );
  XNOR2_X1 U606 ( .A(n510), .B(n509), .ZN(n514) );
  XOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n512) );
  NAND2_X1 U608 ( .A1(n608), .A2(n611), .ZN(n511) );
  XNOR2_X1 U609 ( .A(n512), .B(n511), .ZN(n513) );
  NAND2_X1 U610 ( .A1(n514), .A2(n513), .ZN(n515) );
  NOR2_X1 U611 ( .A1(n603), .A2(n515), .ZN(n516) );
  XNOR2_X1 U612 ( .A(n516), .B(KEYINPUT114), .ZN(n517) );
  NOR2_X1 U613 ( .A1(n556), .A2(n517), .ZN(n518) );
  XOR2_X1 U614 ( .A(KEYINPUT51), .B(n518), .Z(n519) );
  NOR2_X1 U615 ( .A1(n653), .A2(n519), .ZN(n534) );
  XNOR2_X2 U616 ( .A(n522), .B(KEYINPUT33), .ZN(n652) );
  XNOR2_X1 U617 ( .A(KEYINPUT97), .B(n551), .ZN(n524) );
  NAND2_X1 U618 ( .A1(n524), .A2(n550), .ZN(n523) );
  INV_X1 U619 ( .A(n592), .ZN(n636) );
  NOR2_X1 U620 ( .A1(n636), .A2(n525), .ZN(n526) );
  XNOR2_X1 U621 ( .A(n526), .B(KEYINPUT115), .ZN(n530) );
  OR2_X1 U622 ( .A1(n602), .A2(n601), .ZN(n527) );
  NAND2_X1 U623 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U624 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U625 ( .A1(n652), .A2(n531), .ZN(n532) );
  XOR2_X1 U626 ( .A(KEYINPUT116), .B(n532), .Z(n533) );
  NOR2_X1 U627 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U628 ( .A(n535), .B(KEYINPUT52), .ZN(n536) );
  NOR2_X1 U629 ( .A1(n571), .A2(n536), .ZN(n537) );
  NAND2_X1 U630 ( .A1(G952), .A2(n537), .ZN(n651) );
  INV_X1 U631 ( .A(n362), .ZN(n628) );
  NOR2_X1 U632 ( .A1(n579), .A2(n628), .ZN(n538) );
  NAND2_X1 U633 ( .A1(n611), .A2(n538), .ZN(n539) );
  XNOR2_X1 U634 ( .A(KEYINPUT79), .B(n539), .ZN(n547) );
  NAND2_X1 U635 ( .A1(n633), .A2(n602), .ZN(n540) );
  XNOR2_X1 U636 ( .A(n540), .B(KEYINPUT19), .ZN(n584) );
  NAND2_X1 U637 ( .A1(G952), .A2(n737), .ZN(n574) );
  NOR2_X1 U638 ( .A1(G898), .A2(n737), .ZN(n722) );
  NAND2_X1 U639 ( .A1(G902), .A2(n722), .ZN(n541) );
  NAND2_X1 U640 ( .A1(n574), .A2(n541), .ZN(n542) );
  OR2_X1 U641 ( .A1(n544), .A2(n608), .ZN(n545) );
  XOR2_X1 U642 ( .A(KEYINPUT22), .B(KEYINPUT65), .Z(n546) );
  NAND2_X1 U643 ( .A1(n547), .A2(n553), .ZN(n548) );
  XOR2_X1 U644 ( .A(KEYINPUT32), .B(n548), .Z(n750) );
  NAND2_X1 U645 ( .A1(n652), .A2(n557), .ZN(n549) );
  NAND2_X1 U646 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U647 ( .A(KEYINPUT103), .B(n552), .Z(n632) );
  NAND2_X1 U648 ( .A1(n553), .A2(n628), .ZN(n565) );
  NOR2_X1 U649 ( .A1(n603), .A2(n565), .ZN(n554) );
  NAND2_X1 U650 ( .A1(n611), .A2(n554), .ZN(n683) );
  NAND2_X1 U651 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U652 ( .A(KEYINPUT31), .B(n558), .Z(n691) );
  NAND2_X1 U653 ( .A1(n606), .A2(n559), .ZN(n560) );
  NOR2_X1 U654 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U655 ( .A1(n562), .A2(n586), .ZN(n679) );
  NAND2_X1 U656 ( .A1(n691), .A2(n679), .ZN(n563) );
  XNOR2_X1 U657 ( .A(n563), .B(KEYINPUT94), .ZN(n564) );
  NAND2_X1 U658 ( .A1(n564), .A2(n592), .ZN(n568) );
  NOR2_X1 U659 ( .A1(n611), .A2(n565), .ZN(n567) );
  INV_X1 U660 ( .A(n579), .ZN(n566) );
  NAND2_X1 U661 ( .A1(n567), .A2(n566), .ZN(n677) );
  INV_X1 U662 ( .A(n361), .ZN(n727) );
  XNOR2_X1 U663 ( .A(n570), .B(KEYINPUT82), .ZN(n647) );
  INV_X1 U664 ( .A(n571), .ZN(n576) );
  NOR2_X1 U665 ( .A1(G900), .A2(n737), .ZN(n572) );
  NAND2_X1 U666 ( .A1(G902), .A2(n572), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U668 ( .A1(n576), .A2(n575), .ZN(n605) );
  NOR2_X1 U669 ( .A1(n608), .A2(n605), .ZN(n577) );
  XNOR2_X1 U670 ( .A(KEYINPUT68), .B(n577), .ZN(n578) );
  NOR2_X1 U671 ( .A1(n362), .A2(n624), .ZN(n581) );
  XNOR2_X1 U672 ( .A(n581), .B(KEYINPUT43), .ZN(n582) );
  NOR2_X1 U673 ( .A1(n633), .A2(n582), .ZN(n696) );
  INV_X1 U674 ( .A(KEYINPUT80), .ZN(n639) );
  NOR2_X1 U675 ( .A1(n592), .A2(n639), .ZN(n583) );
  NOR2_X1 U676 ( .A1(KEYINPUT73), .A2(n583), .ZN(n590) );
  INV_X1 U677 ( .A(n584), .ZN(n589) );
  XNOR2_X1 U678 ( .A(KEYINPUT28), .B(n587), .ZN(n588) );
  NAND2_X1 U679 ( .A1(n588), .A2(n606), .ZN(n598) );
  NOR2_X1 U680 ( .A1(n589), .A2(n598), .ZN(n688) );
  NAND2_X1 U681 ( .A1(n590), .A2(n688), .ZN(n591) );
  NAND2_X1 U682 ( .A1(n591), .A2(KEYINPUT47), .ZN(n597) );
  INV_X1 U683 ( .A(KEYINPUT73), .ZN(n593) );
  INV_X1 U684 ( .A(KEYINPUT47), .ZN(n594) );
  NAND2_X1 U685 ( .A1(n595), .A2(n688), .ZN(n596) );
  XNOR2_X1 U686 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n599) );
  INV_X1 U687 ( .A(n601), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U689 ( .A(KEYINPUT30), .B(n604), .Z(n614) );
  INV_X1 U690 ( .A(n605), .ZN(n607) );
  AND2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n610) );
  INV_X1 U692 ( .A(n608), .ZN(n609) );
  NAND2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n631) );
  XNOR2_X1 U695 ( .A(KEYINPUT70), .B(KEYINPUT84), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n619), .B(n618), .ZN(n644) );
  NAND2_X1 U697 ( .A1(n644), .A2(n687), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n752), .A2(n751), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(n626), .ZN(n629) );
  NOR2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U703 ( .A(n630), .B(KEYINPUT108), .ZN(n748) );
  INV_X1 U704 ( .A(n748), .ZN(n643) );
  NOR2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U707 ( .A(KEYINPUT105), .B(n635), .Z(n747) );
  NAND2_X1 U708 ( .A1(n636), .A2(KEYINPUT47), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n747), .A2(n637), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U711 ( .A1(n747), .A2(KEYINPUT80), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n642) );
  INV_X1 U713 ( .A(n692), .ZN(n684) );
  NAND2_X1 U714 ( .A1(n644), .A2(n684), .ZN(n695) );
  INV_X1 U715 ( .A(n736), .ZN(n645) );
  NOR2_X1 U716 ( .A1(KEYINPUT2), .A2(n645), .ZN(n646) );
  NOR2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n649) );
  NOR2_X1 U718 ( .A1(n664), .A2(n736), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n649), .A2(n662), .ZN(n650) );
  INV_X1 U720 ( .A(n652), .ZN(n654) );
  NOR2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U722 ( .A(KEYINPUT117), .B(n655), .Z(n656) );
  NOR2_X1 U723 ( .A1(G952), .A2(n737), .ZN(n657) );
  XOR2_X1 U724 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n660) );
  XNOR2_X1 U725 ( .A(n360), .B(KEYINPUT81), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n662), .A2(n661), .ZN(n668) );
  INV_X1 U727 ( .A(KEYINPUT75), .ZN(n663) );
  NOR2_X1 U728 ( .A1(KEYINPUT2), .A2(n666), .ZN(n667) );
  NAND2_X1 U729 ( .A1(n705), .A2(G210), .ZN(n669) );
  XNOR2_X1 U730 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U731 ( .A(KEYINPUT56), .B(KEYINPUT118), .ZN(n672) );
  XOR2_X1 U732 ( .A(n673), .B(KEYINPUT62), .Z(n674) );
  XNOR2_X1 U733 ( .A(n674), .B(KEYINPUT86), .ZN(n675) );
  XNOR2_X1 U734 ( .A(G101), .B(n677), .ZN(G3) );
  NOR2_X1 U735 ( .A1(n399), .A2(n679), .ZN(n678) );
  XOR2_X1 U736 ( .A(G104), .B(n678), .Z(G6) );
  NOR2_X1 U737 ( .A1(n692), .A2(n679), .ZN(n681) );
  XNOR2_X1 U738 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n680) );
  XNOR2_X1 U739 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U740 ( .A(G107), .B(n682), .ZN(G9) );
  XNOR2_X1 U741 ( .A(G110), .B(n683), .ZN(G12) );
  XOR2_X1 U742 ( .A(G128), .B(KEYINPUT29), .Z(n686) );
  NAND2_X1 U743 ( .A1(n688), .A2(n684), .ZN(n685) );
  XNOR2_X1 U744 ( .A(n686), .B(n685), .ZN(G30) );
  NAND2_X1 U745 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n689), .B(G146), .ZN(G48) );
  NOR2_X1 U747 ( .A1(n399), .A2(n691), .ZN(n690) );
  XOR2_X1 U748 ( .A(G113), .B(n690), .Z(G15) );
  NOR2_X1 U749 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U750 ( .A(KEYINPUT110), .B(n693), .Z(n694) );
  XNOR2_X1 U751 ( .A(G116), .B(n694), .ZN(G18) );
  XNOR2_X1 U752 ( .A(G134), .B(n695), .ZN(G36) );
  XNOR2_X1 U753 ( .A(G140), .B(n696), .ZN(n697) );
  XNOR2_X1 U754 ( .A(n697), .B(KEYINPUT111), .ZN(G42) );
  BUF_X1 U755 ( .A(n705), .Z(n714) );
  NAND2_X1 U756 ( .A1(n714), .A2(G469), .ZN(n702) );
  XOR2_X1 U757 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n699) );
  XNOR2_X1 U758 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n698) );
  NOR2_X1 U759 ( .A1(n718), .A2(n703), .ZN(G54) );
  NAND2_X1 U760 ( .A1(n705), .A2(G475), .ZN(n706) );
  XNOR2_X1 U761 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U762 ( .A(n709), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U763 ( .A(n710), .B(KEYINPUT121), .Z(n712) );
  NAND2_X1 U764 ( .A1(n714), .A2(G478), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n718), .A2(n713), .ZN(G63) );
  NAND2_X1 U767 ( .A1(G217), .A2(n714), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n718), .A2(n717), .ZN(G66) );
  XOR2_X1 U770 ( .A(n719), .B(KEYINPUT123), .Z(n720) );
  XNOR2_X1 U771 ( .A(n721), .B(n720), .ZN(n723) );
  NOR2_X1 U772 ( .A1(n723), .A2(n722), .ZN(n731) );
  NAND2_X1 U773 ( .A1(G224), .A2(G953), .ZN(n724) );
  XNOR2_X1 U774 ( .A(n724), .B(KEYINPUT61), .ZN(n725) );
  XNOR2_X1 U775 ( .A(KEYINPUT122), .B(n725), .ZN(n726) );
  NAND2_X1 U776 ( .A1(G898), .A2(n726), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n727), .A2(n737), .ZN(n728) );
  NAND2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U779 ( .A(n731), .B(n730), .ZN(G69) );
  XNOR2_X1 U780 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n735) );
  XNOR2_X1 U781 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n735), .B(n734), .ZN(n740) );
  XNOR2_X1 U783 ( .A(n740), .B(n736), .ZN(n738) );
  NAND2_X1 U784 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U785 ( .A(KEYINPUT126), .B(n739), .ZN(n745) );
  XNOR2_X1 U786 ( .A(G227), .B(n740), .ZN(n741) );
  NAND2_X1 U787 ( .A1(n741), .A2(G900), .ZN(n742) );
  NAND2_X1 U788 ( .A1(n742), .A2(G953), .ZN(n743) );
  XOR2_X1 U789 ( .A(KEYINPUT127), .B(n743), .Z(n744) );
  NAND2_X1 U790 ( .A1(n745), .A2(n744), .ZN(G72) );
  XNOR2_X1 U791 ( .A(n746), .B(G122), .ZN(G24) );
  XNOR2_X1 U792 ( .A(G143), .B(n747), .ZN(G45) );
  XNOR2_X1 U793 ( .A(G125), .B(KEYINPUT37), .ZN(n749) );
  XNOR2_X1 U794 ( .A(n749), .B(n748), .ZN(G27) );
  XOR2_X1 U795 ( .A(n750), .B(G119), .Z(G21) );
  XNOR2_X1 U796 ( .A(G131), .B(n751), .ZN(G33) );
  XNOR2_X1 U797 ( .A(G137), .B(n752), .ZN(G39) );
endmodule

