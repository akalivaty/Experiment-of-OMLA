

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U549 ( .A1(n733), .A2(n732), .ZN(n740) );
  BUF_X1 U550 ( .A(n615), .Z(n616) );
  NOR2_X1 U551 ( .A1(G299), .A2(n709), .ZN(n695) );
  XNOR2_X2 U552 ( .A(n521), .B(n520), .ZN(n617) );
  XNOR2_X1 U553 ( .A(KEYINPUT93), .B(n810), .ZN(n513) );
  NOR2_X1 U554 ( .A1(n768), .A2(n915), .ZN(n514) );
  AND2_X1 U555 ( .A1(n764), .A2(n763), .ZN(n515) );
  OR2_X1 U556 ( .A1(n723), .A2(G301), .ZN(n516) );
  XOR2_X1 U557 ( .A(n699), .B(KEYINPUT26), .Z(n517) );
  XOR2_X1 U558 ( .A(n693), .B(KEYINPUT27), .Z(n518) );
  NOR2_X1 U559 ( .A1(n735), .A2(n970), .ZN(n699) );
  AND2_X1 U560 ( .A1(n794), .A2(n795), .ZN(n696) );
  NOR2_X1 U561 ( .A1(n703), .A2(n702), .ZN(n706) );
  INV_X1 U562 ( .A(KEYINPUT97), .ZN(n741) );
  XNOR2_X1 U563 ( .A(n744), .B(KEYINPUT32), .ZN(n745) );
  INV_X1 U564 ( .A(KEYINPUT86), .ZN(n691) );
  NOR2_X1 U565 ( .A1(G2105), .A2(n524), .ZN(n531) );
  NOR2_X1 U566 ( .A1(G164), .A2(G1384), .ZN(n795) );
  INV_X1 U567 ( .A(KEYINPUT23), .ZN(n532) );
  NAND2_X1 U568 ( .A1(n513), .A2(n811), .ZN(n812) );
  XNOR2_X1 U569 ( .A(n533), .B(n532), .ZN(n534) );
  NOR2_X1 U570 ( .A1(G651), .A2(n649), .ZN(n654) );
  NOR2_X1 U571 ( .A1(n539), .A2(n538), .ZN(n690) );
  BUF_X1 U572 ( .A(n690), .Z(G160) );
  INV_X1 U573 ( .A(G2104), .ZN(n524) );
  INV_X1 U574 ( .A(n531), .ZN(n519) );
  INV_X1 U575 ( .A(n519), .ZN(n889) );
  NAND2_X1 U576 ( .A1(G102), .A2(n889), .ZN(n523) );
  XNOR2_X1 U577 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n521) );
  NOR2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  NAND2_X1 U579 ( .A1(G138), .A2(n617), .ZN(n522) );
  NAND2_X1 U580 ( .A1(n523), .A2(n522), .ZN(n529) );
  INV_X1 U581 ( .A(G2105), .ZN(n525) );
  NOR2_X1 U582 ( .A1(n524), .A2(n525), .ZN(n615) );
  NAND2_X1 U583 ( .A1(G114), .A2(n615), .ZN(n527) );
  NOR2_X2 U584 ( .A1(G2104), .A2(n525), .ZN(n885) );
  NAND2_X1 U585 ( .A1(G126), .A2(n885), .ZN(n526) );
  NAND2_X1 U586 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U587 ( .A1(n529), .A2(n528), .ZN(G164) );
  NAND2_X1 U588 ( .A1(G113), .A2(n615), .ZN(n530) );
  XNOR2_X1 U589 ( .A(n530), .B(KEYINPUT64), .ZN(n535) );
  NAND2_X1 U590 ( .A1(G101), .A2(n531), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U592 ( .A1(G125), .A2(n885), .ZN(n537) );
  NAND2_X1 U593 ( .A1(G137), .A2(n617), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n661) );
  NAND2_X1 U596 ( .A1(G91), .A2(n661), .ZN(n542) );
  INV_X1 U597 ( .A(G651), .ZN(n543) );
  NOR2_X1 U598 ( .A1(G543), .A2(n543), .ZN(n540) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n540), .Z(n653) );
  NAND2_X1 U600 ( .A1(G65), .A2(n653), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n547) );
  XOR2_X1 U602 ( .A(KEYINPUT0), .B(G543), .Z(n649) );
  NOR2_X1 U603 ( .A1(n649), .A2(n543), .ZN(n658) );
  NAND2_X1 U604 ( .A1(G78), .A2(n658), .ZN(n545) );
  NAND2_X1 U605 ( .A1(G53), .A2(n654), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U607 ( .A1(n547), .A2(n546), .ZN(G299) );
  NAND2_X1 U608 ( .A1(n661), .A2(G89), .ZN(n548) );
  XNOR2_X1 U609 ( .A(n548), .B(KEYINPUT4), .ZN(n550) );
  NAND2_X1 U610 ( .A1(G76), .A2(n658), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U612 ( .A(KEYINPUT5), .B(n551), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n654), .A2(G51), .ZN(n552) );
  XOR2_X1 U614 ( .A(KEYINPUT75), .B(n552), .Z(n554) );
  NAND2_X1 U615 ( .A1(n653), .A2(G63), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n555), .Z(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U619 ( .A(KEYINPUT7), .B(n558), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(n559) );
  XNOR2_X1 U621 ( .A(KEYINPUT76), .B(n559), .ZN(G286) );
  XOR2_X1 U622 ( .A(G2446), .B(G2451), .Z(n561) );
  XNOR2_X1 U623 ( .A(G2454), .B(KEYINPUT105), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n561), .B(n560), .ZN(n568) );
  XOR2_X1 U625 ( .A(G2438), .B(G2430), .Z(n563) );
  XNOR2_X1 U626 ( .A(G2435), .B(G2443), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U628 ( .A(n564), .B(G2427), .Z(n566) );
  XNOR2_X1 U629 ( .A(G1341), .B(G1348), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U631 ( .A(n568), .B(n567), .ZN(n569) );
  AND2_X1 U632 ( .A1(n569), .A2(G14), .ZN(G401) );
  AND2_X1 U633 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U634 ( .A(G132), .ZN(G219) );
  INV_X1 U635 ( .A(G69), .ZN(G235) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n829) );
  NAND2_X1 U639 ( .A1(n829), .A2(G567), .ZN(n571) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  NAND2_X1 U641 ( .A1(G56), .A2(n653), .ZN(n572) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(n572), .Z(n578) );
  NAND2_X1 U643 ( .A1(n661), .A2(G81), .ZN(n573) );
  XNOR2_X1 U644 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U645 ( .A1(G68), .A2(n658), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n654), .A2(G43), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n924) );
  INV_X1 U651 ( .A(G860), .ZN(n833) );
  XNOR2_X1 U652 ( .A(KEYINPUT72), .B(n833), .ZN(n603) );
  NOR2_X1 U653 ( .A1(n924), .A2(n603), .ZN(n581) );
  XNOR2_X1 U654 ( .A(n581), .B(KEYINPUT73), .ZN(G153) );
  NAND2_X1 U655 ( .A1(n658), .A2(G77), .ZN(n582) );
  XNOR2_X1 U656 ( .A(n582), .B(KEYINPUT70), .ZN(n584) );
  NAND2_X1 U657 ( .A1(G90), .A2(n661), .ZN(n583) );
  NAND2_X1 U658 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U659 ( .A(n585), .B(KEYINPUT9), .ZN(n587) );
  NAND2_X1 U660 ( .A1(G52), .A2(n654), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U662 ( .A1(G64), .A2(n653), .ZN(n588) );
  XNOR2_X1 U663 ( .A(KEYINPUT69), .B(n588), .ZN(n589) );
  NOR2_X1 U664 ( .A1(n590), .A2(n589), .ZN(G171) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G79), .A2(n658), .ZN(n592) );
  NAND2_X1 U667 ( .A1(G54), .A2(n654), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G92), .A2(n661), .ZN(n594) );
  NAND2_X1 U670 ( .A1(G66), .A2(n653), .ZN(n593) );
  NAND2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n597), .B(KEYINPUT15), .ZN(n840) );
  NOR2_X1 U674 ( .A1(G868), .A2(n840), .ZN(n599) );
  INV_X1 U675 ( .A(G868), .ZN(n673) );
  NOR2_X1 U676 ( .A1(n673), .A2(G301), .ZN(n598) );
  NOR2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U678 ( .A(KEYINPUT74), .B(n600), .ZN(G284) );
  NAND2_X1 U679 ( .A1(G868), .A2(G286), .ZN(n602) );
  NAND2_X1 U680 ( .A1(G299), .A2(n673), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U682 ( .A1(G559), .A2(n603), .ZN(n604) );
  XOR2_X1 U683 ( .A(KEYINPUT77), .B(n604), .Z(n605) );
  INV_X1 U684 ( .A(n840), .ZN(n917) );
  NAND2_X1 U685 ( .A1(n605), .A2(n917), .ZN(n606) );
  XNOR2_X1 U686 ( .A(n606), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n924), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n917), .A2(G868), .ZN(n607) );
  NOR2_X1 U689 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U690 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G123), .A2(n885), .ZN(n610) );
  XNOR2_X1 U692 ( .A(n610), .B(KEYINPUT78), .ZN(n611) );
  XNOR2_X1 U693 ( .A(KEYINPUT18), .B(n611), .ZN(n614) );
  NAND2_X1 U694 ( .A1(G99), .A2(n889), .ZN(n612) );
  XOR2_X1 U695 ( .A(KEYINPUT79), .B(n612), .Z(n613) );
  NAND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G111), .A2(n616), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G135), .A2(n617), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n946) );
  XNOR2_X1 U701 ( .A(n946), .B(G2096), .ZN(n623) );
  INV_X1 U702 ( .A(G2100), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G85), .A2(n661), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G72), .A2(n658), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U707 ( .A(KEYINPUT66), .B(n626), .Z(n632) );
  NAND2_X1 U708 ( .A1(n653), .A2(G60), .ZN(n627) );
  XOR2_X1 U709 ( .A(KEYINPUT67), .B(n627), .Z(n629) );
  NAND2_X1 U710 ( .A1(n654), .A2(G47), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U712 ( .A(KEYINPUT68), .B(n630), .Z(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(G290) );
  NAND2_X1 U714 ( .A1(G88), .A2(n661), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G75), .A2(n658), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G62), .A2(n653), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G50), .A2(n654), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U720 ( .A1(n638), .A2(n637), .ZN(G166) );
  NAND2_X1 U721 ( .A1(G86), .A2(n661), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G61), .A2(n653), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n658), .A2(G73), .ZN(n641) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n641), .Z(n642) );
  NOR2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n654), .A2(G48), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U729 ( .A1(G49), .A2(n654), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U732 ( .A1(n653), .A2(n648), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n649), .A2(G87), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n651), .A2(n650), .ZN(G288) );
  NAND2_X1 U735 ( .A1(G559), .A2(n917), .ZN(n652) );
  XOR2_X1 U736 ( .A(n924), .B(n652), .Z(n834) );
  NAND2_X1 U737 ( .A1(G67), .A2(n653), .ZN(n656) );
  NAND2_X1 U738 ( .A1(G55), .A2(n654), .ZN(n655) );
  NAND2_X1 U739 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U740 ( .A(n657), .B(KEYINPUT81), .ZN(n660) );
  NAND2_X1 U741 ( .A1(G80), .A2(n658), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n661), .A2(G93), .ZN(n662) );
  XOR2_X1 U744 ( .A(KEYINPUT80), .B(n662), .Z(n663) );
  NOR2_X1 U745 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U746 ( .A(KEYINPUT82), .B(n665), .Z(n836) );
  XNOR2_X1 U747 ( .A(n836), .B(G290), .ZN(n668) );
  XNOR2_X1 U748 ( .A(G166), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U749 ( .A(n666), .B(G305), .ZN(n667) );
  XNOR2_X1 U750 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U751 ( .A(n669), .B(G288), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n670), .B(G299), .ZN(n839) );
  XNOR2_X1 U753 ( .A(n834), .B(n839), .ZN(n671) );
  XNOR2_X1 U754 ( .A(KEYINPUT83), .B(n671), .ZN(n672) );
  NOR2_X1 U755 ( .A1(n673), .A2(n672), .ZN(n675) );
  NOR2_X1 U756 ( .A1(n836), .A2(G868), .ZN(n674) );
  NOR2_X1 U757 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n676) );
  XNOR2_X1 U760 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U761 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U762 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U763 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U764 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U765 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NAND2_X1 U766 ( .A1(G120), .A2(G108), .ZN(n681) );
  NOR2_X1 U767 ( .A1(G235), .A2(n681), .ZN(n682) );
  NAND2_X1 U768 ( .A1(n682), .A2(G57), .ZN(n683) );
  XOR2_X1 U769 ( .A(KEYINPUT85), .B(n683), .Z(n837) );
  NAND2_X1 U770 ( .A1(n837), .A2(G567), .ZN(n688) );
  NOR2_X1 U771 ( .A1(G219), .A2(G220), .ZN(n684) );
  XOR2_X1 U772 ( .A(KEYINPUT22), .B(n684), .Z(n685) );
  NOR2_X1 U773 ( .A1(G218), .A2(n685), .ZN(n686) );
  NAND2_X1 U774 ( .A1(G96), .A2(n686), .ZN(n838) );
  NAND2_X1 U775 ( .A1(n838), .A2(G2106), .ZN(n687) );
  NAND2_X1 U776 ( .A1(n688), .A2(n687), .ZN(n913) );
  NAND2_X1 U777 ( .A1(G661), .A2(G483), .ZN(n689) );
  NOR2_X1 U778 ( .A1(n913), .A2(n689), .ZN(n832) );
  NAND2_X1 U779 ( .A1(n832), .A2(G36), .ZN(G176) );
  INV_X1 U780 ( .A(G166), .ZN(G303) );
  NAND2_X1 U781 ( .A1(G40), .A2(n690), .ZN(n692) );
  XNOR2_X2 U782 ( .A(n692), .B(n691), .ZN(n794) );
  NAND2_X2 U783 ( .A1(n795), .A2(n794), .ZN(n735) );
  NOR2_X1 U784 ( .A1(G2084), .A2(n735), .ZN(n717) );
  NAND2_X1 U785 ( .A1(n717), .A2(G8), .ZN(n731) );
  NAND2_X1 U786 ( .A1(G8), .A2(n735), .ZN(n734) );
  NOR2_X1 U787 ( .A1(G1966), .A2(n734), .ZN(n718) );
  NAND2_X1 U788 ( .A1(n696), .A2(G2072), .ZN(n693) );
  NAND2_X1 U789 ( .A1(G1956), .A2(n735), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n518), .A2(n694), .ZN(n709) );
  XNOR2_X1 U791 ( .A(n695), .B(KEYINPUT94), .ZN(n708) );
  NAND2_X1 U792 ( .A1(G1348), .A2(n735), .ZN(n698) );
  NAND2_X1 U793 ( .A1(G2067), .A2(n696), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n704) );
  NOR2_X1 U795 ( .A1(n840), .A2(n704), .ZN(n703) );
  INV_X1 U796 ( .A(G1996), .ZN(n970) );
  NAND2_X1 U797 ( .A1(n735), .A2(G1341), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n517), .A2(n700), .ZN(n701) );
  NOR2_X1 U799 ( .A1(n701), .A2(n924), .ZN(n702) );
  AND2_X1 U800 ( .A1(n840), .A2(n704), .ZN(n705) );
  NOR2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U803 ( .A1(G299), .A2(n709), .ZN(n710) );
  XOR2_X1 U804 ( .A(KEYINPUT28), .B(n710), .Z(n711) );
  NOR2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U806 ( .A(n713), .B(KEYINPUT29), .ZN(n716) );
  XOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .Z(n975) );
  NOR2_X1 U808 ( .A1(n975), .A2(n735), .ZN(n715) );
  NOR2_X1 U809 ( .A1(n696), .A2(G1961), .ZN(n714) );
  NOR2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n723) );
  AND2_X1 U811 ( .A1(n716), .A2(n516), .ZN(n728) );
  NOR2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U813 ( .A1(G8), .A2(n719), .ZN(n720) );
  XNOR2_X1 U814 ( .A(KEYINPUT30), .B(n720), .ZN(n721) );
  XOR2_X1 U815 ( .A(KEYINPUT95), .B(n721), .Z(n722) );
  NOR2_X1 U816 ( .A1(G168), .A2(n722), .ZN(n725) );
  AND2_X1 U817 ( .A1(G301), .A2(n723), .ZN(n724) );
  NOR2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U819 ( .A(n726), .B(KEYINPUT31), .ZN(n727) );
  NOR2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U821 ( .A(n729), .B(KEYINPUT96), .ZN(n733) );
  NOR2_X1 U822 ( .A1(n718), .A2(n733), .ZN(n730) );
  NAND2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n748) );
  INV_X1 U824 ( .A(G286), .ZN(n732) );
  INV_X1 U825 ( .A(n734), .ZN(n761) );
  INV_X1 U826 ( .A(n761), .ZN(n773) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n773), .ZN(n737) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U830 ( .A1(n738), .A2(G303), .ZN(n739) );
  NAND2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U832 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n743), .A2(G8), .ZN(n746) );
  XOR2_X1 U834 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n744) );
  XNOR2_X1 U835 ( .A(n746), .B(n745), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U837 ( .A(n749), .B(KEYINPUT100), .ZN(n760) );
  NOR2_X1 U838 ( .A1(G2090), .A2(G303), .ZN(n750) );
  XNOR2_X1 U839 ( .A(KEYINPUT102), .B(n750), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n751), .A2(G8), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n760), .A2(n752), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n753), .A2(n773), .ZN(n755) );
  INV_X1 U843 ( .A(KEYINPUT103), .ZN(n754) );
  XNOR2_X1 U844 ( .A(n755), .B(n754), .ZN(n770) );
  NOR2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n756) );
  XOR2_X1 U846 ( .A(KEYINPUT101), .B(n756), .Z(n765) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n765), .A2(n757), .ZN(n928) );
  INV_X1 U849 ( .A(KEYINPUT33), .ZN(n758) );
  AND2_X1 U850 ( .A1(n928), .A2(n758), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n919) );
  AND2_X1 U853 ( .A1(n761), .A2(n919), .ZN(n762) );
  OR2_X1 U854 ( .A1(KEYINPUT33), .A2(n762), .ZN(n763) );
  INV_X1 U855 ( .A(n765), .ZN(n766) );
  NOR2_X1 U856 ( .A1(n766), .A2(n773), .ZN(n767) );
  AND2_X1 U857 ( .A1(KEYINPUT33), .A2(n767), .ZN(n768) );
  XNOR2_X1 U858 ( .A(G1981), .B(G305), .ZN(n915) );
  NAND2_X1 U859 ( .A1(n515), .A2(n514), .ZN(n769) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n775) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XOR2_X1 U862 ( .A(n771), .B(KEYINPUT24), .Z(n772) );
  NOR2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n813) );
  NAND2_X1 U865 ( .A1(n885), .A2(G119), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G131), .A2(n617), .ZN(n776) );
  XOR2_X1 U867 ( .A(KEYINPUT89), .B(n776), .Z(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U869 ( .A1(G107), .A2(n616), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G95), .A2(n889), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n901) );
  INV_X1 U873 ( .A(G1991), .ZN(n968) );
  NOR2_X1 U874 ( .A1(n901), .A2(n968), .ZN(n793) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(KEYINPUT91), .Z(n784) );
  NAND2_X1 U876 ( .A1(G105), .A2(n889), .ZN(n783) );
  XNOR2_X1 U877 ( .A(n784), .B(n783), .ZN(n785) );
  XNOR2_X1 U878 ( .A(n785), .B(KEYINPUT90), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n885), .A2(G129), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G117), .A2(n616), .ZN(n789) );
  NAND2_X1 U882 ( .A1(G141), .A2(n617), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n881) );
  NOR2_X1 U885 ( .A1(n881), .A2(n970), .ZN(n792) );
  NOR2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n943) );
  INV_X1 U887 ( .A(n794), .ZN(n796) );
  NOR2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n824) );
  INV_X1 U889 ( .A(n824), .ZN(n797) );
  NOR2_X1 U890 ( .A1(n943), .A2(n797), .ZN(n817) );
  XOR2_X1 U891 ( .A(KEYINPUT92), .B(n817), .Z(n809) );
  NAND2_X1 U892 ( .A1(G104), .A2(n889), .ZN(n799) );
  NAND2_X1 U893 ( .A1(G140), .A2(n617), .ZN(n798) );
  NAND2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U895 ( .A(n800), .B(KEYINPUT87), .ZN(n801) );
  XNOR2_X1 U896 ( .A(n801), .B(KEYINPUT34), .ZN(n807) );
  XNOR2_X1 U897 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n805) );
  NAND2_X1 U898 ( .A1(G116), .A2(n616), .ZN(n803) );
  NAND2_X1 U899 ( .A1(G128), .A2(n885), .ZN(n802) );
  NAND2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U901 ( .A(n805), .B(n804), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U903 ( .A(KEYINPUT36), .B(n808), .Z(n904) );
  XNOR2_X1 U904 ( .A(KEYINPUT37), .B(G2067), .ZN(n814) );
  NOR2_X1 U905 ( .A1(n904), .A2(n814), .ZN(n950) );
  NAND2_X1 U906 ( .A1(n824), .A2(n950), .ZN(n822) );
  NAND2_X1 U907 ( .A1(n809), .A2(n822), .ZN(n810) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n934) );
  NAND2_X1 U909 ( .A1(n934), .A2(n824), .ZN(n811) );
  OR2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n827) );
  NAND2_X1 U911 ( .A1(n904), .A2(n814), .ZN(n942) );
  AND2_X1 U912 ( .A1(n968), .A2(n901), .ZN(n947) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n815) );
  NOR2_X1 U914 ( .A1(n947), .A2(n815), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n818) );
  AND2_X1 U916 ( .A1(n970), .A2(n881), .ZN(n954) );
  NOR2_X1 U917 ( .A1(n818), .A2(n954), .ZN(n820) );
  XNOR2_X1 U918 ( .A(KEYINPUT104), .B(KEYINPUT39), .ZN(n819) );
  XNOR2_X1 U919 ( .A(n820), .B(n819), .ZN(n821) );
  NAND2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n942), .A2(n823), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U924 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U927 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(G188) );
  XOR2_X1 U930 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  XOR2_X1 U931 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  NAND2_X1 U933 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(G145) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  NOR2_X1 U936 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U938 ( .A(G171), .B(n839), .ZN(n843) );
  XNOR2_X1 U939 ( .A(KEYINPUT114), .B(n924), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n844), .B(G286), .ZN(n845) );
  NOR2_X1 U943 ( .A1(G37), .A2(n845), .ZN(G397) );
  XOR2_X1 U944 ( .A(G2100), .B(G2096), .Z(n847) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2090), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1961), .B(G1971), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1981), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U956 ( .A(G1966), .B(G1956), .Z(n857) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U960 ( .A(G2474), .B(KEYINPUT107), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U962 ( .A(G1976), .B(KEYINPUT41), .Z(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U964 ( .A1(n885), .A2(G124), .ZN(n865) );
  XNOR2_X1 U965 ( .A(KEYINPUT108), .B(KEYINPUT44), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n872) );
  NAND2_X1 U967 ( .A1(G112), .A2(n616), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G136), .A2(n617), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G100), .A2(n889), .ZN(n868) );
  XNOR2_X1 U971 ( .A(KEYINPUT109), .B(n868), .ZN(n869) );
  NOR2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U974 ( .A(KEYINPUT110), .B(n873), .Z(G162) );
  NAND2_X1 U975 ( .A1(G118), .A2(n616), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G130), .A2(n885), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G106), .A2(n889), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G142), .A2(n617), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U981 ( .A(KEYINPUT45), .B(n878), .Z(n879) );
  NOR2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n884) );
  XOR2_X1 U983 ( .A(n946), .B(n881), .Z(n882) );
  XNOR2_X1 U984 ( .A(n882), .B(G162), .ZN(n883) );
  XOR2_X1 U985 ( .A(n884), .B(n883), .Z(n896) );
  NAND2_X1 U986 ( .A1(G115), .A2(n616), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G127), .A2(n885), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n888), .B(KEYINPUT47), .ZN(n891) );
  NAND2_X1 U990 ( .A1(G103), .A2(n889), .ZN(n890) );
  NAND2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n894) );
  NAND2_X1 U992 ( .A1(n617), .A2(G139), .ZN(n892) );
  XOR2_X1 U993 ( .A(KEYINPUT112), .B(n892), .Z(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n938) );
  XNOR2_X1 U995 ( .A(G160), .B(n938), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U997 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n898) );
  XNOR2_X1 U998 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U1000 ( .A(n900), .B(n899), .Z(n903) );
  XNOR2_X1 U1001 ( .A(G164), .B(n901), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n906), .ZN(G395) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(G397), .A2(n908), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n913), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(KEYINPUT115), .B(n909), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(G395), .A2(n910), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n913), .ZN(G319) );
  INV_X1 U1014 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1015 ( .A(G16), .B(KEYINPUT56), .Z(n937) );
  XOR2_X1 U1016 ( .A(G168), .B(G1966), .Z(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1018 ( .A(KEYINPUT57), .B(n916), .Z(n932) );
  XNOR2_X1 U1019 ( .A(n917), .B(G1348), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(G1971), .A2(G303), .ZN(n918) );
  NAND2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(G1956), .B(G299), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(G1341), .B(n924), .ZN(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(G1961), .B(G301), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1032 ( .A(KEYINPUT125), .B(n935), .Z(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n967) );
  XOR2_X1 U1034 ( .A(G2072), .B(n938), .Z(n940) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n941), .Z(n961) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n945) );
  XOR2_X1 U1039 ( .A(G160), .B(G2084), .Z(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n952) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(KEYINPUT117), .B(n948), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n958) );
  XOR2_X1 U1045 ( .A(G2090), .B(G162), .Z(n953) );
  NOR2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(n955), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(KEYINPUT51), .B(n956), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(KEYINPUT119), .B(n959), .ZN(n960) );
  NOR2_X1 U1051 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1052 ( .A(KEYINPUT52), .B(n962), .Z(n963) );
  NOR2_X1 U1053 ( .A1(KEYINPUT55), .A2(n963), .ZN(n965) );
  INV_X1 U1054 ( .A(G29), .ZN(n964) );
  NOR2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1056 ( .A1(n967), .A2(n966), .ZN(n994) );
  XOR2_X1 U1057 ( .A(G29), .B(KEYINPUT124), .Z(n992) );
  XNOR2_X1 U1058 ( .A(G2090), .B(G35), .ZN(n984) );
  XNOR2_X1 U1059 ( .A(G25), .B(n968), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n969), .A2(G28), .ZN(n981) );
  XNOR2_X1 U1061 ( .A(G32), .B(n970), .ZN(n974) );
  XNOR2_X1 U1062 ( .A(G2067), .B(G26), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(G33), .B(G2072), .ZN(n971) );
  NOR2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n978) );
  XNOR2_X1 U1066 ( .A(G27), .B(n975), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(KEYINPUT120), .B(n976), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(n979), .B(KEYINPUT121), .ZN(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(KEYINPUT53), .B(n982), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n988) );
  XOR2_X1 U1073 ( .A(G34), .B(KEYINPUT122), .Z(n986) );
  XNOR2_X1 U1074 ( .A(G2084), .B(KEYINPUT54), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(n986), .B(n985), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1077 ( .A(n989), .B(KEYINPUT123), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(n990), .B(KEYINPUT55), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n1021) );
  XOR2_X1 U1081 ( .A(G1966), .B(G21), .Z(n1005) );
  XOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .Z(n995) );
  XNOR2_X1 U1083 ( .A(G4), .B(n995), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(G20), .B(G1956), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(G1981), .B(G6), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G1341), .B(G19), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1090 ( .A(KEYINPUT126), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1091 ( .A(n1003), .B(KEYINPUT60), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(KEYINPUT127), .B(n1006), .ZN(n1008) );
  XOR2_X1 U1094 ( .A(G1961), .B(G5), .Z(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1015) );
  XNOR2_X1 U1096 ( .A(G1976), .B(G23), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G1971), .B(G22), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(G1986), .B(G24), .Z(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1016), .ZN(n1018) );
  INV_X1 U1104 ( .A(G16), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(G11), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(n1022), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

