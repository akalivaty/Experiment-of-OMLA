//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(G134), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G137), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(G137), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT64), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n188), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G134), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT11), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n190), .A2(KEYINPUT64), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n194), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n192), .B2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n193), .A2(G134), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n194), .B2(new_n196), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n195), .A2(KEYINPUT11), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n189), .B1(new_n191), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n207), .A2(KEYINPUT0), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n213), .A3(G128), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n207), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n209), .B1(KEYINPUT0), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n206), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n200), .B2(new_n189), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(G143), .B2(new_n210), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n208), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT1), .B1(new_n212), .B2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n207), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n219), .B(new_n205), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n218), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT66), .B1(new_n230), .B2(G116), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(G119), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n231), .A2(new_n234), .B1(G116), .B2(new_n230), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT2), .B(G113), .Z(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n229), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n235), .A2(new_n236), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n235), .A2(new_n236), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n218), .A2(new_n228), .A3(new_n241), .A4(KEYINPUT68), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n205), .A2(new_n219), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n211), .A2(new_n213), .ZN(new_n245));
  OAI21_X1  g059(.A(G128), .B1(new_n224), .B2(KEYINPUT65), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n222), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n227), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n244), .A2(new_n250), .B1(new_n206), .B2(new_n217), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT68), .B1(new_n251), .B2(new_n241), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT28), .B1(new_n243), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n218), .A2(new_n228), .A3(new_n241), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(G237), .A2(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G210), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(KEYINPUT27), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n253), .A2(new_n256), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n218), .A2(new_n228), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n267), .B1(new_n218), .B2(new_n228), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n237), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n270), .A2(new_n254), .A3(new_n262), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n241), .B1(new_n218), .B2(new_n228), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n255), .B2(new_n254), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n218), .A2(new_n228), .A3(new_n241), .A4(KEYINPUT28), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n262), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n263), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n253), .A2(new_n278), .A3(new_n256), .A4(new_n264), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n266), .A2(new_n276), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G472), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n254), .A2(new_n261), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n270), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n270), .A2(new_n285), .A3(KEYINPUT67), .A4(new_n283), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n270), .A2(new_n285), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n256), .A2(new_n274), .A3(new_n238), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n291), .A2(KEYINPUT31), .B1(new_n262), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n282), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n295), .ZN(new_n297));
  AOI211_X1 g111(.A(KEYINPUT32), .B(new_n297), .C1(new_n290), .C2(new_n293), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n281), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT70), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT71), .B(G217), .Z(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(G234), .B2(new_n277), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT73), .B(G125), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT16), .ZN(new_n304));
  INV_X1    g118(.A(G140), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G125), .A2(G140), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(new_n303), .B2(G140), .ZN(new_n308));
  OAI211_X1 g122(.A(G146), .B(new_n306), .C1(new_n308), .C2(new_n304), .ZN(new_n309));
  XOR2_X1   g123(.A(G125), .B(G140), .Z(new_n310));
  OR2_X1    g124(.A1(new_n310), .A2(G146), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n230), .B2(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n230), .A2(G128), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(KEYINPUT23), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT23), .B1(new_n208), .B2(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n208), .A2(G119), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n312), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G110), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(new_n317), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT24), .B(G110), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n320), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n321), .B1(new_n320), .B2(new_n324), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n309), .B(new_n311), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  AND2_X1   g141(.A1(KEYINPUT73), .A2(G125), .ZN(new_n328));
  NOR2_X1   g142(.A1(KEYINPUT73), .A2(G125), .ZN(new_n329));
  OAI21_X1  g143(.A(G140), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n307), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n304), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n328), .A2(new_n329), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n333), .A2(KEYINPUT16), .A3(G140), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n210), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n309), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n322), .A2(new_n323), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n315), .A2(new_n318), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(G110), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G953), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(G221), .A3(G234), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT75), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT22), .B(G137), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n327), .A2(new_n340), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n345), .B1(new_n327), .B2(new_n340), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT25), .B1(new_n348), .B2(new_n277), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n350));
  NOR4_X1   g164(.A1(new_n346), .A2(new_n347), .A3(new_n350), .A4(G902), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n302), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n277), .B1(new_n301), .B2(G234), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT77), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n348), .A2(new_n356), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT76), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT70), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n281), .B(new_n362), .C1(new_n296), .C2(new_n298), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n300), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(G214), .B1(G237), .B2(G902), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(KEYINPUT88), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n250), .A2(new_n333), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n217), .A2(new_n303), .ZN(new_n368));
  INV_X1    g182(.A(G224), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G953), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT7), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n367), .B(new_n368), .C1(KEYINPUT90), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(KEYINPUT90), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n373), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(G107), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(KEYINPUT3), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(G107), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT81), .ZN(new_n386));
  INV_X1    g200(.A(G107), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n377), .B(G101), .C1(new_n383), .C2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n239), .B2(new_n240), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n385), .A2(KEYINPUT81), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n386), .B1(new_n393), .B2(new_n388), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT82), .B(G101), .Z(new_n395));
  NAND2_X1  g209(.A1(new_n379), .A2(new_n381), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n384), .A4(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n387), .A2(G104), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(new_n379), .B2(new_n381), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n401), .A2(new_n394), .A3(KEYINPUT83), .A4(new_n395), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n394), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n377), .B1(new_n404), .B2(G101), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT84), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n380), .B2(G107), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(new_n400), .ZN(new_n410));
  OAI21_X1  g224(.A(G101), .B1(new_n388), .B2(new_n408), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G101), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n381), .B2(KEYINPUT84), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n388), .A2(new_n384), .A3(new_n408), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(KEYINPUT85), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n399), .B2(new_n402), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n230), .A2(G116), .ZN(new_n419));
  OAI21_X1  g233(.A(G113), .B1(new_n419), .B2(KEYINPUT5), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n420), .B1(new_n235), .B2(KEYINPUT5), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n239), .A2(new_n421), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n392), .A2(new_n406), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G122), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n424), .B(KEYINPUT8), .Z(new_n425));
  NOR3_X1   g239(.A1(new_n410), .A2(new_n411), .A3(new_n407), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT85), .B1(new_n414), .B2(new_n415), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n403), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n425), .B1(new_n429), .B2(new_n422), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n231), .A2(new_n234), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT5), .A3(new_n419), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n420), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n235), .A2(KEYINPUT89), .A3(KEYINPUT5), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n418), .B1(new_n436), .B2(new_n239), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n423), .A2(new_n424), .B1(new_n430), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(G902), .B1(new_n376), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n424), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n403), .A2(new_n422), .A3(new_n428), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n391), .B1(new_n403), .B2(new_n405), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n383), .A2(new_n389), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT4), .B1(new_n445), .B2(new_n413), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n399), .B2(new_n402), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n441), .B(new_n424), .C1(new_n447), .C2(new_n391), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(KEYINPUT6), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(new_n440), .C1(new_n442), .C2(new_n443), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n367), .A2(new_n368), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n371), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G210), .B1(G237), .B2(G902), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n439), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n439), .B2(new_n454), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n366), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n308), .A2(G146), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n311), .ZN(new_n460));
  INV_X1    g274(.A(G237), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n341), .A3(G214), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n212), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n257), .A2(G143), .A3(G214), .ZN(new_n464));
  NAND2_X1  g278(.A1(KEYINPUT18), .A2(G131), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n465), .A2(KEYINPUT92), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(KEYINPUT92), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n463), .A2(new_n464), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n463), .A2(new_n464), .ZN(new_n470));
  INV_X1    g284(.A(new_n465), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI211_X1 g286(.A(KEYINPUT91), .B(new_n465), .C1(new_n463), .C2(new_n464), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n460), .B(new_n468), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n464), .ZN(new_n475));
  AOI21_X1  g289(.A(G143), .B1(new_n257), .B2(G214), .ZN(new_n476));
  OAI21_X1  g290(.A(G131), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT17), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n463), .A2(new_n204), .A3(new_n464), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n470), .A2(KEYINPUT17), .A3(G131), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n335), .A2(new_n480), .A3(new_n309), .A4(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(G113), .B(G122), .Z(new_n483));
  XOR2_X1   g297(.A(KEYINPUT93), .B(G104), .Z(new_n484));
  XOR2_X1   g298(.A(new_n483), .B(new_n484), .Z(new_n485));
  NAND3_X1  g299(.A1(new_n474), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT94), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n474), .A2(new_n482), .A3(KEYINPUT94), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n474), .A2(new_n482), .ZN(new_n491));
  INV_X1    g305(.A(new_n485), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT95), .A3(new_n277), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n488), .A2(new_n489), .B1(new_n492), .B2(new_n491), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(G902), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n498), .A3(G475), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n310), .A2(KEYINPUT19), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(KEYINPUT19), .B2(new_n308), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n210), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n477), .A2(new_n479), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n309), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n474), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n492), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n490), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT20), .ZN(new_n508));
  INV_X1    g322(.A(G475), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n277), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n488), .A2(new_n489), .B1(new_n505), .B2(new_n492), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n277), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT20), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT96), .ZN(new_n515));
  INV_X1    g329(.A(G122), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G116), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n233), .A2(G122), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G107), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n518), .A3(new_n387), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT13), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n208), .B2(G143), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n208), .A2(G143), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n212), .A2(G128), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(new_n523), .ZN(new_n528));
  OAI21_X1  g342(.A(G134), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n525), .A3(new_n187), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n522), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n525), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G134), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n530), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT14), .B1(new_n516), .B2(G116), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT14), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n233), .A3(G122), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n537), .A3(new_n517), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G107), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n534), .A2(new_n521), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n515), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT9), .B(G234), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n301), .A2(G953), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n531), .A2(new_n540), .A3(new_n515), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n544), .ZN(new_n547));
  INV_X1    g361(.A(new_n545), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n547), .B1(new_n548), .B2(new_n541), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n549), .A3(new_n277), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n546), .A2(new_n549), .A3(KEYINPUT97), .A4(new_n277), .ZN(new_n553));
  INV_X1    g367(.A(G478), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(KEYINPUT15), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n550), .B(new_n551), .C1(KEYINPUT15), .C2(new_n554), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n341), .A2(G952), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(G234), .B2(G237), .ZN(new_n560));
  AOI211_X1 g374(.A(new_n277), .B(new_n341), .C1(G234), .C2(G237), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT21), .B(G898), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n499), .A2(new_n514), .A3(new_n558), .A4(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n458), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n418), .A2(new_n250), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n245), .B1(new_n221), .B2(new_n208), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n249), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT83), .B1(new_n445), .B2(new_n395), .ZN(new_n571));
  INV_X1    g385(.A(new_n402), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n428), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT86), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n418), .A2(KEYINPUT86), .A3(new_n570), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n568), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n206), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n567), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n429), .A2(new_n249), .A3(new_n248), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT86), .B1(new_n418), .B2(new_n570), .ZN(new_n581));
  AND4_X1   g395(.A1(KEYINPUT86), .A2(new_n403), .A3(new_n428), .A4(new_n570), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT12), .A3(new_n206), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n341), .A2(G227), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT80), .ZN(new_n587));
  XNOR2_X1  g401(.A(G110), .B(G140), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n589), .B(new_n590), .Z(new_n591));
  NAND2_X1  g405(.A1(new_n217), .A2(new_n390), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n250), .A2(KEYINPUT10), .ZN(new_n593));
  OAI22_X1  g407(.A1(new_n447), .A2(new_n592), .B1(new_n429), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n575), .A2(new_n576), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT87), .B(KEYINPUT10), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n591), .B1(new_n597), .B2(new_n578), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n585), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n596), .B1(new_n581), .B2(new_n582), .ZN(new_n600));
  INV_X1    g414(.A(new_n594), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n578), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n596), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n575), .B2(new_n576), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n604), .A2(new_n206), .A3(new_n594), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n591), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G469), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n277), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n598), .B1(new_n578), .B2(new_n597), .ZN(new_n610));
  INV_X1    g424(.A(new_n591), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n605), .B1(new_n584), .B2(new_n579), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n610), .B(G469), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n608), .A2(new_n277), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G221), .B1(new_n543), .B2(G902), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n566), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n364), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n395), .ZN(G3));
  NAND2_X1  g434(.A1(new_n616), .A2(new_n617), .ZN(new_n621));
  AOI21_X1  g435(.A(G902), .B1(new_n290), .B2(new_n293), .ZN(new_n622));
  INV_X1    g436(.A(G472), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT98), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n292), .A2(new_n262), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n229), .A2(KEYINPUT30), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n218), .A2(new_n228), .A3(new_n267), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n284), .B1(new_n629), .B2(new_n237), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n626), .B1(new_n630), .B2(new_n283), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n288), .B2(new_n289), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n625), .B(G472), .C1(new_n632), .C2(G902), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n297), .B1(new_n290), .B2(new_n293), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n360), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n624), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n365), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n439), .A2(new_n454), .ZN(new_n638));
  INV_X1    g452(.A(new_n455), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n439), .A2(new_n454), .A3(new_n455), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n546), .A2(new_n549), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n554), .A2(G902), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n550), .A2(new_n554), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n499), .A2(new_n514), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n642), .A2(new_n649), .A3(new_n564), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n621), .A2(new_n636), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT34), .B(G104), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  AND3_X1   g467(.A1(new_n510), .A2(KEYINPUT99), .A3(new_n513), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT99), .B1(new_n510), .B2(new_n513), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n558), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n657), .A2(new_n499), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n656), .A2(new_n658), .A3(new_n642), .A4(new_n564), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n621), .A2(new_n659), .A3(new_n636), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n387), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT100), .B(KEYINPUT35), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  INV_X1    g477(.A(new_n634), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n327), .A2(new_n340), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT36), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n345), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n665), .B(new_n667), .Z(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n355), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n352), .A2(new_n670), .ZN(new_n671));
  AND4_X1   g485(.A1(new_n664), .A2(new_n624), .A3(new_n633), .A4(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n617), .ZN(new_n673));
  AOI21_X1  g487(.A(G902), .B1(new_n599), .B2(new_n606), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n614), .B1(new_n674), .B2(new_n608), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n673), .B1(new_n675), .B2(new_n613), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n672), .A2(new_n676), .A3(new_n566), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  INV_X1    g493(.A(new_n642), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n352), .A2(new_n670), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n300), .A2(new_n363), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n560), .B1(new_n561), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n656), .A2(new_n658), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n676), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XNOR2_X1  g504(.A(new_n685), .B(KEYINPUT39), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n621), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n640), .A2(new_n641), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n681), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT32), .B1(new_n632), .B2(new_n297), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n634), .A2(new_n282), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n254), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n629), .B2(new_n237), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n703), .A2(new_n262), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n277), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n243), .A2(new_n252), .A3(new_n261), .ZN(new_n706));
  OAI21_X1  g520(.A(G472), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n499), .A2(new_n514), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n365), .A3(new_n657), .ZN(new_n710));
  OR3_X1    g524(.A1(new_n698), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n694), .A2(new_n695), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n212), .ZN(G45));
  NAND2_X1  g527(.A1(new_n649), .A2(new_n686), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n676), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n683), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT101), .B(G146), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G48));
  NAND2_X1  g533(.A1(new_n607), .A2(new_n277), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G469), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n617), .A3(new_n609), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n650), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n361), .A3(new_n300), .A4(new_n363), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT41), .B(G113), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT102), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n724), .B(new_n726), .ZN(G15));
  NOR2_X1   g541(.A1(new_n722), .A2(new_n659), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n361), .A3(new_n300), .A4(new_n363), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  NOR2_X1   g544(.A1(new_n722), .A2(new_n680), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n565), .A2(new_n681), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n300), .A3(new_n363), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  AND3_X1   g548(.A1(new_n721), .A2(new_n617), .A3(new_n609), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n622), .A2(new_n623), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n253), .A2(new_n256), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT103), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n253), .A2(new_n739), .A3(new_n256), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n262), .A3(new_n740), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n288), .A2(new_n289), .B1(KEYINPUT31), .B2(new_n291), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n297), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n736), .A2(new_n743), .A3(new_n360), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n696), .A2(new_n709), .A3(new_n365), .A4(new_n657), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n563), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n735), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NOR3_X1   g562(.A1(new_n736), .A2(new_n743), .A3(new_n681), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n735), .A2(new_n642), .A3(new_n715), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  NAND2_X1  g565(.A1(new_n299), .A2(new_n361), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n640), .A2(new_n617), .A3(new_n641), .A4(new_n365), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n616), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n752), .A2(new_n755), .A3(new_n756), .A4(new_n714), .ZN(new_n757));
  AOI211_X1 g571(.A(new_n360), .B(new_n753), .C1(new_n675), .C2(new_n613), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n300), .A3(new_n363), .A4(new_n715), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT42), .B1(new_n759), .B2(KEYINPUT104), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n362), .B1(new_n701), .B2(new_n281), .ZN(new_n761));
  INV_X1    g575(.A(new_n363), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT104), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n715), .A4(new_n758), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n757), .B1(new_n760), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n204), .ZN(G33));
  AND3_X1   g581(.A1(new_n758), .A2(new_n300), .A3(new_n363), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n687), .B(KEYINPUT105), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  NAND2_X1  g585(.A1(new_n647), .A2(new_n648), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n514), .A3(new_n499), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT43), .Z(new_n774));
  NAND3_X1  g588(.A1(new_n624), .A2(new_n633), .A3(new_n664), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(new_n671), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n640), .A2(new_n641), .A3(new_n365), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n608), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n615), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT46), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n609), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n617), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(new_n691), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(KEYINPUT106), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(KEYINPUT106), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n781), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  OR3_X1    g610(.A1(new_n714), .A2(new_n361), .A3(new_n780), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n791), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n791), .A2(new_n798), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n763), .B(new_n797), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n305), .ZN(G42));
  NAND2_X1  g616(.A1(new_n721), .A2(new_n609), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(KEYINPUT49), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT107), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n361), .A2(new_n617), .A3(new_n366), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n697), .A2(new_n773), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n803), .A2(KEYINPUT49), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n805), .A2(new_n708), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n724), .A2(new_n729), .A3(new_n733), .A4(new_n747), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n759), .A2(KEYINPUT104), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n765), .A3(new_n756), .ZN(new_n812));
  INV_X1    g626(.A(new_n757), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n681), .A2(new_n685), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT108), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n558), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n556), .A2(KEYINPUT108), .A3(new_n557), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n815), .A2(new_n499), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(new_n300), .A3(new_n363), .A4(new_n656), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n749), .A2(new_n715), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n770), .B1(new_n823), .B2(new_n755), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n624), .A2(new_n633), .A3(new_n635), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n696), .A2(new_n366), .A3(new_n564), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n817), .A2(new_n514), .A3(new_n499), .A4(new_n818), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(new_n676), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT109), .B1(new_n677), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n649), .A2(new_n696), .A3(new_n366), .A4(new_n564), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n826), .A2(new_n833), .A3(new_n676), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n364), .B2(new_n618), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n677), .A2(KEYINPUT109), .A3(new_n830), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT110), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n621), .A2(new_n636), .A3(new_n832), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n300), .A2(new_n361), .A3(new_n363), .ZN(new_n840));
  INV_X1    g654(.A(new_n618), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT109), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n826), .A2(new_n676), .A3(new_n829), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n624), .A2(new_n633), .A3(new_n664), .A4(new_n671), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n618), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n843), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  AND4_X1   g661(.A1(KEYINPUT110), .A2(new_n842), .A3(new_n847), .A4(new_n837), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n814), .B(new_n825), .C1(new_n838), .C2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n750), .B1(new_n683), .B2(new_n688), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n717), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n745), .B1(new_n701), .B2(new_n707), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n671), .A2(new_n685), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n616), .A2(KEYINPUT112), .A3(new_n617), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT112), .B1(new_n676), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n616), .A2(new_n617), .A3(new_n854), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT112), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT113), .A3(new_n855), .A4(new_n853), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n851), .A2(new_n863), .A3(KEYINPUT52), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(new_n851), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT53), .B1(new_n849), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n842), .A2(new_n847), .A3(new_n837), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT110), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n836), .A2(KEYINPUT110), .A3(new_n837), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n824), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n858), .A2(new_n862), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n621), .A2(new_n714), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n763), .A2(new_n875), .A3(new_n682), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n689), .A2(new_n876), .A3(new_n750), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n873), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n717), .B1(new_n850), .B2(KEYINPUT111), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT111), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n750), .B(new_n880), .C1(new_n683), .C2(new_n688), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(KEYINPUT52), .A3(new_n863), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n872), .A2(new_n883), .A3(new_n884), .A4(new_n814), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n867), .A2(KEYINPUT54), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n884), .B1(new_n849), .B2(new_n866), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n825), .B1(new_n838), .B2(new_n848), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT114), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT114), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n872), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n812), .A2(new_n813), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n895));
  INV_X1    g709(.A(new_n810), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT115), .B1(new_n766), .B2(new_n810), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n883), .A2(KEYINPUT53), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n887), .B(new_n888), .C1(new_n893), .C2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT116), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n886), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n774), .A2(new_n560), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n722), .A2(new_n780), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n752), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT48), .Z(new_n907));
  XOR2_X1   g721(.A(new_n559), .B(KEYINPUT117), .Z(new_n908));
  NAND4_X1  g722(.A1(new_n904), .A2(new_n361), .A3(new_n560), .A4(new_n708), .ZN(new_n909));
  INV_X1    g723(.A(new_n649), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n903), .A2(new_n744), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n913), .B2(new_n731), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n909), .A2(new_n709), .A3(new_n772), .ZN(new_n915));
  INV_X1    g729(.A(new_n749), .ZN(new_n916));
  INV_X1    g730(.A(new_n744), .ZN(new_n917));
  NOR4_X1   g731(.A1(new_n917), .A2(new_n697), .A3(new_n722), .A4(new_n365), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n918), .A2(new_n903), .A3(KEYINPUT50), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT50), .B1(new_n918), .B2(new_n903), .ZN(new_n920));
  OAI221_X1 g734(.A(new_n915), .B1(new_n916), .B2(new_n905), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n799), .B(new_n800), .C1(new_n617), .C2(new_n803), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n912), .A2(new_n780), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n907), .B(new_n914), .C1(new_n924), .C2(KEYINPUT51), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(KEYINPUT51), .B2(new_n924), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n897), .A2(new_n898), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n884), .B1(new_n878), .B2(new_n882), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n890), .A2(new_n927), .A3(new_n892), .A4(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n929), .A2(KEYINPUT116), .A3(new_n887), .A4(new_n888), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n902), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n931), .A2(new_n932), .B1(G952), .B2(G953), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n809), .B1(new_n933), .B2(new_n934), .ZN(G75));
  NOR2_X1   g749(.A1(new_n341), .A2(G952), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n929), .A2(new_n888), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(G902), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT56), .B1(new_n940), .B2(G210), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n449), .A2(new_n451), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n453), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n937), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT56), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n944), .B(KEYINPUT119), .ZN(new_n947));
  INV_X1    g761(.A(G210), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n946), .B(new_n947), .C1(new_n939), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT120), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n949), .A2(KEYINPUT120), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(G51));
  NAND2_X1  g766(.A1(new_n870), .A2(new_n871), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n891), .B1(new_n953), .B2(new_n825), .ZN(new_n954));
  AOI211_X1 g768(.A(KEYINPUT114), .B(new_n824), .C1(new_n870), .C2(new_n871), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n899), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n888), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT54), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(KEYINPUT122), .A3(new_n900), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n938), .A2(new_n960), .A3(KEYINPUT54), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n614), .B(KEYINPUT121), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT57), .Z(new_n963));
  NAND3_X1  g777(.A1(new_n959), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n607), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n939), .A2(new_n785), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n936), .B1(new_n965), .B2(new_n966), .ZN(G54));
  NAND3_X1  g781(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n968), .A2(new_n511), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n511), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n936), .ZN(G60));
  INV_X1    g785(.A(new_n645), .ZN(new_n972));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT59), .Z(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n959), .A2(new_n961), .A3(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n976), .A2(new_n937), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n900), .A2(new_n901), .ZN(new_n978));
  INV_X1    g792(.A(new_n886), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n930), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n974), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT123), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n982), .A2(new_n983), .A3(new_n972), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n974), .B1(new_n902), .B2(new_n930), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT123), .B1(new_n985), .B2(new_n645), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n977), .A2(new_n984), .A3(new_n986), .ZN(G63));
  NOR2_X1   g801(.A1(new_n956), .A2(new_n957), .ZN(new_n988));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT124), .Z(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT60), .ZN(new_n991));
  OR3_X1    g805(.A1(new_n988), .A2(new_n668), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n357), .A2(new_n358), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n988), .B2(new_n991), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n992), .A2(new_n937), .A3(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(G66));
  OAI21_X1  g811(.A(G953), .B1(new_n562), .B2(new_n369), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT125), .Z(new_n999));
  NAND2_X1  g813(.A1(new_n953), .A2(new_n896), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n999), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n942), .B1(G898), .B2(new_n341), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(G69));
  XNOR2_X1  g818(.A(new_n629), .B(new_n501), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(G900), .B2(G953), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n879), .A2(new_n881), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n801), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n752), .A2(new_n745), .ZN(new_n1010));
  OAI22_X1  g824(.A1(new_n793), .A2(new_n794), .B1(new_n781), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1009), .A2(new_n894), .A3(new_n770), .A4(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1007), .B1(new_n1012), .B2(G953), .ZN(new_n1013));
  AOI211_X1 g827(.A(new_n780), .B(new_n693), .C1(new_n910), .C2(new_n828), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n801), .B1(new_n840), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g829(.A1(new_n1008), .A2(new_n712), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n1016), .A2(KEYINPUT62), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(KEYINPUT62), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1015), .A2(new_n795), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n1019), .A2(new_n341), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1013), .B1(new_n1020), .B2(new_n1005), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n341), .B1(G227), .B2(G900), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1021), .B(new_n1022), .ZN(G72));
  XOR2_X1   g837(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1024));
  NOR2_X1   g838(.A1(new_n623), .A2(new_n277), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(new_n1012), .B2(new_n1000), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n271), .B(KEYINPUT127), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n936), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n867), .A2(new_n885), .ZN(new_n1030));
  INV_X1    g844(.A(new_n271), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n704), .A2(new_n1031), .A3(new_n1026), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1029), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n704), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1026), .B1(new_n1019), .B2(new_n1000), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(G57));
endmodule


