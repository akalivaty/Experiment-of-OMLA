//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  XOR2_X1   g000(.A(G183gat), .B(G211gat), .Z(new_n202));
  XOR2_X1   g001(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n203));
  OAI21_X1  g002(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G71gat), .B(G78gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT95), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G231gat), .A2(G233gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G127gat), .B(G155gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n215), .A2(new_n216), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n203), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n215), .A2(new_n216), .ZN(new_n221));
  INV_X1    g020(.A(new_n203), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OR3_X1    g023(.A1(new_n224), .A2(KEYINPUT90), .A3(G1gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT90), .B1(new_n224), .B2(G1gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n228), .B(KEYINPUT91), .C1(G1gat), .C2(new_n226), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n229), .B(G8gat), .Z(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n211), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(KEYINPUT21), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n220), .A2(new_n223), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n220), .B2(new_n223), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n202), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n223), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n233), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n223), .A3(new_n234), .ZN(new_n240));
  INV_X1    g039(.A(new_n202), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G190gat), .B(G218gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(G99gat), .A2(G106gat), .ZN(new_n245));
  INV_X1    g044(.A(G85gat), .ZN(new_n246));
  INV_X1    g045(.A(G92gat), .ZN(new_n247));
  AOI22_X1  g046(.A1(KEYINPUT8), .A2(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n246), .B2(new_n247), .ZN(new_n250));
  NAND4_X1  g049(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n248), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G99gat), .B(G106gat), .Z(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  INV_X1    g053(.A(KEYINPUT17), .ZN(new_n255));
  NOR3_X1   g054(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n257), .A2(new_n258), .B1(G29gat), .B2(G36gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT87), .B(G50gat), .ZN(new_n260));
  INV_X1    g059(.A(G43gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G50gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G43gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT15), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT88), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n261), .A2(G50gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(new_n269), .A3(KEYINPUT15), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n267), .A2(KEYINPUT88), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n259), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n259), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n270), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n273), .A2(KEYINPUT89), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT89), .B1(new_n273), .B2(new_n275), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n255), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n275), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(new_n255), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n254), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT89), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n273), .A2(KEYINPUT89), .A3(new_n275), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n254), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n283), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n244), .B1(new_n282), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT99), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT99), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n292), .B(new_n244), .C1(new_n282), .C2(new_n289), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT96), .ZN(new_n295));
  XNOR2_X1  g094(.A(G134gat), .B(G162gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT17), .B1(new_n285), .B2(new_n286), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n288), .B1(new_n298), .B2(new_n280), .ZN(new_n299));
  INV_X1    g098(.A(new_n283), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n276), .A2(new_n277), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n254), .ZN(new_n302));
  INV_X1    g101(.A(new_n244), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n291), .A2(new_n293), .A3(new_n297), .A4(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n297), .B(KEYINPUT97), .Z(new_n306));
  AOI21_X1  g105(.A(new_n306), .B1(new_n290), .B2(new_n304), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G120gat), .B(G148gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(G176gat), .B(G204gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n232), .A2(KEYINPUT10), .A3(new_n254), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n211), .A2(new_n288), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n288), .A2(new_n209), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n316), .B2(KEYINPUT10), .ZN(new_n317));
  NAND2_X1  g116(.A1(G230gat), .A2(G233gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT100), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n318), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n312), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n317), .A2(new_n318), .ZN(new_n325));
  INV_X1    g124(.A(new_n312), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n243), .A2(new_n309), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT93), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT34), .ZN(new_n332));
  INV_X1    g131(.A(G169gat), .ZN(new_n333));
  INV_X1    g132(.A(G176gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT23), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(G169gat), .B2(G176gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  AND4_X1   g137(.A1(KEYINPUT25), .A2(new_n335), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT65), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT65), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n349));
  AND3_X1   g148(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n350), .B1(new_n341), .B2(new_n340), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NOR3_X1   g153(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT27), .B(G183gat), .ZN(new_n360));
  INV_X1    g159(.A(G190gat), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT28), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G183gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT27), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G183gat), .ZN(new_n366));
  AND4_X1   g165(.A1(KEYINPUT28), .A2(new_n364), .A3(new_n366), .A4(new_n361), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n341), .B(new_n359), .C1(new_n362), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n354), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G120gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G113gat), .ZN(new_n371));
  INV_X1    g170(.A(G113gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G120gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT66), .ZN(new_n377));
  INV_X1    g176(.A(G127gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G134gat), .ZN(new_n379));
  INV_X1    g178(.A(G134gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(G127gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(G127gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(G134gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT66), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n376), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT67), .B1(new_n379), .B2(new_n381), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT1), .B1(new_n371), .B2(new_n373), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT67), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(new_n384), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n369), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n386), .A2(new_n391), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n354), .A2(new_n394), .A3(new_n368), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n332), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT68), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n332), .A3(new_n397), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n398), .A2(new_n399), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G15gat), .B(G43gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n393), .A2(G227gat), .A3(G233gat), .A4(new_n395), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(KEYINPUT32), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n411), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n404), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n402), .A2(new_n403), .A3(new_n412), .A4(new_n413), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n417), .A2(KEYINPUT69), .A3(KEYINPUT36), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT36), .B1(new_n417), .B2(KEYINPUT69), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G197gat), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n421), .A2(G204gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(G204gat), .ZN(new_n423));
  INV_X1    g222(.A(G211gat), .ZN(new_n424));
  INV_X1    g223(.A(G218gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n422), .B(new_n423), .C1(new_n426), .C2(KEYINPUT22), .ZN(new_n427));
  XOR2_X1   g226(.A(G211gat), .B(G218gat), .Z(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT70), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n342), .A2(new_n343), .ZN(new_n432));
  AND2_X1   g231(.A1(G169gat), .A2(G176gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n333), .A2(new_n334), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n336), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n335), .A3(new_n435), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n436), .A2(new_n349), .B1(new_n347), .B2(new_n339), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n358), .A2(new_n357), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n341), .B1(new_n438), .B2(new_n355), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n360), .A2(new_n361), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT28), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n360), .A2(KEYINPUT28), .A3(new_n361), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n439), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n431), .B1(new_n437), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT29), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n354), .A2(KEYINPUT70), .A3(new_n368), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT71), .ZN(new_n449));
  NAND2_X1  g248(.A1(G226gat), .A2(G233gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n450), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n369), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n449), .B1(new_n448), .B2(new_n450), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n430), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n445), .A2(new_n447), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n452), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n369), .A2(new_n446), .A3(new_n450), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n430), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G8gat), .B(G36gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(G64gat), .B(G92gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n465), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n456), .A2(new_n461), .A3(KEYINPUT30), .A4(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n456), .A2(new_n461), .A3(new_n467), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n469), .A2(KEYINPUT72), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT72), .B1(new_n469), .B2(new_n470), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n466), .B(new_n468), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT0), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT77), .ZN(new_n476));
  XOR2_X1   g275(.A(G57gat), .B(G85gat), .Z(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT5), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT76), .ZN(new_n481));
  OR2_X1    g280(.A1(G155gat), .A2(G162gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(G155gat), .A2(G162gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(KEYINPUT74), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT74), .ZN(new_n485));
  AND2_X1   g284(.A1(G155gat), .A2(G162gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(G155gat), .A2(G162gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n483), .A2(KEYINPUT2), .ZN(new_n489));
  AND2_X1   g288(.A1(G141gat), .A2(G148gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(G141gat), .A2(G148gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n484), .A2(new_n488), .A3(new_n489), .A4(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(G141gat), .A2(G148gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(G141gat), .A2(G148gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n489), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT73), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n483), .B1(new_n487), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n486), .A2(KEYINPUT73), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n392), .A2(new_n481), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n493), .A2(new_n500), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT76), .B1(new_n394), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n394), .A2(new_n503), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G225gat), .A2(G233gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n480), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n502), .A2(new_n510), .A3(new_n504), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT3), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT75), .B1(new_n501), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n493), .A2(new_n500), .A3(new_n512), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n394), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT75), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n503), .A2(new_n516), .A3(KEYINPUT3), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n394), .A2(new_n503), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n508), .B1(new_n519), .B2(KEYINPUT4), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n511), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n509), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n502), .A2(new_n504), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT4), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n510), .B1(new_n394), .B2(new_n503), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n524), .A2(new_n518), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n479), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n479), .A3(new_n527), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT78), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT78), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n533), .A3(new_n530), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n528), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n536));
  AOI211_X1 g335(.A(new_n530), .B(new_n479), .C1(new_n522), .C2(new_n527), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(new_n535), .B2(KEYINPUT79), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n473), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G78gat), .B(G106gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(new_n263), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT80), .B(KEYINPUT31), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(G22gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(G228gat), .A2(G233gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n429), .A2(new_n446), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n501), .B1(new_n546), .B2(new_n512), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n514), .A2(new_n446), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT82), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n549), .B2(new_n430), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n546), .B(KEYINPUT81), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(KEYINPUT3), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(new_n501), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n430), .A2(new_n548), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n545), .ZN(new_n555));
  OAI221_X1 g354(.A(new_n544), .B1(new_n545), .B2(new_n550), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n544), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n551), .A2(KEYINPUT3), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n555), .B1(new_n558), .B2(new_n503), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n550), .A2(new_n545), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n420), .B1(new_n539), .B2(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n564), .A2(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(KEYINPUT83), .ZN(new_n566));
  INV_X1    g365(.A(new_n531), .ZN(new_n567));
  INV_X1    g366(.A(new_n528), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n537), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n455), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(new_n451), .A3(new_n453), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n429), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n458), .A2(new_n459), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n430), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT38), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n465), .B1(new_n462), .B2(KEYINPUT37), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n569), .B(new_n469), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n460), .B1(new_n571), .B2(new_n430), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n467), .B1(new_n581), .B2(new_n573), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n462), .A2(KEYINPUT37), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n577), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n563), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n506), .A2(new_n508), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT39), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n518), .A2(new_n525), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n510), .B1(new_n502), .B2(new_n504), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n508), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n478), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n587), .B(new_n508), .C1(new_n589), .C2(new_n590), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(KEYINPUT40), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT84), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n592), .A2(new_n596), .A3(KEYINPUT40), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT40), .B1(new_n592), .B2(new_n593), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(new_n528), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n473), .A2(KEYINPUT85), .A3(new_n598), .A4(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT85), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n468), .B1(new_n581), .B2(new_n467), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n469), .A2(new_n470), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT72), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n469), .A2(KEYINPUT72), .A3(new_n470), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n598), .A2(new_n600), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n585), .B1(new_n601), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n565), .A2(new_n566), .A3(new_n612), .ZN(new_n613));
  OR4_X1    g412(.A1(KEYINPUT35), .A2(new_n417), .A3(new_n562), .A4(new_n569), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n614), .A2(new_n473), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n417), .A2(new_n562), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n529), .A2(new_n533), .A3(new_n530), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n533), .B1(new_n529), .B2(new_n530), .ZN(new_n619));
  OAI211_X1 g418(.A(KEYINPUT79), .B(new_n568), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n537), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n608), .B(new_n616), .C1(new_n617), .C2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT86), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT35), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n624), .B1(new_n623), .B2(KEYINPUT35), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n615), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n613), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n230), .B1(new_n298), .B2(new_n280), .ZN(new_n629));
  NAND2_X1  g428(.A1(G229gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n301), .A2(new_n231), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n629), .A2(KEYINPUT18), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n630), .B(KEYINPUT13), .Z(new_n633));
  NOR2_X1   g432(.A1(new_n301), .A2(new_n231), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n287), .A2(new_n230), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G113gat), .B(G141gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT11), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(new_n333), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G197gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n632), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT18), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n643), .A2(KEYINPUT92), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT92), .B1(new_n643), .B2(new_n644), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n644), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n632), .A3(new_n636), .ZN(new_n649));
  INV_X1    g448(.A(new_n641), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n331), .B1(new_n628), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n647), .A2(new_n651), .ZN(new_n655));
  AOI211_X1 g454(.A(KEYINPUT93), .B(new_n655), .C1(new_n613), .C2(new_n627), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n330), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n536), .A2(new_n538), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT101), .B(G1gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1324gat));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  NAND3_X1  g463(.A1(new_n658), .A2(new_n473), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n658), .A2(new_n473), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n668), .B2(G8gat), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n665), .B2(new_n669), .ZN(G1325gat));
  INV_X1    g469(.A(G15gat), .ZN(new_n671));
  INV_X1    g470(.A(new_n417), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n658), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n420), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n673), .B1(new_n676), .B2(new_n671), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n658), .A2(new_n562), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NOR3_X1   g479(.A1(new_n243), .A2(new_n309), .A3(new_n328), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n653), .B2(new_n656), .ZN(new_n682));
  OR3_X1    g481(.A1(new_n682), .A2(G29gat), .A3(new_n659), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n627), .A2(KEYINPUT102), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n615), .B(new_n686), .C1(new_n625), .C2(new_n626), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n564), .A2(new_n611), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n305), .A2(new_n308), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(KEYINPUT44), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n613), .B2(new_n627), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n243), .A2(new_n655), .A3(new_n328), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698), .B2(new_n659), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n699), .ZN(G1328gat));
  NOR2_X1   g499(.A1(new_n608), .A2(G36gat), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n681), .B(new_n701), .C1(new_n653), .C2(new_n656), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(KEYINPUT46), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n698), .A2(new_n608), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(G36gat), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n702), .B2(KEYINPUT46), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n702), .A2(new_n707), .A3(KEYINPUT46), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n705), .B(new_n706), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n708), .ZN(new_n711));
  OAI21_X1  g510(.A(G36gat), .B1(new_n698), .B2(new_n608), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(KEYINPUT46), .B2(new_n702), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT104), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(G1329gat));
  OAI21_X1  g514(.A(G43gat), .B1(new_n698), .B2(new_n420), .ZN(new_n716));
  OR2_X1    g515(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n672), .A2(new_n261), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n716), .B(new_n717), .C1(new_n682), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1330gat));
  XNOR2_X1  g520(.A(new_n682), .B(KEYINPUT106), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n563), .A2(new_n260), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT48), .ZN(new_n725));
  INV_X1    g524(.A(new_n260), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n698), .A2(new_n563), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n728));
  OR3_X1    g527(.A1(new_n698), .A2(KEYINPUT107), .A3(new_n563), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n722), .A2(new_n723), .B1(new_n260), .B2(new_n727), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n725), .A2(new_n730), .B1(new_n731), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g531(.A1(new_n243), .A2(new_n655), .A3(new_n309), .A4(new_n328), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n564), .A2(new_n611), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n627), .B2(KEYINPUT102), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n733), .B1(new_n735), .B2(new_n687), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n660), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT108), .B(G57gat), .Z(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1332gat));
  XNOR2_X1  g538(.A(new_n473), .B(KEYINPUT109), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n743), .B2(new_n742), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT110), .ZN(G1333gat));
  AOI21_X1  g546(.A(G71gat), .B1(new_n736), .B2(new_n672), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n674), .A2(G71gat), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n736), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n562), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT111), .B(G78gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n243), .A2(new_n652), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n693), .A2(new_n328), .A3(new_n696), .A4(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756), .B2(new_n659), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n614), .A2(new_n473), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n623), .A2(KEYINPUT35), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT86), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT35), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n688), .B1(new_n763), .B2(new_n686), .ZN(new_n764));
  INV_X1    g563(.A(new_n687), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n758), .B(new_n690), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n755), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n758), .B1(new_n689), .B2(new_n690), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(KEYINPUT113), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(new_n772));
  INV_X1    g571(.A(new_n755), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n309), .B1(new_n735), .B2(new_n687), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n758), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n691), .A2(KEYINPUT112), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n772), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n771), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n660), .A2(new_n246), .A3(new_n328), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n757), .B1(new_n780), .B2(new_n781), .ZN(G1336gat));
  AOI21_X1  g581(.A(KEYINPUT44), .B1(new_n689), .B2(new_n690), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n755), .A2(new_n328), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n783), .A2(new_n695), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n741), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(new_n786), .B2(G92gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n741), .A2(new_n247), .A3(new_n328), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n780), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n772), .B2(new_n777), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n247), .B1(new_n785), .B2(new_n473), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n790), .B(KEYINPUT52), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT52), .B1(new_n791), .B2(new_n792), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT114), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n789), .A2(new_n793), .A3(new_n795), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n756), .B2(new_n420), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n329), .A2(G99gat), .A3(new_n417), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n780), .B2(new_n798), .ZN(G1338gat));
  INV_X1    g598(.A(G106gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n785), .B2(new_n562), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(KEYINPUT53), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n329), .A2(new_n563), .A3(G106gat), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n780), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT51), .B1(new_n775), .B2(new_n776), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n803), .B1(new_n770), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G106gat), .B1(new_n756), .B2(new_n563), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT115), .B1(new_n809), .B2(KEYINPUT53), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n804), .B1(new_n772), .B2(new_n777), .ZN(new_n811));
  OAI211_X1 g610(.A(KEYINPUT115), .B(KEYINPUT53), .C1(new_n811), .C2(new_n801), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n805), .B1(new_n810), .B2(new_n813), .ZN(G1339gat));
  NOR2_X1   g613(.A1(new_n330), .A2(new_n652), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n630), .B1(new_n629), .B2(new_n631), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n634), .A2(new_n635), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n816), .A2(new_n817), .B1(new_n818), .B2(new_n633), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n816), .A2(new_n817), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n640), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n309), .A2(new_n647), .A3(new_n328), .A4(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT92), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n648), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n643), .A2(KEYINPUT92), .A3(new_n644), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n826), .A2(new_n642), .B1(new_n305), .B2(new_n308), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n827), .A2(new_n821), .B1(new_n652), .B2(new_n309), .ZN(new_n828));
  INV_X1    g627(.A(new_n327), .ZN(new_n829));
  XNOR2_X1  g628(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n326), .B1(new_n320), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n317), .A2(new_n319), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(KEYINPUT54), .A3(new_n325), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n325), .A2(KEYINPUT54), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT116), .B1(new_n836), .B2(new_n832), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n831), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n829), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT55), .B(new_n831), .C1(new_n835), .C2(new_n837), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n831), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n833), .A2(new_n834), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n836), .A2(KEYINPUT116), .A3(new_n832), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT118), .B1(new_n847), .B2(KEYINPUT55), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n840), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n822), .B1(new_n828), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n243), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n815), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n659), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n616), .A3(new_n740), .ZN(new_n854));
  OAI21_X1  g653(.A(G113gat), .B1(new_n854), .B2(new_n655), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n652), .A2(new_n372), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT120), .Z(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n854), .B2(new_n857), .ZN(G1340gat));
  NOR2_X1   g657(.A1(new_n854), .A2(new_n329), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(new_n370), .ZN(G1341gat));
  NOR2_X1   g659(.A1(new_n854), .A2(new_n851), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(new_n378), .ZN(G1342gat));
  NOR4_X1   g661(.A1(new_n852), .A2(new_n659), .A3(new_n473), .A4(new_n309), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n380), .A3(new_n616), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT56), .Z(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n854), .B2(new_n309), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1343gat));
  OAI21_X1  g666(.A(KEYINPUT57), .B1(new_n852), .B2(new_n563), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n741), .A2(new_n659), .A3(new_n674), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n690), .A2(new_n821), .A3(new_n647), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n655), .B2(new_n690), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n327), .B1(new_n847), .B2(KEYINPUT55), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n841), .A2(new_n842), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n847), .A2(KEYINPUT118), .A3(KEYINPUT55), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n243), .B1(new_n877), .B2(new_n822), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n870), .B(new_n562), .C1(new_n878), .C2(new_n815), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n868), .A2(new_n869), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT121), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n868), .A2(new_n879), .A3(new_n882), .A4(new_n869), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n652), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G141gat), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n674), .A2(new_n563), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n655), .A2(G141gat), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n853), .A2(new_n740), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT58), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n853), .A2(new_n740), .A3(new_n886), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n884), .A2(G141gat), .B1(new_n893), .B2(new_n887), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT122), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  XOR2_X1   g695(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n897));
  AND2_X1   g696(.A1(new_n888), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G141gat), .B1(new_n880), .B2(new_n655), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n900), .B(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n891), .A2(new_n896), .A3(new_n902), .ZN(G1344gat));
  INV_X1    g702(.A(G148gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n893), .A2(new_n904), .A3(new_n328), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n881), .A2(new_n328), .A3(new_n883), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(KEYINPUT59), .A3(new_n904), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n868), .A2(new_n879), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n328), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n869), .B(KEYINPUT125), .ZN(new_n910));
  OAI21_X1  g709(.A(G148gat), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(KEYINPUT59), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n905), .B1(new_n907), .B2(new_n912), .ZN(G1345gat));
  NAND3_X1  g712(.A1(new_n881), .A2(new_n243), .A3(new_n883), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G155gat), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n851), .A2(G155gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n892), .B2(new_n916), .ZN(G1346gat));
  INV_X1    g716(.A(G162gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n863), .A2(new_n918), .A3(new_n886), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n881), .A2(new_n690), .A3(new_n883), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n918), .ZN(G1347gat));
  NOR3_X1   g720(.A1(new_n852), .A2(new_n660), .A3(new_n740), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(new_n616), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n333), .A3(new_n652), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  INV_X1    g726(.A(new_n852), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n659), .A2(new_n473), .A3(new_n616), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n655), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n926), .A2(new_n927), .A3(new_n932), .ZN(G1348gat));
  NAND3_X1  g732(.A1(new_n923), .A2(new_n334), .A3(new_n328), .ZN(new_n934));
  OAI21_X1  g733(.A(G176gat), .B1(new_n931), .B2(new_n329), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1349gat));
  NAND3_X1  g735(.A1(new_n923), .A2(new_n360), .A3(new_n243), .ZN(new_n937));
  OAI21_X1  g736(.A(G183gat), .B1(new_n931), .B2(new_n851), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n931), .B2(new_n309), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n941), .A2(KEYINPUT127), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(KEYINPUT127), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n923), .A2(new_n361), .A3(new_n690), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(G1351gat));
  NAND2_X1  g747(.A1(new_n922), .A2(new_n886), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n652), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n420), .A2(new_n659), .A3(new_n473), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n908), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n655), .A2(new_n421), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(G1352gat));
  NOR3_X1   g755(.A1(new_n949), .A2(G204gat), .A3(new_n329), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n909), .B2(new_n952), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n950), .A2(new_n424), .A3(new_n243), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n954), .A2(new_n243), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n425), .A3(new_n690), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n954), .A2(new_n690), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n425), .ZN(G1355gat));
endmodule


