

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772;

  INV_X1 U383 ( .A(G953), .ZN(n628) );
  INV_X1 U384 ( .A(n570), .ZN(n692) );
  NOR2_X1 U385 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U386 ( .A(KEYINPUT24), .B(G110), .Z(n362) );
  XOR2_X1 U387 ( .A(n538), .B(n537), .Z(n363) );
  NOR2_X2 U388 ( .A1(n381), .A2(n608), .ZN(n380) );
  XNOR2_X2 U389 ( .A(n606), .B(KEYINPUT32), .ZN(n769) );
  AND2_X2 U390 ( .A1(n605), .A2(n369), .ZN(n601) );
  XNOR2_X2 U391 ( .A(n407), .B(n406), .ZN(n771) );
  XNOR2_X2 U392 ( .A(n383), .B(KEYINPUT16), .ZN(n397) );
  XNOR2_X2 U393 ( .A(n555), .B(KEYINPUT1), .ZN(n685) );
  NOR2_X1 U394 ( .A1(n612), .A2(n431), .ZN(n404) );
  XNOR2_X1 U395 ( .A(n476), .B(n475), .ZN(n535) );
  NOR2_X1 U396 ( .A1(G953), .A2(n670), .ZN(n673) );
  AND2_X2 U397 ( .A1(n401), .A2(n664), .ZN(n738) );
  AND2_X1 U398 ( .A1(n386), .A2(n411), .ZN(n385) );
  NOR2_X1 U399 ( .A1(n547), .A2(n548), .ZN(n439) );
  NOR2_X1 U400 ( .A1(n562), .A2(n650), .ZN(n563) );
  XNOR2_X1 U401 ( .A(n425), .B(n424), .ZN(n768) );
  NAND2_X1 U402 ( .A1(n393), .A2(n391), .ZN(n569) );
  XNOR2_X1 U403 ( .A(n404), .B(n372), .ZN(n600) );
  NOR2_X1 U404 ( .A1(n586), .A2(n394), .ZN(n395) );
  XNOR2_X1 U405 ( .A(n535), .B(n534), .ZN(n689) );
  XNOR2_X1 U406 ( .A(n570), .B(KEYINPUT6), .ZN(n602) );
  XNOR2_X1 U407 ( .A(n750), .B(n366), .ZN(n374) );
  XOR2_X2 U408 ( .A(n510), .B(n498), .Z(n485) );
  XNOR2_X1 U409 ( .A(n479), .B(n447), .ZN(n509) );
  XNOR2_X1 U410 ( .A(n446), .B(G128), .ZN(n479) );
  XOR2_X1 U411 ( .A(G902), .B(KEYINPUT15), .Z(n619) );
  OR2_X1 U412 ( .A1(n388), .A2(n370), .ZN(n384) );
  BUF_X1 U413 ( .A(n716), .Z(n364) );
  XNOR2_X1 U414 ( .A(n374), .B(n487), .ZN(n716) );
  NAND2_X1 U415 ( .A1(n385), .A2(n384), .ZN(n666) );
  NOR2_X1 U416 ( .A1(G237), .A2(G902), .ZN(n489) );
  XNOR2_X1 U417 ( .A(n435), .B(G101), .ZN(n453) );
  INV_X1 U418 ( .A(KEYINPUT4), .ZN(n435) );
  XOR2_X1 U419 ( .A(G137), .B(G140), .Z(n472) );
  NOR2_X1 U420 ( .A1(n557), .A2(n558), .ZN(n593) );
  AND2_X1 U421 ( .A1(n443), .A2(n363), .ZN(n389) );
  NAND2_X1 U422 ( .A1(n716), .A2(n488), .ZN(n373) );
  NAND2_X1 U423 ( .A1(n378), .A2(n377), .ZN(n376) );
  XNOR2_X1 U424 ( .A(n420), .B(n503), .ZN(n625) );
  XNOR2_X1 U425 ( .A(n421), .B(n497), .ZN(n420) );
  NAND2_X1 U426 ( .A1(n616), .A2(KEYINPUT44), .ZN(n382) );
  INV_X1 U427 ( .A(KEYINPUT64), .ZN(n607) );
  XNOR2_X1 U428 ( .A(n410), .B(G146), .ZN(n486) );
  INV_X1 U429 ( .A(G125), .ZN(n410) );
  NOR2_X1 U430 ( .A1(n413), .A2(n412), .ZN(n411) );
  INV_X1 U431 ( .A(n661), .ZN(n412) );
  NOR2_X1 U432 ( .A1(n662), .A2(KEYINPUT79), .ZN(n413) );
  INV_X1 U433 ( .A(KEYINPUT38), .ZN(n402) );
  XNOR2_X1 U434 ( .A(n616), .B(n615), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n768), .B(n423), .ZN(n377) );
  INV_X1 U436 ( .A(KEYINPUT44), .ZN(n423) );
  XNOR2_X1 U437 ( .A(n486), .B(n471), .ZN(n494) );
  XNOR2_X1 U438 ( .A(n470), .B(KEYINPUT68), .ZN(n471) );
  INV_X1 U439 ( .A(KEYINPUT10), .ZN(n470) );
  INV_X1 U440 ( .A(G143), .ZN(n446) );
  INV_X1 U441 ( .A(n602), .ZN(n609) );
  XNOR2_X1 U442 ( .A(KEYINPUT30), .B(KEYINPUT102), .ZN(n537) );
  INV_X1 U443 ( .A(KEYINPUT67), .ZN(n436) );
  XNOR2_X1 U444 ( .A(n452), .B(n428), .ZN(n555) );
  INV_X1 U445 ( .A(G469), .ZN(n428) );
  NOR2_X1 U446 ( .A1(n737), .A2(G902), .ZN(n476) );
  XNOR2_X1 U447 ( .A(n453), .B(n434), .ZN(n482) );
  XNOR2_X1 U448 ( .A(G110), .B(KEYINPUT70), .ZN(n434) );
  XNOR2_X1 U449 ( .A(n472), .B(n445), .ZN(n448) );
  BUF_X1 U450 ( .A(n666), .Z(n758) );
  XNOR2_X1 U451 ( .A(n613), .B(KEYINPUT34), .ZN(n427) );
  XNOR2_X1 U452 ( .A(n553), .B(n493), .ZN(n375) );
  XNOR2_X1 U453 ( .A(n505), .B(n504), .ZN(n558) );
  XNOR2_X1 U454 ( .A(n429), .B(n456), .ZN(n633) );
  XNOR2_X1 U455 ( .A(n455), .B(n461), .ZN(n429) );
  XOR2_X1 U456 ( .A(KEYINPUT84), .B(n629), .Z(n724) );
  INV_X1 U457 ( .A(KEYINPUT40), .ZN(n406) );
  XOR2_X1 U458 ( .A(KEYINPUT69), .B(G131), .Z(n499) );
  INV_X1 U459 ( .A(KEYINPUT79), .ZN(n387) );
  XNOR2_X1 U460 ( .A(n382), .B(n607), .ZN(n381) );
  NOR2_X1 U461 ( .A1(G237), .A2(G953), .ZN(n459) );
  XNOR2_X1 U462 ( .A(KEYINPUT91), .B(KEYINPUT11), .ZN(n422) );
  XNOR2_X1 U463 ( .A(G143), .B(G122), .ZN(n495) );
  XOR2_X1 U464 ( .A(KEYINPUT12), .B(G140), .Z(n496) );
  NAND2_X1 U465 ( .A1(n363), .A2(n396), .ZN(n394) );
  NOR2_X1 U466 ( .A1(n674), .A2(n444), .ZN(n443) );
  NAND2_X1 U467 ( .A1(n593), .A2(n432), .ZN(n431) );
  INV_X1 U468 ( .A(n592), .ZN(n432) );
  XOR2_X1 U469 ( .A(G137), .B(KEYINPUT89), .Z(n458) );
  XNOR2_X1 U470 ( .A(n453), .B(n405), .ZN(n398) );
  XNOR2_X1 U471 ( .A(n494), .B(n472), .ZN(n756) );
  XNOR2_X1 U472 ( .A(n442), .B(KEYINPUT86), .ZN(n441) );
  INV_X1 U473 ( .A(KEYINPUT23), .ZN(n442) );
  XNOR2_X1 U474 ( .A(n400), .B(n399), .ZN(n511) );
  INV_X1 U475 ( .A(KEYINPUT8), .ZN(n399) );
  NAND2_X1 U476 ( .A1(n628), .A2(G234), .ZN(n400) );
  INV_X1 U477 ( .A(G134), .ZN(n447) );
  NOR2_X1 U478 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U479 ( .A(n418), .B(n542), .ZN(n702) );
  NAND2_X1 U480 ( .A1(n415), .A2(n555), .ZN(n543) );
  XNOR2_X1 U481 ( .A(n416), .B(n478), .ZN(n415) );
  NOR2_X1 U482 ( .A1(n549), .A2(n570), .ZN(n416) );
  INV_X1 U483 ( .A(KEYINPUT0), .ZN(n433) );
  INV_X1 U484 ( .A(KEYINPUT25), .ZN(n534) );
  XNOR2_X1 U485 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U486 ( .A(G104), .B(G107), .ZN(n450) );
  XNOR2_X1 U487 ( .A(n482), .B(n448), .ZN(n449) );
  XNOR2_X1 U488 ( .A(n718), .B(n717), .ZN(n719) );
  NAND2_X1 U489 ( .A1(n568), .A2(n430), .ZN(n662) );
  XOR2_X1 U490 ( .A(KEYINPUT42), .B(n544), .Z(n770) );
  NAND2_X1 U491 ( .A1(n417), .A2(n414), .ZN(n544) );
  INV_X1 U492 ( .A(n543), .ZN(n414) );
  INV_X1 U493 ( .A(n702), .ZN(n417) );
  INV_X1 U494 ( .A(KEYINPUT35), .ZN(n424) );
  NAND2_X1 U495 ( .A1(n427), .A2(n426), .ZN(n425) );
  INV_X1 U496 ( .A(n614), .ZN(n426) );
  XOR2_X1 U497 ( .A(KEYINPUT96), .B(n521), .Z(n652) );
  NOR2_X1 U498 ( .A1(n559), .A2(n430), .ZN(n560) );
  XOR2_X1 U499 ( .A(n633), .B(KEYINPUT62), .Z(n635) );
  XNOR2_X1 U500 ( .A(KEYINPUT80), .B(KEYINPUT39), .ZN(n365) );
  XOR2_X1 U501 ( .A(n486), .B(KEYINPUT17), .Z(n366) );
  XNOR2_X1 U502 ( .A(n755), .B(G146), .ZN(n456) );
  XOR2_X1 U503 ( .A(n458), .B(n457), .Z(n367) );
  XOR2_X1 U504 ( .A(n491), .B(n490), .Z(n368) );
  NOR2_X1 U505 ( .A1(n685), .A2(n692), .ZN(n369) );
  NAND2_X1 U506 ( .A1(n662), .A2(KEYINPUT79), .ZN(n370) );
  AND2_X1 U507 ( .A1(n390), .A2(n363), .ZN(n371) );
  INV_X2 U508 ( .A(G113), .ZN(n405) );
  XOR2_X1 U509 ( .A(n594), .B(KEYINPUT71), .Z(n372) );
  INV_X1 U510 ( .A(n365), .ZN(n396) );
  XNOR2_X1 U511 ( .A(n509), .B(n499), .ZN(n755) );
  XNOR2_X2 U512 ( .A(n373), .B(n368), .ZN(n540) );
  NOR2_X2 U513 ( .A1(n375), .A2(n584), .ZN(n409) );
  NOR2_X1 U514 ( .A1(n543), .A2(n375), .ZN(n651) );
  NAND2_X1 U515 ( .A1(n380), .A2(n376), .ZN(n618) );
  NAND2_X1 U516 ( .A1(n379), .A2(n768), .ZN(n378) );
  XNOR2_X1 U517 ( .A(n398), .B(n383), .ZN(n455) );
  XNOR2_X2 U518 ( .A(n454), .B(G119), .ZN(n383) );
  NAND2_X1 U519 ( .A1(n388), .A2(n387), .ZN(n386) );
  XNOR2_X1 U520 ( .A(n438), .B(KEYINPUT48), .ZN(n388) );
  NAND2_X1 U521 ( .A1(n390), .A2(n389), .ZN(n392) );
  INV_X1 U522 ( .A(n586), .ZN(n390) );
  XNOR2_X2 U523 ( .A(n536), .B(KEYINPUT88), .ZN(n586) );
  NAND2_X1 U524 ( .A1(n392), .A2(n365), .ZN(n391) );
  NAND2_X1 U525 ( .A1(n395), .A2(n443), .ZN(n393) );
  NOR2_X1 U526 ( .A1(n771), .A2(n770), .ZN(n546) );
  NAND2_X1 U527 ( .A1(n569), .A2(n652), .ZN(n407) );
  XNOR2_X2 U528 ( .A(n397), .B(n485), .ZN(n750) );
  XOR2_X2 U529 ( .A(G107), .B(G122), .Z(n510) );
  NAND2_X1 U530 ( .A1(n439), .A2(n563), .ZN(n438) );
  XNOR2_X1 U531 ( .A(n408), .B(n756), .ZN(n737) );
  XNOR2_X2 U532 ( .A(n409), .B(n433), .ZN(n612) );
  NAND2_X1 U533 ( .A1(n622), .A2(n621), .ZN(n401) );
  NAND2_X1 U534 ( .A1(n540), .A2(n675), .ZN(n553) );
  NOR2_X1 U535 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U536 ( .A(n535), .B(KEYINPUT25), .ZN(n599) );
  NAND2_X1 U537 ( .A1(n477), .A2(n539), .ZN(n549) );
  XNOR2_X1 U538 ( .A(n469), .B(n441), .ZN(n440) );
  XNOR2_X1 U539 ( .A(n440), .B(n473), .ZN(n408) );
  NAND2_X1 U540 ( .A1(n738), .A2(G210), .ZN(n720) );
  XNOR2_X2 U541 ( .A(n601), .B(KEYINPUT99), .ZN(n767) );
  NAND2_X1 U542 ( .A1(n541), .A2(n675), .ZN(n678) );
  XNOR2_X1 U543 ( .A(n540), .B(n402), .ZN(n541) );
  NAND2_X2 U544 ( .A1(n767), .A2(n769), .ZN(n616) );
  NAND2_X1 U545 ( .A1(n403), .A2(n724), .ZN(n636) );
  XNOR2_X1 U546 ( .A(n634), .B(n635), .ZN(n403) );
  NOR2_X2 U547 ( .A1(n600), .A2(n599), .ZN(n605) );
  XNOR2_X2 U548 ( .A(n405), .B(G104), .ZN(n498) );
  INV_X1 U549 ( .A(n593), .ZN(n677) );
  NAND2_X1 U550 ( .A1(n419), .A2(n593), .ZN(n418) );
  INV_X1 U551 ( .A(n678), .ZN(n419) );
  XNOR2_X1 U552 ( .A(n494), .B(n422), .ZN(n421) );
  NAND2_X1 U553 ( .A1(n684), .A2(n685), .ZN(n610) );
  XNOR2_X2 U554 ( .A(n462), .B(G472), .ZN(n570) );
  XNOR2_X2 U555 ( .A(n618), .B(n617), .ZN(n746) );
  XNOR2_X2 U556 ( .A(G116), .B(KEYINPUT3), .ZN(n454) );
  INV_X1 U557 ( .A(n540), .ZN(n430) );
  NAND2_X1 U558 ( .A1(n684), .A2(n555), .ZN(n536) );
  XNOR2_X2 U559 ( .A(n437), .B(n436), .ZN(n684) );
  NOR2_X2 U560 ( .A1(n689), .A2(n592), .ZN(n437) );
  NAND2_X1 U561 ( .A1(n371), .A2(n539), .ZN(n559) );
  INV_X1 U562 ( .A(n539), .ZN(n444) );
  XNOR2_X1 U563 ( .A(n546), .B(n545), .ZN(n547) );
  AND2_X1 U564 ( .A1(G227), .A2(n628), .ZN(n445) );
  INV_X1 U565 ( .A(KEYINPUT46), .ZN(n545) );
  INV_X1 U566 ( .A(n660), .ZN(n562) );
  INV_X1 U567 ( .A(KEYINPUT81), .ZN(n615) );
  XNOR2_X1 U568 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U569 ( .A(n367), .B(n460), .ZN(n461) );
  XNOR2_X1 U570 ( .A(n502), .B(n501), .ZN(n503) );
  INV_X1 U571 ( .A(KEYINPUT75), .ZN(n490) );
  INV_X1 U572 ( .A(KEYINPUT19), .ZN(n493) );
  XNOR2_X1 U573 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U574 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U575 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U576 ( .A(n456), .B(n451), .ZN(n727) );
  NOR2_X1 U577 ( .A1(G902), .A2(n727), .ZN(n452) );
  XNOR2_X1 U578 ( .A(KEYINPUT73), .B(KEYINPUT5), .ZN(n457) );
  XNOR2_X1 U579 ( .A(n459), .B(KEYINPUT74), .ZN(n500) );
  NAND2_X1 U580 ( .A1(G210), .A2(n500), .ZN(n460) );
  NOR2_X1 U581 ( .A1(n633), .A2(G902), .ZN(n462) );
  INV_X1 U582 ( .A(G952), .ZN(n710) );
  NOR2_X1 U583 ( .A1(G953), .A2(n710), .ZN(n571) );
  NAND2_X1 U584 ( .A1(G953), .A2(G902), .ZN(n572) );
  NOR2_X1 U585 ( .A1(G900), .A2(n572), .ZN(n463) );
  NOR2_X1 U586 ( .A1(n571), .A2(n463), .ZN(n465) );
  NAND2_X1 U587 ( .A1(G234), .A2(G237), .ZN(n464) );
  XOR2_X1 U588 ( .A(KEYINPUT14), .B(n464), .Z(n575) );
  NOR2_X1 U589 ( .A1(n465), .A2(n575), .ZN(n539) );
  INV_X1 U590 ( .A(n619), .ZN(n488) );
  NAND2_X1 U591 ( .A1(n488), .A2(G234), .ZN(n466) );
  XNOR2_X1 U592 ( .A(n466), .B(KEYINPUT20), .ZN(n474) );
  NAND2_X1 U593 ( .A1(G221), .A2(n474), .ZN(n467) );
  XNOR2_X1 U594 ( .A(KEYINPUT21), .B(n467), .ZN(n688) );
  XNOR2_X1 U595 ( .A(G128), .B(G119), .ZN(n468) );
  XNOR2_X1 U596 ( .A(n362), .B(n468), .ZN(n469) );
  AND2_X1 U597 ( .A1(n511), .A2(G221), .ZN(n473) );
  NAND2_X1 U598 ( .A1(G217), .A2(n474), .ZN(n475) );
  NOR2_X1 U599 ( .A1(n688), .A2(n599), .ZN(n477) );
  XNOR2_X1 U600 ( .A(KEYINPUT104), .B(KEYINPUT28), .ZN(n478) );
  AND2_X1 U601 ( .A1(G224), .A2(n628), .ZN(n480) );
  XNOR2_X1 U602 ( .A(n482), .B(n481), .ZN(n484) );
  INV_X1 U603 ( .A(KEYINPUT18), .ZN(n483) );
  XNOR2_X1 U604 ( .A(n484), .B(n483), .ZN(n487) );
  XOR2_X1 U605 ( .A(KEYINPUT72), .B(n489), .Z(n492) );
  NAND2_X1 U606 ( .A1(n492), .A2(G210), .ZN(n491) );
  NAND2_X1 U607 ( .A1(n492), .A2(G214), .ZN(n675) );
  INV_X1 U608 ( .A(n651), .ZN(n645) );
  NAND2_X1 U609 ( .A1(n645), .A2(KEYINPUT76), .ZN(n523) );
  XNOR2_X1 U610 ( .A(KEYINPUT13), .B(G475), .ZN(n505) );
  XNOR2_X1 U611 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U612 ( .A(n499), .B(n498), .ZN(n502) );
  NAND2_X1 U613 ( .A1(n500), .A2(G214), .ZN(n501) );
  NOR2_X1 U614 ( .A1(G902), .A2(n625), .ZN(n504) );
  XNOR2_X1 U615 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n517) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(KEYINPUT92), .Z(n507) );
  XNOR2_X1 U617 ( .A(G116), .B(KEYINPUT7), .ZN(n506) );
  XNOR2_X1 U618 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U619 ( .A(n509), .B(n508), .ZN(n515) );
  XOR2_X1 U620 ( .A(n510), .B(KEYINPUT93), .Z(n513) );
  NAND2_X1 U621 ( .A1(G217), .A2(n511), .ZN(n512) );
  XNOR2_X1 U622 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U623 ( .A(n515), .B(n514), .ZN(n733) );
  NOR2_X1 U624 ( .A1(G902), .A2(n733), .ZN(n516) );
  XNOR2_X1 U625 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U626 ( .A(G478), .B(n518), .ZN(n557) );
  INV_X1 U627 ( .A(n557), .ZN(n520) );
  NOR2_X1 U628 ( .A1(n558), .A2(n520), .ZN(n519) );
  XOR2_X1 U629 ( .A(KEYINPUT97), .B(n519), .Z(n641) );
  NAND2_X1 U630 ( .A1(n558), .A2(n520), .ZN(n521) );
  NOR2_X1 U631 ( .A1(n641), .A2(n652), .ZN(n679) );
  INV_X1 U632 ( .A(n679), .ZN(n590) );
  OR2_X1 U633 ( .A1(n590), .A2(KEYINPUT77), .ZN(n522) );
  NAND2_X1 U634 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U635 ( .A1(n524), .A2(KEYINPUT47), .ZN(n526) );
  OR2_X1 U636 ( .A1(KEYINPUT76), .A2(n645), .ZN(n525) );
  NAND2_X1 U637 ( .A1(n526), .A2(n525), .ZN(n531) );
  NAND2_X1 U638 ( .A1(n651), .A2(n590), .ZN(n527) );
  NAND2_X1 U639 ( .A1(KEYINPUT76), .A2(n527), .ZN(n528) );
  NOR2_X1 U640 ( .A1(KEYINPUT77), .A2(n528), .ZN(n529) );
  NOR2_X1 U641 ( .A1(KEYINPUT47), .A2(n529), .ZN(n530) );
  NOR2_X1 U642 ( .A1(n531), .A2(n530), .ZN(n533) );
  NAND2_X1 U643 ( .A1(KEYINPUT77), .A2(n590), .ZN(n532) );
  NAND2_X1 U644 ( .A1(n533), .A2(n532), .ZN(n548) );
  XOR2_X1 U645 ( .A(KEYINPUT87), .B(n688), .Z(n592) );
  NAND2_X1 U646 ( .A1(n692), .A2(n675), .ZN(n538) );
  INV_X1 U647 ( .A(n541), .ZN(n674) );
  XNOR2_X1 U648 ( .A(KEYINPUT105), .B(KEYINPUT41), .ZN(n542) );
  NOR2_X1 U649 ( .A1(n609), .A2(n549), .ZN(n550) );
  XNOR2_X1 U650 ( .A(n550), .B(KEYINPUT100), .ZN(n551) );
  NAND2_X1 U651 ( .A1(n551), .A2(n652), .ZN(n564) );
  XNOR2_X1 U652 ( .A(KEYINPUT106), .B(n564), .ZN(n552) );
  XNOR2_X1 U653 ( .A(n554), .B(KEYINPUT36), .ZN(n556) );
  NAND2_X1 U654 ( .A1(n556), .A2(n685), .ZN(n660) );
  NAND2_X1 U655 ( .A1(n558), .A2(n557), .ZN(n614) );
  XNOR2_X1 U656 ( .A(n560), .B(KEYINPUT103), .ZN(n561) );
  NOR2_X1 U657 ( .A1(n614), .A2(n561), .ZN(n650) );
  XOR2_X1 U658 ( .A(KEYINPUT43), .B(KEYINPUT101), .Z(n567) );
  NOR2_X1 U659 ( .A1(n685), .A2(n564), .ZN(n565) );
  NAND2_X1 U660 ( .A1(n565), .A2(n675), .ZN(n566) );
  XNOR2_X1 U661 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U662 ( .A1(n641), .A2(n569), .ZN(n661) );
  OR2_X1 U663 ( .A1(n570), .A2(n610), .ZN(n697) );
  INV_X1 U664 ( .A(n571), .ZN(n574) );
  OR2_X1 U665 ( .A1(n572), .A2(G898), .ZN(n573) );
  NAND2_X1 U666 ( .A1(n574), .A2(n573), .ZN(n576) );
  INV_X1 U667 ( .A(n575), .ZN(n707) );
  NAND2_X1 U668 ( .A1(n576), .A2(n707), .ZN(n578) );
  INV_X1 U669 ( .A(KEYINPUT85), .ZN(n577) );
  NAND2_X1 U670 ( .A1(n578), .A2(n577), .ZN(n583) );
  INV_X1 U671 ( .A(G902), .ZN(n580) );
  NOR2_X1 U672 ( .A1(G898), .A2(n628), .ZN(n752) );
  NAND2_X1 U673 ( .A1(n752), .A2(KEYINPUT85), .ZN(n579) );
  NOR2_X1 U674 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U675 ( .A1(n581), .A2(n707), .ZN(n582) );
  NAND2_X1 U676 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U677 ( .A1(n697), .A2(n612), .ZN(n585) );
  XNOR2_X1 U678 ( .A(n585), .B(KEYINPUT31), .ZN(n656) );
  INV_X1 U679 ( .A(n612), .ZN(n588) );
  NOR2_X1 U680 ( .A1(n586), .A2(n692), .ZN(n587) );
  NAND2_X1 U681 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U682 ( .A(KEYINPUT90), .B(n589), .ZN(n642) );
  NAND2_X1 U683 ( .A1(n656), .A2(n642), .ZN(n591) );
  NAND2_X1 U684 ( .A1(n591), .A2(n590), .ZN(n598) );
  XNOR2_X1 U685 ( .A(KEYINPUT22), .B(KEYINPUT65), .ZN(n594) );
  NOR2_X1 U686 ( .A1(n602), .A2(n600), .ZN(n596) );
  NOR2_X1 U687 ( .A1(n685), .A2(n689), .ZN(n595) );
  NAND2_X1 U688 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U689 ( .A(KEYINPUT98), .B(n597), .ZN(n772) );
  NAND2_X1 U690 ( .A1(n598), .A2(n772), .ZN(n608) );
  INV_X1 U691 ( .A(n685), .ZN(n603) );
  NOR2_X1 U692 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U693 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U694 ( .A(n611), .B(KEYINPUT33), .ZN(n682) );
  NOR2_X1 U695 ( .A1(n612), .A2(n682), .ZN(n613) );
  INV_X1 U696 ( .A(KEYINPUT45), .ZN(n617) );
  NOR2_X2 U697 ( .A1(n666), .A2(n746), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n623), .A2(n619), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n619), .A2(KEYINPUT2), .ZN(n620) );
  XNOR2_X1 U700 ( .A(KEYINPUT66), .B(n620), .ZN(n621) );
  NAND2_X1 U701 ( .A1(KEYINPUT2), .A2(n623), .ZN(n664) );
  NAND2_X1 U702 ( .A1(n738), .A2(G475), .ZN(n627) );
  XOR2_X1 U703 ( .A(KEYINPUT59), .B(KEYINPUT121), .Z(n624) );
  XNOR2_X1 U704 ( .A(n627), .B(n626), .ZN(n630) );
  NOR2_X1 U705 ( .A1(G952), .A2(n628), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n724), .ZN(n632) );
  INV_X1 U707 ( .A(KEYINPUT60), .ZN(n631) );
  XNOR2_X1 U708 ( .A(n632), .B(n631), .ZN(G60) );
  NAND2_X1 U709 ( .A1(n738), .A2(G472), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n636), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U711 ( .A(G104), .B(KEYINPUT107), .ZN(n638) );
  INV_X1 U712 ( .A(n652), .ZN(n654) );
  NOR2_X1 U713 ( .A1(n654), .A2(n642), .ZN(n637) );
  XNOR2_X1 U714 ( .A(n638), .B(n637), .ZN(G6) );
  XOR2_X1 U715 ( .A(KEYINPUT108), .B(KEYINPUT26), .Z(n640) );
  XNOR2_X1 U716 ( .A(G107), .B(KEYINPUT27), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n640), .B(n639), .ZN(n644) );
  INV_X1 U718 ( .A(n641), .ZN(n657) );
  NOR2_X1 U719 ( .A1(n642), .A2(n657), .ZN(n643) );
  XOR2_X1 U720 ( .A(n644), .B(n643), .Z(G9) );
  NOR2_X1 U721 ( .A1(n645), .A2(n657), .ZN(n649) );
  XOR2_X1 U722 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n647) );
  XNOR2_X1 U723 ( .A(G128), .B(KEYINPUT29), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U725 ( .A(n649), .B(n648), .ZN(G30) );
  XOR2_X1 U726 ( .A(G143), .B(n650), .Z(G45) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n653), .B(G146), .ZN(G48) );
  NOR2_X1 U729 ( .A1(n654), .A2(n656), .ZN(n655) );
  XOR2_X1 U730 ( .A(G113), .B(n655), .Z(G15) );
  NOR2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U732 ( .A(G116), .B(n658), .Z(G18) );
  XOR2_X1 U733 ( .A(G125), .B(KEYINPUT37), .Z(n659) );
  XNOR2_X1 U734 ( .A(n660), .B(n659), .ZN(G27) );
  XNOR2_X1 U735 ( .A(G134), .B(n661), .ZN(G36) );
  XNOR2_X1 U736 ( .A(G140), .B(n662), .ZN(G42) );
  INV_X1 U737 ( .A(KEYINPUT2), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n746), .A2(n667), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(KEYINPUT78), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n665), .A2(n664), .ZN(n669) );
  AND2_X1 U741 ( .A1(n758), .A2(n667), .ZN(n668) );
  NOR2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U743 ( .A1(n702), .A2(n682), .ZN(n671) );
  XOR2_X1 U744 ( .A(KEYINPUT116), .B(n671), .Z(n672) );
  NAND2_X1 U745 ( .A1(n673), .A2(n672), .ZN(n712) );
  NOR2_X1 U746 ( .A1(n541), .A2(n675), .ZN(n676) );
  NOR2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n704) );
  XOR2_X1 U751 ( .A(KEYINPUT50), .B(KEYINPUT112), .Z(n687) );
  OR2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U753 ( .A(n687), .B(n686), .ZN(n695) );
  NAND2_X1 U754 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U755 ( .A(KEYINPUT49), .B(n690), .ZN(n691) );
  NOR2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U757 ( .A(n693), .B(KEYINPUT111), .ZN(n694) );
  NOR2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U759 ( .A(KEYINPUT113), .B(n696), .ZN(n698) );
  NAND2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U761 ( .A(n699), .B(KEYINPUT51), .ZN(n700) );
  XNOR2_X1 U762 ( .A(KEYINPUT114), .B(n700), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U765 ( .A(n705), .B(KEYINPUT115), .ZN(n706) );
  XNOR2_X1 U766 ( .A(n706), .B(KEYINPUT52), .ZN(n708) );
  NAND2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U768 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U769 ( .A(KEYINPUT53), .B(n713), .ZN(G75) );
  XNOR2_X1 U770 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n714) );
  XNOR2_X1 U771 ( .A(n714), .B(KEYINPUT55), .ZN(n715) );
  XOR2_X1 U772 ( .A(n715), .B(KEYINPUT117), .Z(n718) );
  XNOR2_X1 U773 ( .A(n364), .B(KEYINPUT54), .ZN(n717) );
  XNOR2_X1 U774 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U775 ( .A1(n721), .A2(n724), .ZN(n723) );
  XOR2_X1 U776 ( .A(KEYINPUT118), .B(KEYINPUT56), .Z(n722) );
  XNOR2_X1 U777 ( .A(n723), .B(n722), .ZN(G51) );
  INV_X1 U778 ( .A(n724), .ZN(n741) );
  XOR2_X1 U779 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n726) );
  XNOR2_X1 U780 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n725) );
  XNOR2_X1 U781 ( .A(n726), .B(n725), .ZN(n728) );
  XNOR2_X1 U782 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U783 ( .A1(n738), .A2(G469), .ZN(n729) );
  XOR2_X1 U784 ( .A(n730), .B(n729), .Z(n731) );
  NOR2_X1 U785 ( .A1(n741), .A2(n731), .ZN(G54) );
  NAND2_X1 U786 ( .A1(n738), .A2(G478), .ZN(n735) );
  XOR2_X1 U787 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n732) );
  NOR2_X1 U788 ( .A1(n741), .A2(n736), .ZN(G63) );
  XNOR2_X1 U789 ( .A(n737), .B(KEYINPUT124), .ZN(n740) );
  NAND2_X1 U790 ( .A1(G217), .A2(n738), .ZN(n739) );
  XNOR2_X1 U791 ( .A(n740), .B(n739), .ZN(n742) );
  NOR2_X1 U792 ( .A1(n742), .A2(n741), .ZN(G66) );
  INV_X1 U793 ( .A(G898), .ZN(n745) );
  NAND2_X1 U794 ( .A1(G953), .A2(G224), .ZN(n743) );
  XOR2_X1 U795 ( .A(KEYINPUT61), .B(n743), .Z(n744) );
  NOR2_X1 U796 ( .A1(n745), .A2(n744), .ZN(n748) );
  NOR2_X1 U797 ( .A1(G953), .A2(n746), .ZN(n747) );
  NOR2_X1 U798 ( .A1(n748), .A2(n747), .ZN(n754) );
  XOR2_X1 U799 ( .A(G101), .B(G110), .Z(n749) );
  XNOR2_X1 U800 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U801 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U802 ( .A(n754), .B(n753), .Z(G69) );
  XOR2_X1 U803 ( .A(KEYINPUT4), .B(n756), .Z(n757) );
  XOR2_X1 U804 ( .A(n755), .B(n757), .Z(n760) );
  XNOR2_X1 U805 ( .A(n760), .B(n758), .ZN(n759) );
  NOR2_X1 U806 ( .A1(G953), .A2(n759), .ZN(n765) );
  XNOR2_X1 U807 ( .A(KEYINPUT125), .B(n760), .ZN(n761) );
  XNOR2_X1 U808 ( .A(G227), .B(n761), .ZN(n763) );
  NAND2_X1 U809 ( .A1(G900), .A2(G953), .ZN(n762) );
  NOR2_X1 U810 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U811 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U812 ( .A(KEYINPUT126), .B(n766), .ZN(G72) );
  XNOR2_X1 U813 ( .A(n767), .B(G110), .ZN(G12) );
  XNOR2_X1 U814 ( .A(G122), .B(n768), .ZN(G24) );
  XNOR2_X1 U815 ( .A(n769), .B(G119), .ZN(G21) );
  XOR2_X1 U816 ( .A(n770), .B(G137), .Z(G39) );
  XOR2_X1 U817 ( .A(n771), .B(G131), .Z(G33) );
  XNOR2_X1 U818 ( .A(n772), .B(G101), .ZN(G3) );
endmodule

