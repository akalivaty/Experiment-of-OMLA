

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U557 ( .A1(n666), .A2(n665), .ZN(n681) );
  XOR2_X1 U558 ( .A(KEYINPUT17), .B(n525), .Z(n890) );
  NOR2_X2 U559 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X2 U560 ( .A(n654), .B(KEYINPUT29), .ZN(n657) );
  NOR2_X1 U561 ( .A1(n534), .A2(n533), .ZN(n592) );
  NOR2_X1 U562 ( .A1(n588), .A2(n587), .ZN(n589) );
  AND2_X2 U563 ( .A1(n671), .A2(n672), .ZN(n660) );
  NOR2_X1 U564 ( .A1(n664), .A2(n597), .ZN(n599) );
  XOR2_X1 U565 ( .A(KEYINPUT84), .B(n529), .Z(n524) );
  INV_X1 U566 ( .A(KEYINPUT28), .ZN(n617) );
  INV_X1 U567 ( .A(KEYINPUT30), .ZN(n598) );
  XNOR2_X1 U568 ( .A(n531), .B(KEYINPUT66), .ZN(n891) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n530), .ZN(n894) );
  NOR2_X1 U570 ( .A1(G651), .A2(n581), .ZN(n802) );
  XNOR2_X1 U571 ( .A(n762), .B(KEYINPUT103), .ZN(n763) );
  BUF_X1 U572 ( .A(n592), .Z(G164) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  NAND2_X1 U574 ( .A1(G138), .A2(n890), .ZN(n526) );
  XNOR2_X1 U575 ( .A(n526), .B(KEYINPUT85), .ZN(n534) );
  INV_X1 U576 ( .A(G2105), .ZN(n530) );
  NAND2_X1 U577 ( .A1(G126), .A2(n894), .ZN(n528) );
  AND2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  NAND2_X1 U579 ( .A1(G114), .A2(n895), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n529) );
  AND2_X1 U581 ( .A1(G2104), .A2(n530), .ZN(n531) );
  NAND2_X1 U582 ( .A1(G102), .A2(n891), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n524), .A2(n532), .ZN(n533) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n798) );
  NAND2_X1 U585 ( .A1(n798), .A2(G89), .ZN(n535) );
  XNOR2_X1 U586 ( .A(n535), .B(KEYINPUT4), .ZN(n537) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n581) );
  INV_X1 U588 ( .A(G651), .ZN(n539) );
  NOR2_X1 U589 ( .A1(n581), .A2(n539), .ZN(n794) );
  NAND2_X1 U590 ( .A1(G76), .A2(n794), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U592 ( .A(n538), .B(KEYINPUT5), .ZN(n546) );
  XNOR2_X1 U593 ( .A(KEYINPUT75), .B(KEYINPUT6), .ZN(n544) );
  NOR2_X1 U594 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n540), .Z(n795) );
  NAND2_X1 U596 ( .A1(G63), .A2(n795), .ZN(n542) );
  NAND2_X1 U597 ( .A1(G51), .A2(n802), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U599 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U601 ( .A(KEYINPUT7), .B(n547), .ZN(G168) );
  NAND2_X1 U602 ( .A1(G64), .A2(n795), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G52), .A2(n802), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U605 ( .A1(G77), .A2(n794), .ZN(n551) );
  NAND2_X1 U606 ( .A1(G90), .A2(n798), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U608 ( .A(KEYINPUT9), .B(n552), .Z(n553) );
  XNOR2_X1 U609 ( .A(KEYINPUT68), .B(n553), .ZN(n554) );
  NOR2_X1 U610 ( .A1(n555), .A2(n554), .ZN(G171) );
  NAND2_X1 U611 ( .A1(G75), .A2(n794), .ZN(n557) );
  NAND2_X1 U612 ( .A1(G88), .A2(n798), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G62), .A2(n795), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G50), .A2(n802), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U617 ( .A1(n561), .A2(n560), .ZN(G166) );
  INV_X1 U618 ( .A(G166), .ZN(G303) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U620 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n563) );
  NAND2_X1 U621 ( .A1(G73), .A2(n794), .ZN(n562) );
  XNOR2_X1 U622 ( .A(n563), .B(n562), .ZN(n570) );
  NAND2_X1 U623 ( .A1(G61), .A2(n795), .ZN(n565) );
  NAND2_X1 U624 ( .A1(G48), .A2(n802), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G86), .A2(n798), .ZN(n566) );
  XOR2_X1 U627 ( .A(KEYINPUT80), .B(n566), .Z(n567) );
  NOR2_X1 U628 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(G305) );
  NAND2_X1 U630 ( .A1(G72), .A2(n794), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G85), .A2(n798), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U633 ( .A1(G60), .A2(n795), .ZN(n573) );
  XNOR2_X1 U634 ( .A(KEYINPUT67), .B(n573), .ZN(n574) );
  NOR2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n802), .A2(G47), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(G290) );
  NAND2_X1 U638 ( .A1(G49), .A2(n802), .ZN(n579) );
  NAND2_X1 U639 ( .A1(G74), .A2(G651), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U641 ( .A1(n795), .A2(n580), .ZN(n583) );
  NAND2_X1 U642 ( .A1(n581), .A2(G87), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(G288) );
  NAND2_X1 U644 ( .A1(G125), .A2(n894), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G113), .A2(n895), .ZN(n584) );
  AND2_X1 U646 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U647 ( .A1(G101), .A2(n891), .ZN(n586) );
  XNOR2_X1 U648 ( .A(n586), .B(KEYINPUT23), .ZN(n588) );
  AND2_X1 U649 ( .A1(G137), .A2(n890), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X2 U651 ( .A(n591), .B(KEYINPUT65), .ZN(G160) );
  NAND2_X1 U652 ( .A1(G160), .A2(G40), .ZN(n693) );
  INV_X1 U653 ( .A(n693), .ZN(n594) );
  NOR2_X1 U654 ( .A1(G1384), .A2(n592), .ZN(n593) );
  XNOR2_X1 U655 ( .A(n593), .B(KEYINPUT64), .ZN(n692) );
  NAND2_X2 U656 ( .A1(n594), .A2(n692), .ZN(n667) );
  NAND2_X1 U657 ( .A1(n667), .A2(G8), .ZN(n595) );
  XNOR2_X1 U658 ( .A(n595), .B(KEYINPUT94), .ZN(n685) );
  NOR2_X1 U659 ( .A1(n685), .A2(G1966), .ZN(n664) );
  NOR2_X1 U660 ( .A1(G2084), .A2(n667), .ZN(n596) );
  XOR2_X1 U661 ( .A(KEYINPUT96), .B(n596), .Z(n661) );
  NAND2_X1 U662 ( .A1(G8), .A2(n661), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n599), .B(n598), .ZN(n600) );
  NOR2_X1 U664 ( .A1(G168), .A2(n600), .ZN(n604) );
  XNOR2_X1 U665 ( .A(G2078), .B(KEYINPUT25), .ZN(n952) );
  NOR2_X1 U666 ( .A1(n667), .A2(n952), .ZN(n602) );
  INV_X1 U667 ( .A(n667), .ZN(n642) );
  INV_X1 U668 ( .A(G1961), .ZN(n1005) );
  NOR2_X1 U669 ( .A1(n642), .A2(n1005), .ZN(n601) );
  NOR2_X1 U670 ( .A1(n602), .A2(n601), .ZN(n655) );
  NOR2_X1 U671 ( .A1(G171), .A2(n655), .ZN(n603) );
  NOR2_X1 U672 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U673 ( .A(KEYINPUT31), .B(n605), .Z(n671) );
  NAND2_X1 U674 ( .A1(G65), .A2(n795), .ZN(n607) );
  NAND2_X1 U675 ( .A1(G53), .A2(n802), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U677 ( .A1(G78), .A2(n794), .ZN(n609) );
  NAND2_X1 U678 ( .A1(G91), .A2(n798), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U680 ( .A1(n611), .A2(n610), .ZN(n979) );
  INV_X1 U681 ( .A(G2072), .ZN(n954) );
  NOR2_X2 U682 ( .A1(n667), .A2(n954), .ZN(n613) );
  XOR2_X1 U683 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n612) );
  XNOR2_X1 U684 ( .A(n613), .B(n612), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n667), .A2(G1956), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U687 ( .A(n616), .B(KEYINPUT98), .Z(n619) );
  NOR2_X2 U688 ( .A1(n979), .A2(n619), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(n617), .ZN(n653) );
  NAND2_X1 U690 ( .A1(n979), .A2(n619), .ZN(n651) );
  NAND2_X1 U691 ( .A1(G81), .A2(n798), .ZN(n620) );
  XNOR2_X1 U692 ( .A(n620), .B(KEYINPUT12), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n621), .B(KEYINPUT72), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G68), .A2(n794), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U696 ( .A(KEYINPUT13), .B(n624), .ZN(n630) );
  NAND2_X1 U697 ( .A1(G56), .A2(n795), .ZN(n625) );
  XOR2_X1 U698 ( .A(KEYINPUT14), .B(n625), .Z(n628) );
  NAND2_X1 U699 ( .A1(G43), .A2(n802), .ZN(n626) );
  XNOR2_X1 U700 ( .A(KEYINPUT73), .B(n626), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n630), .A2(n629), .ZN(n993) );
  INV_X1 U703 ( .A(G1996), .ZN(n960) );
  NOR2_X1 U704 ( .A1(n667), .A2(n960), .ZN(n631) );
  XOR2_X1 U705 ( .A(n631), .B(KEYINPUT26), .Z(n633) );
  NAND2_X1 U706 ( .A1(n667), .A2(G1341), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U708 ( .A1(n993), .A2(n634), .ZN(n646) );
  NAND2_X1 U709 ( .A1(G66), .A2(n795), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G54), .A2(n802), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U712 ( .A1(G79), .A2(n794), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G92), .A2(n798), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n641), .B(KEYINPUT15), .ZN(n978) );
  NAND2_X1 U717 ( .A1(G1348), .A2(n667), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n642), .A2(G2067), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n647) );
  NOR2_X1 U720 ( .A1(n978), .A2(n647), .ZN(n645) );
  OR2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n978), .A2(n647), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  AND2_X1 U726 ( .A1(G171), .A2(n655), .ZN(n656) );
  XNOR2_X1 U727 ( .A(KEYINPUT99), .B(n658), .ZN(n672) );
  INV_X1 U728 ( .A(KEYINPUT100), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(n666) );
  INV_X1 U730 ( .A(n661), .ZN(n662) );
  AND2_X1 U731 ( .A1(G8), .A2(n662), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n685), .A2(G1971), .ZN(n669) );
  NOR2_X1 U734 ( .A1(G2090), .A2(n667), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U736 ( .A1(n670), .A2(G303), .ZN(n674) );
  AND2_X1 U737 ( .A1(n671), .A2(n674), .ZN(n673) );
  NAND2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n678) );
  INV_X1 U739 ( .A(n674), .ZN(n675) );
  OR2_X1 U740 ( .A1(n675), .A2(G286), .ZN(n676) );
  AND2_X1 U741 ( .A1(n676), .A2(G8), .ZN(n677) );
  NAND2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U743 ( .A(n679), .B(KEYINPUT32), .Z(n680) );
  NOR2_X2 U744 ( .A1(n681), .A2(n680), .ZN(n745) );
  NAND2_X1 U745 ( .A1(G8), .A2(G166), .ZN(n682) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XOR2_X1 U747 ( .A(KEYINPUT101), .B(n683), .Z(n684) );
  NOR2_X1 U748 ( .A1(n745), .A2(n684), .ZN(n686) );
  INV_X1 U749 ( .A(n685), .ZN(n754) );
  OR2_X1 U750 ( .A1(n686), .A2(n754), .ZN(n691) );
  NOR2_X1 U751 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XOR2_X1 U752 ( .A(n687), .B(KEYINPUT24), .Z(n688) );
  XNOR2_X1 U753 ( .A(KEYINPUT95), .B(n688), .ZN(n689) );
  NAND2_X1 U754 ( .A1(n689), .A2(n754), .ZN(n690) );
  NAND2_X1 U755 ( .A1(n691), .A2(n690), .ZN(n728) );
  NOR2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n729) );
  XOR2_X1 U757 ( .A(n729), .B(KEYINPUT91), .Z(n711) );
  NAND2_X1 U758 ( .A1(G119), .A2(n894), .ZN(n695) );
  NAND2_X1 U759 ( .A1(G107), .A2(n895), .ZN(n694) );
  NAND2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U761 ( .A1(G131), .A2(n890), .ZN(n696) );
  XNOR2_X1 U762 ( .A(KEYINPUT89), .B(n696), .ZN(n697) );
  NOR2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U764 ( .A1(G95), .A2(n891), .ZN(n699) );
  NAND2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n886) );
  NAND2_X1 U766 ( .A1(G1991), .A2(n886), .ZN(n701) );
  XNOR2_X1 U767 ( .A(n701), .B(KEYINPUT90), .ZN(n710) );
  NAND2_X1 U768 ( .A1(G129), .A2(n894), .ZN(n703) );
  NAND2_X1 U769 ( .A1(G117), .A2(n895), .ZN(n702) );
  NAND2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U771 ( .A1(n891), .A2(G105), .ZN(n704) );
  XOR2_X1 U772 ( .A(KEYINPUT38), .B(n704), .Z(n705) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U774 ( .A1(n890), .A2(G141), .ZN(n707) );
  NAND2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n885) );
  NAND2_X1 U776 ( .A1(G1996), .A2(n885), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n941) );
  AND2_X1 U778 ( .A1(n711), .A2(n941), .ZN(n734) );
  XOR2_X1 U779 ( .A(KEYINPUT92), .B(n734), .Z(n723) );
  NAND2_X1 U780 ( .A1(G140), .A2(n890), .ZN(n713) );
  NAND2_X1 U781 ( .A1(G104), .A2(n891), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U783 ( .A(KEYINPUT34), .B(n714), .ZN(n720) );
  NAND2_X1 U784 ( .A1(n895), .A2(G116), .ZN(n715) );
  XOR2_X1 U785 ( .A(KEYINPUT87), .B(n715), .Z(n717) );
  NAND2_X1 U786 ( .A1(n894), .A2(G128), .ZN(n716) );
  NAND2_X1 U787 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U788 ( .A(KEYINPUT35), .B(n718), .Z(n719) );
  NOR2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U790 ( .A(KEYINPUT36), .B(n721), .Z(n904) );
  XOR2_X1 U791 ( .A(G2067), .B(KEYINPUT37), .Z(n730) );
  AND2_X1 U792 ( .A1(n904), .A2(n730), .ZN(n946) );
  NAND2_X1 U793 ( .A1(n946), .A2(n729), .ZN(n722) );
  XNOR2_X1 U794 ( .A(n722), .B(KEYINPUT88), .ZN(n731) );
  NAND2_X1 U795 ( .A1(n723), .A2(n731), .ZN(n724) );
  XNOR2_X1 U796 ( .A(KEYINPUT93), .B(n724), .ZN(n727) );
  XNOR2_X1 U797 ( .A(G1986), .B(G290), .ZN(n989) );
  NAND2_X1 U798 ( .A1(n729), .A2(n989), .ZN(n725) );
  XNOR2_X1 U799 ( .A(n725), .B(KEYINPUT86), .ZN(n726) );
  AND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n756) );
  NAND2_X1 U801 ( .A1(n728), .A2(n756), .ZN(n744) );
  INV_X1 U802 ( .A(n729), .ZN(n741) );
  NOR2_X1 U803 ( .A1(n904), .A2(n730), .ZN(n942) );
  INV_X1 U804 ( .A(n731), .ZN(n738) );
  NOR2_X1 U805 ( .A1(G1996), .A2(n885), .ZN(n929) );
  NOR2_X1 U806 ( .A1(G1986), .A2(G290), .ZN(n732) );
  NOR2_X1 U807 ( .A1(G1991), .A2(n886), .ZN(n934) );
  NOR2_X1 U808 ( .A1(n732), .A2(n934), .ZN(n733) );
  NOR2_X1 U809 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U810 ( .A1(n929), .A2(n735), .ZN(n736) );
  XOR2_X1 U811 ( .A(KEYINPUT39), .B(n736), .Z(n737) );
  NOR2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U813 ( .A1(n942), .A2(n739), .ZN(n740) );
  NOR2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U815 ( .A(n742), .B(KEYINPUT102), .Z(n743) );
  AND2_X1 U816 ( .A1(n744), .A2(n743), .ZN(n761) );
  XNOR2_X1 U817 ( .A(G1981), .B(G305), .ZN(n975) );
  INV_X1 U818 ( .A(n745), .ZN(n749) );
  NOR2_X1 U819 ( .A1(G1976), .A2(G288), .ZN(n982) );
  NOR2_X1 U820 ( .A1(G1971), .A2(G303), .ZN(n985) );
  NOR2_X1 U821 ( .A1(n982), .A2(n985), .ZN(n747) );
  INV_X1 U822 ( .A(KEYINPUT33), .ZN(n746) );
  AND2_X1 U823 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U824 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n987) );
  AND2_X1 U826 ( .A1(n987), .A2(n754), .ZN(n750) );
  OR2_X1 U827 ( .A1(KEYINPUT33), .A2(n750), .ZN(n751) );
  NAND2_X1 U828 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U829 ( .A1(n975), .A2(n753), .ZN(n759) );
  AND2_X1 U830 ( .A1(n982), .A2(KEYINPUT33), .ZN(n755) );
  NAND2_X1 U831 ( .A1(n755), .A2(n754), .ZN(n757) );
  AND2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U833 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U834 ( .A1(n761), .A2(n760), .ZN(n764) );
  INV_X1 U835 ( .A(KEYINPUT40), .ZN(n762) );
  XNOR2_X1 U836 ( .A(n764), .B(n763), .ZN(G329) );
  INV_X1 U837 ( .A(G57), .ZN(G237) );
  INV_X1 U838 ( .A(G132), .ZN(G219) );
  NAND2_X1 U839 ( .A1(G94), .A2(G452), .ZN(n766) );
  XNOR2_X1 U840 ( .A(n766), .B(KEYINPUT69), .ZN(G173) );
  XOR2_X1 U841 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n768) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U843 ( .A(n768), .B(n767), .ZN(G223) );
  INV_X1 U844 ( .A(G223), .ZN(n831) );
  NAND2_X1 U845 ( .A1(n831), .A2(G567), .ZN(n769) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n769), .Z(G234) );
  INV_X1 U847 ( .A(G860), .ZN(n793) );
  NOR2_X1 U848 ( .A1(n993), .A2(n793), .ZN(n770) );
  XOR2_X1 U849 ( .A(KEYINPUT74), .B(n770), .Z(G153) );
  INV_X1 U850 ( .A(G171), .ZN(G301) );
  NAND2_X1 U851 ( .A1(G868), .A2(G301), .ZN(n772) );
  INV_X1 U852 ( .A(G868), .ZN(n813) );
  NAND2_X1 U853 ( .A1(n978), .A2(n813), .ZN(n771) );
  NAND2_X1 U854 ( .A1(n772), .A2(n771), .ZN(G284) );
  INV_X1 U855 ( .A(n979), .ZN(G299) );
  NOR2_X1 U856 ( .A1(G286), .A2(n813), .ZN(n774) );
  NOR2_X1 U857 ( .A1(G868), .A2(G299), .ZN(n773) );
  NOR2_X1 U858 ( .A1(n774), .A2(n773), .ZN(G297) );
  NAND2_X1 U859 ( .A1(n793), .A2(G559), .ZN(n775) );
  INV_X1 U860 ( .A(n978), .ZN(n791) );
  NAND2_X1 U861 ( .A1(n775), .A2(n791), .ZN(n776) );
  XNOR2_X1 U862 ( .A(n776), .B(KEYINPUT16), .ZN(n777) );
  XNOR2_X1 U863 ( .A(KEYINPUT76), .B(n777), .ZN(G148) );
  NOR2_X1 U864 ( .A1(n978), .A2(n813), .ZN(n778) );
  XNOR2_X1 U865 ( .A(n778), .B(KEYINPUT77), .ZN(n779) );
  NOR2_X1 U866 ( .A1(G559), .A2(n779), .ZN(n781) );
  NOR2_X1 U867 ( .A1(G868), .A2(n993), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(G282) );
  NAND2_X1 U869 ( .A1(n894), .A2(G123), .ZN(n782) );
  XNOR2_X1 U870 ( .A(n782), .B(KEYINPUT18), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G111), .A2(n895), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U873 ( .A1(G135), .A2(n890), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G99), .A2(n891), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n933) );
  XOR2_X1 U877 ( .A(G2096), .B(n933), .Z(n789) );
  NOR2_X1 U878 ( .A1(G2100), .A2(n789), .ZN(n790) );
  XOR2_X1 U879 ( .A(KEYINPUT78), .B(n790), .Z(G156) );
  NAND2_X1 U880 ( .A1(G559), .A2(n791), .ZN(n792) );
  XOR2_X1 U881 ( .A(n993), .B(n792), .Z(n811) );
  NAND2_X1 U882 ( .A1(n793), .A2(n811), .ZN(n805) );
  NAND2_X1 U883 ( .A1(G80), .A2(n794), .ZN(n797) );
  NAND2_X1 U884 ( .A1(G67), .A2(n795), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U886 ( .A1(G93), .A2(n798), .ZN(n799) );
  XNOR2_X1 U887 ( .A(KEYINPUT79), .B(n799), .ZN(n800) );
  NOR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U889 ( .A1(n802), .A2(G55), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n814) );
  XNOR2_X1 U891 ( .A(n805), .B(n814), .ZN(G145) );
  XNOR2_X1 U892 ( .A(G288), .B(KEYINPUT19), .ZN(n807) );
  XNOR2_X1 U893 ( .A(n979), .B(G166), .ZN(n806) );
  XNOR2_X1 U894 ( .A(n807), .B(n806), .ZN(n808) );
  XNOR2_X1 U895 ( .A(n808), .B(G290), .ZN(n809) );
  XNOR2_X1 U896 ( .A(n809), .B(n814), .ZN(n810) );
  XNOR2_X1 U897 ( .A(n810), .B(G305), .ZN(n859) );
  XNOR2_X1 U898 ( .A(n811), .B(n859), .ZN(n812) );
  NAND2_X1 U899 ( .A1(n812), .A2(G868), .ZN(n816) );
  NAND2_X1 U900 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n816), .A2(n815), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2084), .A2(G2078), .ZN(n818) );
  XOR2_X1 U903 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n817) );
  XNOR2_X1 U904 ( .A(n818), .B(n817), .ZN(n819) );
  NAND2_X1 U905 ( .A1(G2090), .A2(n819), .ZN(n820) );
  XNOR2_X1 U906 ( .A(KEYINPUT21), .B(n820), .ZN(n821) );
  NAND2_X1 U907 ( .A1(n821), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U908 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U909 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U910 ( .A1(G220), .A2(G219), .ZN(n822) );
  XOR2_X1 U911 ( .A(KEYINPUT22), .B(n822), .Z(n823) );
  NOR2_X1 U912 ( .A1(G218), .A2(n823), .ZN(n824) );
  NAND2_X1 U913 ( .A1(G96), .A2(n824), .ZN(n836) );
  NAND2_X1 U914 ( .A1(n836), .A2(G2106), .ZN(n828) );
  NAND2_X1 U915 ( .A1(G69), .A2(G120), .ZN(n825) );
  NOR2_X1 U916 ( .A1(G237), .A2(n825), .ZN(n826) );
  NAND2_X1 U917 ( .A1(G108), .A2(n826), .ZN(n837) );
  NAND2_X1 U918 ( .A1(n837), .A2(G567), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(n838) );
  NAND2_X1 U920 ( .A1(G483), .A2(G661), .ZN(n829) );
  NOR2_X1 U921 ( .A1(n838), .A2(n829), .ZN(n830) );
  XOR2_X1 U922 ( .A(KEYINPUT83), .B(n830), .Z(n835) );
  NAND2_X1 U923 ( .A1(n835), .A2(G36), .ZN(G176) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n831), .ZN(G217) );
  NAND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n832) );
  XOR2_X1 U926 ( .A(KEYINPUT104), .B(n832), .Z(n833) );
  NAND2_X1 U927 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  INV_X1 U936 ( .A(n838), .ZN(G319) );
  XOR2_X1 U937 ( .A(KEYINPUT105), .B(G2678), .Z(n840) );
  XNOR2_X1 U938 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2090), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2096), .B(G2100), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n848) );
  XOR2_X1 U946 ( .A(G2084), .B(G2078), .Z(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1976), .B(G1956), .Z(n850) );
  XNOR2_X1 U949 ( .A(G1966), .B(G1961), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U951 ( .A(G1991), .B(G1986), .Z(n852) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1971), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U954 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U955 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U957 ( .A(G1981), .B(G2474), .Z(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(G229) );
  XNOR2_X1 U959 ( .A(n859), .B(KEYINPUT113), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n978), .B(G286), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n993), .B(G171), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n864) );
  NOR2_X1 U964 ( .A1(G37), .A2(n864), .ZN(G397) );
  NAND2_X1 U965 ( .A1(G100), .A2(n891), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n865), .B(KEYINPUT108), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G112), .A2(n895), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n868), .B(KEYINPUT109), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G136), .A2(n890), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n894), .A2(G124), .ZN(n871) );
  XOR2_X1 U973 ( .A(KEYINPUT44), .B(n871), .Z(n872) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(G162) );
  XOR2_X1 U975 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n875) );
  XNOR2_X1 U976 ( .A(n933), .B(KEYINPUT111), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n884) );
  NAND2_X1 U978 ( .A1(G130), .A2(n894), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G118), .A2(n895), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G142), .A2(n890), .ZN(n879) );
  NAND2_X1 U982 ( .A1(G106), .A2(n891), .ZN(n878) );
  NAND2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U984 ( .A(n880), .B(KEYINPUT45), .Z(n881) );
  NOR2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U986 ( .A(n884), .B(n883), .Z(n889) );
  XNOR2_X1 U987 ( .A(G160), .B(n885), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U989 ( .A(n889), .B(n888), .Z(n903) );
  NAND2_X1 U990 ( .A1(G139), .A2(n890), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G103), .A2(n891), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n900) );
  NAND2_X1 U993 ( .A1(G127), .A2(n894), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G115), .A2(n895), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(KEYINPUT110), .B(n901), .Z(n924) );
  XNOR2_X1 U999 ( .A(G164), .B(n924), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(G162), .B(n904), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(KEYINPUT112), .B(n908), .ZN(G395) );
  XOR2_X1 U1005 ( .A(G2451), .B(G2430), .Z(n910) );
  XNOR2_X1 U1006 ( .A(G2438), .B(G2443), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n916) );
  XOR2_X1 U1008 ( .A(G2435), .B(G2454), .Z(n912) );
  XNOR2_X1 U1009 ( .A(G1341), .B(G1348), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n914) );
  XOR2_X1 U1011 ( .A(G2446), .B(G2427), .Z(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1013 ( .A(n916), .B(n915), .Z(n917) );
  NAND2_X1 U1014 ( .A1(G14), .A2(n917), .ZN(n923) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n923), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1019 ( .A1(G397), .A2(G395), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  INV_X1 U1023 ( .A(n923), .ZN(G401) );
  INV_X1 U1024 ( .A(KEYINPUT55), .ZN(n950) );
  XNOR2_X1 U1025 ( .A(KEYINPUT116), .B(KEYINPUT52), .ZN(n948) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n926) );
  XNOR2_X1 U1027 ( .A(G2072), .B(n924), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1029 ( .A(KEYINPUT50), .B(n927), .ZN(n932) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n930), .Z(n931) );
  NAND2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1035 ( .A(KEYINPUT114), .B(n935), .Z(n937) );
  XOR2_X1 U1036 ( .A(G160), .B(G2084), .Z(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n938), .B(KEYINPUT115), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n948), .B(n947), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1045 ( .A1(n951), .A2(G29), .ZN(n1037) );
  XNOR2_X1 U1046 ( .A(G27), .B(n952), .ZN(n965) );
  XNOR2_X1 U1047 ( .A(KEYINPUT117), .B(G2067), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(n953), .B(G26), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(G33), .B(n954), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n955), .A2(G28), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G25), .B(G1991), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n963) );
  XOR2_X1 U1054 ( .A(KEYINPUT118), .B(n960), .Z(n961) );
  XNOR2_X1 U1055 ( .A(G32), .B(n961), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n966), .B(KEYINPUT53), .ZN(n969) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n967) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n967), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(G35), .B(G2090), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1064 ( .A(KEYINPUT55), .B(n972), .Z(n973) );
  NOR2_X1 U1065 ( .A1(G29), .A2(n973), .ZN(n1033) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n1004) );
  XOR2_X1 U1067 ( .A(G1966), .B(G168), .Z(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1069 ( .A(KEYINPUT57), .B(n976), .Z(n1002) );
  XOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT119), .Z(n977) );
  XNOR2_X1 U1071 ( .A(n978), .B(n977), .ZN(n999) );
  XNOR2_X1 U1072 ( .A(n979), .B(G1956), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(G1971), .A2(G303), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT120), .B(n982), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n991) );
  INV_X1 U1077 ( .A(n985), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(KEYINPUT121), .B(n992), .ZN(n997) );
  XNOR2_X1 U1082 ( .A(G301), .B(G1961), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(n993), .B(G1341), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(KEYINPUT122), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1031) );
  INV_X1 U1090 ( .A(G16), .ZN(n1029) );
  XNOR2_X1 U1091 ( .A(n1005), .B(G5), .ZN(n1025) );
  XNOR2_X1 U1092 ( .A(G1348), .B(KEYINPUT59), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(n1006), .B(G4), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G20), .B(G1956), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1013), .Z(n1015) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G21), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT123), .B(n1016), .ZN(n1023) );
  XNOR2_X1 U1104 ( .A(G1971), .B(G22), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(G23), .B(G1976), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1107 ( .A(G1986), .B(G24), .Z(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1112 ( .A(n1026), .B(KEYINPUT61), .ZN(n1027) );
  XOR2_X1 U1113 ( .A(KEYINPUT124), .B(n1027), .Z(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1117 ( .A1(G11), .A2(n1034), .ZN(n1035) );
  XNOR2_X1 U1118 ( .A(KEYINPUT125), .B(n1035), .ZN(n1036) );
  NAND2_X1 U1119 ( .A1(n1037), .A2(n1036), .ZN(n1039) );
  XOR2_X1 U1120 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1038) );
  XNOR2_X1 U1121 ( .A(n1039), .B(n1038), .ZN(G311) );
  XNOR2_X1 U1122 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

