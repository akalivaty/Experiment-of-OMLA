

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777;

  NOR2_X2 U373 ( .A1(n654), .A2(n777), .ZN(n607) );
  XNOR2_X1 U374 ( .A(n561), .B(n560), .ZN(n585) );
  NOR2_X1 U375 ( .A1(n645), .A2(n750), .ZN(n647) );
  OR2_X2 U376 ( .A1(n373), .A2(n372), .ZN(n742) );
  NOR2_X2 U377 ( .A1(n662), .A2(n402), .ZN(n623) );
  XNOR2_X2 U378 ( .A(n356), .B(KEYINPUT121), .ZN(n355) );
  AND2_X2 U379 ( .A1(n737), .A2(n736), .ZN(n356) );
  XNOR2_X2 U380 ( .A(n763), .B(G146), .ZN(n454) );
  NOR2_X2 U381 ( .A1(n537), .A2(n541), .ZN(n538) );
  NOR2_X2 U382 ( .A1(n616), .A2(n703), .ZN(n617) );
  XNOR2_X1 U383 ( .A(n637), .B(n636), .ZN(n732) );
  NAND2_X1 U384 ( .A1(n397), .A2(n393), .ZN(n662) );
  INV_X1 U385 ( .A(n611), .ZN(n353) );
  NOR2_X1 U386 ( .A1(n525), .A2(n524), .ZN(n686) );
  AND2_X1 U387 ( .A1(n409), .A2(n406), .ZN(n405) );
  OR2_X1 U388 ( .A1(n615), .A2(n614), .ZN(n703) );
  XNOR2_X1 U389 ( .A(n521), .B(n520), .ZN(n536) );
  XNOR2_X1 U390 ( .A(n449), .B(n450), .ZN(n519) );
  XNOR2_X1 U391 ( .A(n513), .B(n425), .ZN(n764) );
  XNOR2_X1 U392 ( .A(n426), .B(G146), .ZN(n513) );
  XNOR2_X1 U393 ( .A(n512), .B(n443), .ZN(n499) );
  INV_X1 U394 ( .A(KEYINPUT68), .ZN(n385) );
  NAND2_X1 U395 ( .A1(n354), .A2(n364), .ZN(n747) );
  NOR2_X1 U396 ( .A1(n371), .A2(n638), .ZN(n354) );
  XNOR2_X2 U397 ( .A(n635), .B(KEYINPUT65), .ZN(n639) );
  XNOR2_X1 U398 ( .A(n459), .B(G140), .ZN(n425) );
  NOR2_X1 U399 ( .A1(n712), .A2(n407), .ZN(n406) );
  NAND2_X1 U400 ( .A1(n408), .A2(n411), .ZN(n407) );
  XNOR2_X1 U401 ( .A(n472), .B(n471), .ZN(n545) );
  XNOR2_X1 U402 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U403 ( .A1(n748), .A2(G902), .ZN(n472) );
  INV_X1 U404 ( .A(n592), .ZN(n610) );
  NAND2_X1 U405 ( .A1(n610), .A2(n401), .ZN(n400) );
  INV_X1 U406 ( .A(G134), .ZN(n443) );
  AND2_X1 U407 ( .A1(n630), .A2(n629), .ZN(n634) );
  XNOR2_X1 U408 ( .A(G113), .B(KEYINPUT3), .ZN(n447) );
  XNOR2_X1 U409 ( .A(n382), .B(n381), .ZN(n477) );
  INV_X1 U410 ( .A(KEYINPUT90), .ZN(n381) );
  INV_X1 U411 ( .A(G234), .ZN(n413) );
  XNOR2_X1 U412 ( .A(n418), .B(n499), .ZN(n763) );
  XNOR2_X1 U413 ( .A(n481), .B(n442), .ZN(n418) );
  XNOR2_X1 U414 ( .A(KEYINPUT4), .B(G137), .ZN(n442) );
  OR2_X1 U415 ( .A1(G237), .A2(G902), .ZN(n522) );
  NAND2_X1 U416 ( .A1(n544), .A2(n543), .ZN(n712) );
  INV_X1 U417 ( .A(G902), .ZN(n501) );
  XNOR2_X1 U418 ( .A(n489), .B(n488), .ZN(n648) );
  XNOR2_X1 U419 ( .A(n437), .B(G107), .ZN(n517) );
  XNOR2_X1 U420 ( .A(G104), .B(G110), .ZN(n437) );
  XNOR2_X1 U421 ( .A(G101), .B(G140), .ZN(n388) );
  INV_X1 U422 ( .A(KEYINPUT77), .ZN(n438) );
  XNOR2_X1 U423 ( .A(n432), .B(n519), .ZN(n757) );
  XNOR2_X1 U424 ( .A(n517), .B(n518), .ZN(n432) );
  XNOR2_X1 U425 ( .A(n391), .B(n390), .ZN(n518) );
  INV_X1 U426 ( .A(KEYINPUT16), .ZN(n390) );
  AND2_X1 U427 ( .A1(n694), .A2(n693), .ZN(n422) );
  INV_X1 U428 ( .A(KEYINPUT106), .ZN(n424) );
  XNOR2_X1 U429 ( .A(n433), .B(n587), .ZN(n596) );
  XNOR2_X1 U430 ( .A(n586), .B(KEYINPUT74), .ZN(n587) );
  INV_X1 U431 ( .A(KEYINPUT22), .ZN(n586) );
  NAND2_X1 U432 ( .A1(n596), .A2(n614), .ZN(n611) );
  BUF_X1 U433 ( .A(n545), .Z(n696) );
  NOR2_X1 U434 ( .A1(n610), .A2(n401), .ZN(n399) );
  NAND2_X1 U435 ( .A1(n353), .A2(n400), .ZN(n394) );
  AND2_X1 U436 ( .A1(n396), .A2(n612), .ZN(n395) );
  INV_X1 U437 ( .A(G953), .ZN(n758) );
  XNOR2_X1 U438 ( .A(n416), .B(n415), .ZN(n748) );
  XNOR2_X1 U439 ( .A(n465), .B(n463), .ZN(n415) );
  XNOR2_X1 U440 ( .A(n464), .B(n417), .ZN(n416) );
  XNOR2_X1 U441 ( .A(n497), .B(n389), .ZN(n500) );
  XNOR2_X1 U442 ( .A(n496), .B(n498), .ZN(n389) );
  INV_X1 U443 ( .A(G478), .ZN(n370) );
  INV_X1 U444 ( .A(G475), .ZN(n369) );
  XNOR2_X1 U445 ( .A(n757), .B(n430), .ZN(n657) );
  XNOR2_X1 U446 ( .A(n431), .B(n514), .ZN(n430) );
  XNOR2_X1 U447 ( .A(n513), .B(n435), .ZN(n514) );
  XNOR2_X1 U448 ( .A(n515), .B(n516), .ZN(n431) );
  INV_X1 U449 ( .A(G210), .ZN(n368) );
  INV_X1 U450 ( .A(KEYINPUT15), .ZN(n466) );
  NAND2_X1 U451 ( .A1(G234), .A2(G237), .ZN(n475) );
  NOR2_X1 U452 ( .A1(n700), .A2(n383), .ZN(n701) );
  NOR2_X1 U453 ( .A1(G953), .A2(G237), .ZN(n486) );
  XNOR2_X1 U454 ( .A(G143), .B(G104), .ZN(n482) );
  XNOR2_X1 U455 ( .A(G113), .B(G122), .ZN(n480) );
  XNOR2_X1 U456 ( .A(G119), .B(G116), .ZN(n448) );
  XNOR2_X1 U457 ( .A(KEYINPUT75), .B(G122), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n577), .B(n374), .ZN(n541) );
  INV_X1 U459 ( .A(KEYINPUT38), .ZN(n374) );
  XNOR2_X1 U460 ( .A(n589), .B(n420), .ZN(n592) );
  INV_X1 U461 ( .A(KEYINPUT6), .ZN(n420) );
  NAND2_X1 U462 ( .A1(n584), .A2(KEYINPUT0), .ZN(n411) );
  NAND2_X1 U463 ( .A1(n403), .A2(n357), .ZN(n410) );
  AND2_X1 U464 ( .A1(n378), .A2(n377), .ZN(n478) );
  INV_X1 U465 ( .A(G900), .ZN(n377) );
  XNOR2_X1 U466 ( .A(n581), .B(KEYINPUT101), .ZN(n378) );
  INV_X1 U467 ( .A(n709), .ZN(n419) );
  INV_X1 U468 ( .A(KEYINPUT30), .ZN(n379) );
  NOR2_X1 U469 ( .A1(n545), .A2(n697), .ZN(n613) );
  XNOR2_X1 U470 ( .A(n764), .B(n434), .ZN(n464) );
  XOR2_X1 U471 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n461) );
  XNOR2_X1 U472 ( .A(G119), .B(G128), .ZN(n457) );
  XOR2_X1 U473 ( .A(G110), .B(G137), .Z(n458) );
  XNOR2_X1 U474 ( .A(n414), .B(n412), .ZN(n462) );
  XNOR2_X1 U475 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n414) );
  NOR2_X1 U476 ( .A1(n413), .A2(G953), .ZN(n412) );
  XNOR2_X1 U477 ( .A(G116), .B(G107), .ZN(n494) );
  INV_X1 U478 ( .A(G125), .ZN(n426) );
  BUF_X1 U479 ( .A(n536), .Z(n577) );
  XNOR2_X1 U480 ( .A(n376), .B(KEYINPUT41), .ZN(n707) );
  NOR2_X1 U481 ( .A1(n714), .A2(n712), .ZN(n376) );
  INV_X1 U482 ( .A(KEYINPUT34), .ZN(n386) );
  XNOR2_X1 U483 ( .A(n423), .B(KEYINPUT78), .ZN(n677) );
  NOR2_X1 U484 ( .A1(n562), .A2(n585), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n492), .B(n491), .ZN(n542) );
  XNOR2_X1 U486 ( .A(n504), .B(n503), .ZN(n544) );
  BUF_X1 U487 ( .A(n421), .Z(n383) );
  NAND2_X1 U488 ( .A1(n366), .A2(n365), .ZN(n643) );
  NOR2_X1 U489 ( .A1(n638), .A2(n367), .ZN(n365) );
  INV_X1 U490 ( .A(G472), .ZN(n367) );
  INV_X1 U491 ( .A(G469), .ZN(n372) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n444) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n517), .B(n388), .ZN(n441) );
  BUF_X1 U495 ( .A(n677), .Z(n384) );
  INV_X1 U496 ( .A(KEYINPUT100), .ZN(n588) );
  NAND2_X1 U497 ( .A1(n353), .A2(n398), .ZN(n397) );
  NAND2_X1 U498 ( .A1(n394), .A2(n395), .ZN(n393) );
  AND2_X1 U499 ( .A1(n399), .A2(n612), .ZN(n398) );
  INV_X1 U500 ( .A(G217), .ZN(n371) );
  NAND2_X1 U501 ( .A1(n364), .A2(n363), .ZN(n744) );
  NOR2_X1 U502 ( .A1(n638), .A2(n370), .ZN(n363) );
  NOR2_X1 U503 ( .A1(n652), .A2(n750), .ZN(n653) );
  NOR2_X1 U504 ( .A1(n660), .A2(n750), .ZN(n661) );
  NOR2_X1 U505 ( .A1(n584), .A2(KEYINPUT0), .ZN(n357) );
  XOR2_X1 U506 ( .A(n455), .B(G472), .Z(n358) );
  INV_X1 U507 ( .A(KEYINPUT86), .ZN(n401) );
  XOR2_X1 U508 ( .A(n650), .B(n649), .Z(n359) );
  INV_X1 U509 ( .A(n639), .ZN(n366) );
  NAND2_X1 U510 ( .A1(n360), .A2(n364), .ZN(n651) );
  NOR2_X1 U511 ( .A1(n638), .A2(n369), .ZN(n360) );
  NAND2_X1 U512 ( .A1(n364), .A2(n361), .ZN(n373) );
  INV_X1 U513 ( .A(n638), .ZN(n361) );
  INV_X2 U514 ( .A(n639), .ZN(n364) );
  NAND2_X1 U515 ( .A1(n362), .A2(n366), .ZN(n659) );
  NOR2_X1 U516 ( .A1(n638), .A2(n368), .ZN(n362) );
  NOR2_X1 U517 ( .A1(n612), .A2(n547), .ZN(n549) );
  XNOR2_X1 U518 ( .A(n380), .B(n379), .ZN(n526) );
  XNOR2_X1 U519 ( .A(n387), .B(n386), .ZN(n601) );
  NAND2_X1 U520 ( .A1(n585), .A2(KEYINPUT0), .ZN(n409) );
  XNOR2_X2 U521 ( .A(n375), .B(KEYINPUT33), .ZN(n719) );
  NAND2_X1 U522 ( .A1(n422), .A2(n610), .ZN(n375) );
  NOR2_X1 U523 ( .A1(n574), .A2(n561), .ZN(n523) );
  XNOR2_X1 U524 ( .A(n686), .B(KEYINPUT85), .ZN(n533) );
  NOR2_X1 U525 ( .A1(n589), .A2(n419), .ZN(n380) );
  NAND2_X1 U526 ( .A1(n476), .A2(G902), .ZN(n382) );
  XNOR2_X2 U527 ( .A(n385), .B(G131), .ZN(n481) );
  NAND2_X1 U528 ( .A1(n719), .A2(n620), .ZN(n387) );
  AND2_X1 U529 ( .A1(n392), .A2(n621), .ZN(n402) );
  NAND2_X1 U530 ( .A1(n683), .A2(n665), .ZN(n392) );
  XNOR2_X1 U531 ( .A(n617), .B(KEYINPUT31), .ZN(n683) );
  NAND2_X1 U532 ( .A1(n400), .A2(KEYINPUT86), .ZN(n396) );
  NAND2_X1 U533 ( .A1(n404), .A2(n410), .ZN(n616) );
  INV_X1 U534 ( .A(n585), .ZN(n403) );
  AND2_X1 U535 ( .A1(n409), .A2(n411), .ZN(n404) );
  NAND2_X1 U536 ( .A1(n405), .A2(n410), .ZN(n433) );
  INV_X1 U537 ( .A(n697), .ZN(n408) );
  NAND2_X1 U538 ( .A1(n493), .A2(G221), .ZN(n417) );
  XNOR2_X2 U539 ( .A(G143), .B(G128), .ZN(n512) );
  NAND2_X1 U540 ( .A1(n421), .A2(n546), .ZN(n547) );
  NOR2_X1 U541 ( .A1(n618), .A2(n383), .ZN(n619) );
  NAND2_X1 U542 ( .A1(n694), .A2(n421), .ZN(n615) );
  INV_X2 U543 ( .A(n589), .ZN(n421) );
  XNOR2_X2 U544 ( .A(n456), .B(n358), .ZN(n589) );
  INV_X1 U545 ( .A(n693), .ZN(n614) );
  NAND2_X1 U546 ( .A1(n677), .A2(n621), .ZN(n563) );
  XNOR2_X1 U547 ( .A(n553), .B(n424), .ZN(n562) );
  XNOR2_X2 U548 ( .A(n427), .B(KEYINPUT45), .ZN(n725) );
  NAND2_X1 U549 ( .A1(n428), .A2(n624), .ZN(n427) );
  XNOR2_X1 U550 ( .A(n429), .B(KEYINPUT87), .ZN(n428) );
  NAND2_X1 U551 ( .A1(n623), .A2(n622), .ZN(n429) );
  NAND2_X1 U552 ( .A1(n657), .A2(n628), .ZN(n521) );
  XNOR2_X2 U553 ( .A(n540), .B(n539), .ZN(n774) );
  OR2_X2 U554 ( .A1(n573), .A2(n679), .ZN(n540) );
  AND2_X2 U555 ( .A1(n625), .A2(n725), .ZN(n436) );
  XNOR2_X1 U556 ( .A(n764), .B(n487), .ZN(n488) );
  XOR2_X1 U557 ( .A(n461), .B(n460), .Z(n434) );
  AND2_X1 U558 ( .A1(G224), .A2(n758), .ZN(n435) );
  INV_X1 U559 ( .A(KEYINPUT10), .ZN(n459) );
  BUF_X1 U560 ( .A(n613), .Z(n694) );
  XNOR2_X1 U561 ( .A(n490), .B(G475), .ZN(n491) );
  INV_X1 U562 ( .A(KEYINPUT63), .ZN(n646) );
  NAND2_X1 U563 ( .A1(G227), .A2(n758), .ZN(n439) );
  XNOR2_X1 U564 ( .A(n454), .B(n444), .ZN(n739) );
  NAND2_X1 U565 ( .A1(n739), .A2(n501), .ZN(n446) );
  XOR2_X1 U566 ( .A(KEYINPUT71), .B(G469), .Z(n445) );
  XNOR2_X2 U567 ( .A(n446), .B(n445), .ZN(n550) );
  XNOR2_X2 U568 ( .A(n550), .B(KEYINPUT1), .ZN(n693) );
  XNOR2_X1 U569 ( .A(n693), .B(KEYINPUT88), .ZN(n594) );
  INV_X1 U570 ( .A(n594), .ZN(n525) );
  XNOR2_X1 U571 ( .A(n447), .B(G101), .ZN(n450) );
  XNOR2_X1 U572 ( .A(n448), .B(KEYINPUT72), .ZN(n449) );
  NAND2_X1 U573 ( .A1(n486), .A2(G210), .ZN(n451) );
  XNOR2_X1 U574 ( .A(n451), .B(KEYINPUT5), .ZN(n452) );
  XNOR2_X1 U575 ( .A(n519), .B(n452), .ZN(n453) );
  XNOR2_X1 U576 ( .A(n454), .B(n453), .ZN(n641) );
  OR2_X2 U577 ( .A1(n641), .A2(G902), .ZN(n456) );
  INV_X1 U578 ( .A(KEYINPUT73), .ZN(n455) );
  XNOR2_X1 U579 ( .A(n458), .B(n457), .ZN(n465) );
  XNOR2_X1 U580 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n460) );
  XNOR2_X1 U581 ( .A(KEYINPUT81), .B(n462), .ZN(n493) );
  XOR2_X1 U582 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n463) );
  XOR2_X1 U583 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n468) );
  XNOR2_X1 U584 ( .A(n466), .B(G902), .ZN(n631) );
  INV_X1 U585 ( .A(n631), .ZN(n628) );
  NAND2_X1 U586 ( .A1(G234), .A2(n628), .ZN(n467) );
  XNOR2_X1 U587 ( .A(n468), .B(n467), .ZN(n473) );
  NAND2_X1 U588 ( .A1(G217), .A2(n473), .ZN(n470) );
  INV_X1 U589 ( .A(KEYINPUT25), .ZN(n469) );
  NAND2_X1 U590 ( .A1(n473), .A2(G221), .ZN(n474) );
  XNOR2_X1 U591 ( .A(n474), .B(KEYINPUT21), .ZN(n697) );
  XNOR2_X1 U592 ( .A(n475), .B(KEYINPUT14), .ZN(n476) );
  NAND2_X1 U593 ( .A1(G952), .A2(n476), .ZN(n724) );
  NOR2_X1 U594 ( .A1(G953), .A2(n724), .ZN(n583) );
  NAND2_X1 U595 ( .A1(G953), .A2(n477), .ZN(n581) );
  NOR2_X1 U596 ( .A1(n583), .A2(n478), .ZN(n527) );
  NOR2_X1 U597 ( .A1(n697), .A2(n527), .ZN(n479) );
  XNOR2_X1 U598 ( .A(KEYINPUT70), .B(n479), .ZN(n546) );
  NAND2_X1 U599 ( .A1(n696), .A2(n546), .ZN(n505) );
  XNOR2_X1 U600 ( .A(n481), .B(n480), .ZN(n485) );
  XOR2_X1 U601 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n483) );
  XNOR2_X1 U602 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U603 ( .A(n485), .B(n484), .Z(n489) );
  NAND2_X1 U604 ( .A1(G214), .A2(n486), .ZN(n487) );
  NOR2_X1 U605 ( .A1(G902), .A2(n648), .ZN(n492) );
  XNOR2_X1 U606 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n490) );
  XNOR2_X1 U607 ( .A(KEYINPUT9), .B(KEYINPUT97), .ZN(n498) );
  NAND2_X1 U608 ( .A1(n493), .A2(G217), .ZN(n497) );
  XOR2_X1 U609 ( .A(KEYINPUT7), .B(G122), .Z(n495) );
  XNOR2_X1 U610 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U611 ( .A(n499), .B(n500), .ZN(n745) );
  NAND2_X1 U612 ( .A1(n745), .A2(n501), .ZN(n504) );
  XNOR2_X1 U613 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n502) );
  XNOR2_X1 U614 ( .A(n502), .B(G478), .ZN(n503) );
  NAND2_X1 U615 ( .A1(n542), .A2(n544), .ZN(n679) );
  NOR2_X1 U616 ( .A1(n505), .A2(n679), .ZN(n506) );
  NAND2_X1 U617 ( .A1(n610), .A2(n506), .ZN(n574) );
  INV_X1 U618 ( .A(KEYINPUT18), .ZN(n507) );
  NAND2_X1 U619 ( .A1(KEYINPUT89), .A2(n507), .ZN(n510) );
  INV_X1 U620 ( .A(KEYINPUT89), .ZN(n508) );
  NAND2_X1 U621 ( .A1(n508), .A2(KEYINPUT18), .ZN(n509) );
  NAND2_X1 U622 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U623 ( .A(n512), .B(n511), .ZN(n515) );
  XOR2_X1 U624 ( .A(KEYINPUT4), .B(KEYINPUT17), .Z(n516) );
  NAND2_X1 U625 ( .A1(n522), .A2(G210), .ZN(n520) );
  INV_X1 U626 ( .A(n536), .ZN(n532) );
  NAND2_X1 U627 ( .A1(G214), .A2(n522), .ZN(n709) );
  NAND2_X1 U628 ( .A1(n532), .A2(n709), .ZN(n561) );
  XOR2_X1 U629 ( .A(KEYINPUT36), .B(n523), .Z(n524) );
  NAND2_X1 U630 ( .A1(n550), .A2(n613), .ZN(n618) );
  XNOR2_X1 U631 ( .A(n618), .B(KEYINPUT103), .ZN(n529) );
  NOR2_X1 U632 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U633 ( .A1(n529), .A2(n528), .ZN(n537) );
  INV_X1 U634 ( .A(n544), .ZN(n530) );
  NAND2_X1 U635 ( .A1(n542), .A2(n530), .ZN(n599) );
  NOR2_X1 U636 ( .A1(n537), .A2(n599), .ZN(n531) );
  NAND2_X1 U637 ( .A1(n532), .A2(n531), .ZN(n675) );
  NAND2_X1 U638 ( .A1(n533), .A2(n675), .ZN(n535) );
  OR2_X1 U639 ( .A1(n542), .A2(n544), .ZN(n684) );
  NAND2_X1 U640 ( .A1(n684), .A2(n679), .ZN(n621) );
  INV_X1 U641 ( .A(n621), .ZN(n715) );
  NOR2_X1 U642 ( .A1(n715), .A2(KEYINPUT80), .ZN(n534) );
  NOR2_X1 U643 ( .A1(n535), .A2(n534), .ZN(n559) );
  XNOR2_X1 U644 ( .A(n538), .B(KEYINPUT39), .ZN(n573) );
  XOR2_X1 U645 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n539) );
  INV_X1 U646 ( .A(KEYINPUT42), .ZN(n555) );
  INV_X1 U647 ( .A(n541), .ZN(n710) );
  NAND2_X1 U648 ( .A1(n710), .A2(n709), .ZN(n714) );
  INV_X1 U649 ( .A(n542), .ZN(n543) );
  INV_X1 U650 ( .A(n545), .ZN(n612) );
  XNOR2_X1 U651 ( .A(KEYINPUT105), .B(KEYINPUT28), .ZN(n548) );
  XNOR2_X1 U652 ( .A(n549), .B(n548), .ZN(n552) );
  XOR2_X1 U653 ( .A(n550), .B(KEYINPUT104), .Z(n551) );
  NOR2_X1 U654 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U655 ( .A1(n707), .A2(n562), .ZN(n554) );
  XNOR2_X1 U656 ( .A(n555), .B(n554), .ZN(n775) );
  NAND2_X1 U657 ( .A1(n774), .A2(n775), .ZN(n557) );
  XOR2_X1 U658 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n556) );
  XNOR2_X1 U659 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U660 ( .A1(n559), .A2(n558), .ZN(n570) );
  XOR2_X1 U661 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n560) );
  XNOR2_X1 U662 ( .A(n563), .B(KEYINPUT47), .ZN(n564) );
  NAND2_X1 U663 ( .A1(n564), .A2(KEYINPUT80), .ZN(n568) );
  NAND2_X1 U664 ( .A1(n384), .A2(KEYINPUT47), .ZN(n566) );
  INV_X1 U665 ( .A(KEYINPUT80), .ZN(n565) );
  NAND2_X1 U666 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U667 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X2 U668 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X1 U669 ( .A(KEYINPUT48), .B(KEYINPUT69), .ZN(n571) );
  XNOR2_X1 U670 ( .A(n572), .B(n571), .ZN(n728) );
  NOR2_X1 U671 ( .A1(n684), .A2(n573), .ZN(n689) );
  NOR2_X1 U672 ( .A1(n693), .A2(n574), .ZN(n575) );
  NAND2_X1 U673 ( .A1(n575), .A2(n709), .ZN(n576) );
  XNOR2_X1 U674 ( .A(n576), .B(KEYINPUT43), .ZN(n578) );
  NAND2_X1 U675 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U676 ( .A(n579), .B(KEYINPUT102), .ZN(n776) );
  INV_X1 U677 ( .A(n776), .ZN(n580) );
  OR2_X1 U678 ( .A1(n689), .A2(n580), .ZN(n727) );
  NOR2_X1 U679 ( .A1(n728), .A2(n727), .ZN(n625) );
  NOR2_X1 U680 ( .A1(n581), .A2(G898), .ZN(n582) );
  NOR2_X1 U681 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U682 ( .A(n611), .B(n588), .ZN(n591) );
  AND2_X1 U683 ( .A1(n696), .A2(n589), .ZN(n590) );
  AND2_X1 U684 ( .A1(n591), .A2(n590), .ZN(n654) );
  AND2_X1 U685 ( .A1(n696), .A2(n592), .ZN(n593) );
  AND2_X1 U686 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U687 ( .A1(n596), .A2(n595), .ZN(n598) );
  INV_X1 U688 ( .A(KEYINPUT32), .ZN(n597) );
  XNOR2_X1 U689 ( .A(n598), .B(n597), .ZN(n777) );
  INV_X1 U690 ( .A(n616), .ZN(n620) );
  INV_X1 U691 ( .A(n599), .ZN(n600) );
  NAND2_X1 U692 ( .A1(n601), .A2(n600), .ZN(n603) );
  XNOR2_X1 U693 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n602) );
  XNOR2_X2 U694 ( .A(n603), .B(n602), .ZN(n655) );
  INV_X1 U695 ( .A(n655), .ZN(n604) );
  NAND2_X1 U696 ( .A1(n607), .A2(n604), .ZN(n606) );
  INV_X1 U697 ( .A(KEYINPUT44), .ZN(n605) );
  NAND2_X1 U698 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U699 ( .A1(n607), .A2(KEYINPUT44), .ZN(n608) );
  NAND2_X1 U700 ( .A1(n609), .A2(n608), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n665) );
  NAND2_X1 U702 ( .A1(n655), .A2(KEYINPUT44), .ZN(n622) );
  NOR2_X1 U703 ( .A1(KEYINPUT83), .A2(n628), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n436), .A2(n626), .ZN(n630) );
  INV_X1 U705 ( .A(KEYINPUT2), .ZN(n627) );
  OR2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n436), .A2(n631), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n632), .A2(KEYINPUT83), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n436), .A2(KEYINPUT2), .ZN(n637) );
  INV_X1 U711 ( .A(KEYINPUT76), .ZN(n636) );
  BUF_X2 U712 ( .A(n732), .Z(n638) );
  XNOR2_X1 U713 ( .A(KEYINPUT108), .B(KEYINPUT62), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n645) );
  INV_X1 U716 ( .A(G952), .ZN(n644) );
  AND2_X1 U717 ( .A1(n644), .A2(G953), .ZN(n750) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(G57) );
  XOR2_X1 U719 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n650) );
  XNOR2_X1 U720 ( .A(n648), .B(KEYINPUT123), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n651), .B(n359), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U723 ( .A(n654), .B(G110), .Z(G12) );
  XOR2_X1 U724 ( .A(n655), .B(G122), .Z(G24) );
  XNOR2_X1 U725 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n661), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U729 ( .A(G101), .B(n662), .ZN(n663) );
  XNOR2_X1 U730 ( .A(n663), .B(KEYINPUT109), .ZN(G3) );
  NOR2_X1 U731 ( .A1(n665), .A2(n679), .ZN(n664) );
  XOR2_X1 U732 ( .A(G104), .B(n664), .Z(G6) );
  NOR2_X1 U733 ( .A1(n665), .A2(n684), .ZN(n670) );
  XOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n667) );
  XNOR2_X1 U735 ( .A(G107), .B(KEYINPUT26), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U737 ( .A(KEYINPUT110), .B(n668), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n670), .B(n669), .ZN(G9) );
  XOR2_X1 U739 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n673) );
  INV_X1 U740 ( .A(n684), .ZN(n671) );
  NAND2_X1 U741 ( .A1(n671), .A2(n384), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U743 ( .A(G128), .B(n674), .ZN(G30) );
  XNOR2_X1 U744 ( .A(G143), .B(n675), .ZN(G45) );
  INV_X1 U745 ( .A(n679), .ZN(n676) );
  NAND2_X1 U746 ( .A1(n384), .A2(n676), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n678), .B(G146), .ZN(G48) );
  NOR2_X1 U748 ( .A1(n679), .A2(n683), .ZN(n681) );
  XNOR2_X1 U749 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U751 ( .A(G113), .B(n682), .ZN(G15) );
  NOR2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U753 ( .A(G116), .B(n685), .Z(G18) );
  XOR2_X1 U754 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n688) );
  XNOR2_X1 U755 ( .A(G125), .B(n686), .ZN(n687) );
  XNOR2_X1 U756 ( .A(n688), .B(n687), .ZN(G27) );
  XOR2_X1 U757 ( .A(G134), .B(n689), .Z(n690) );
  XNOR2_X1 U758 ( .A(KEYINPUT116), .B(n690), .ZN(G36) );
  INV_X1 U759 ( .A(n707), .ZN(n691) );
  NAND2_X1 U760 ( .A1(n719), .A2(n691), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n692), .B(KEYINPUT120), .ZN(n737) );
  XNOR2_X1 U762 ( .A(KEYINPUT51), .B(KEYINPUT118), .ZN(n706) );
  NOR2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U764 ( .A(KEYINPUT50), .B(n695), .Z(n702) );
  XOR2_X1 U765 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n699) );
  NAND2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U767 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U770 ( .A(n706), .B(n705), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n721) );
  NOR2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U774 ( .A(KEYINPUT119), .B(n713), .Z(n717) );
  NOR2_X1 U775 ( .A1(n715), .A2(n714), .ZN(n716) );
  OR2_X1 U776 ( .A1(n717), .A2(n716), .ZN(n718) );
  AND2_X1 U777 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U778 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U779 ( .A(n722), .B(KEYINPUT52), .ZN(n723) );
  NOR2_X1 U780 ( .A1(n724), .A2(n723), .ZN(n735) );
  INV_X1 U781 ( .A(n725), .ZN(n751) );
  XNOR2_X1 U782 ( .A(KEYINPUT2), .B(KEYINPUT79), .ZN(n729) );
  NAND2_X1 U783 ( .A1(n751), .A2(n729), .ZN(n726) );
  XNOR2_X1 U784 ( .A(n726), .B(KEYINPUT82), .ZN(n731) );
  OR2_X1 U785 ( .A1(n728), .A2(n727), .ZN(n765) );
  NAND2_X1 U786 ( .A1(n765), .A2(n729), .ZN(n730) );
  NAND2_X1 U787 ( .A1(n731), .A2(n730), .ZN(n733) );
  NOR2_X1 U788 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U789 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X2 U790 ( .A1(G953), .A2(n355), .ZN(n738) );
  XNOR2_X1 U791 ( .A(KEYINPUT53), .B(n738), .ZN(G75) );
  XOR2_X1 U792 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n740) );
  XOR2_X1 U793 ( .A(n740), .B(n739), .Z(n741) );
  XNOR2_X1 U794 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U795 ( .A1(n750), .A2(n743), .ZN(G54) );
  XOR2_X1 U796 ( .A(n745), .B(n744), .Z(n746) );
  NOR2_X1 U797 ( .A1(n750), .A2(n746), .ZN(G63) );
  XNOR2_X1 U798 ( .A(n748), .B(n747), .ZN(n749) );
  NOR2_X1 U799 ( .A1(n750), .A2(n749), .ZN(G66) );
  NOR2_X1 U800 ( .A1(n751), .A2(G953), .ZN(n756) );
  NAND2_X1 U801 ( .A1(G953), .A2(G224), .ZN(n752) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n752), .ZN(n753) );
  NAND2_X1 U803 ( .A1(n753), .A2(G898), .ZN(n754) );
  XOR2_X1 U804 ( .A(KEYINPUT124), .B(n754), .Z(n755) );
  NOR2_X1 U805 ( .A1(n756), .A2(n755), .ZN(n762) );
  XOR2_X1 U806 ( .A(n757), .B(KEYINPUT125), .Z(n760) );
  NOR2_X1 U807 ( .A1(G898), .A2(n758), .ZN(n759) );
  NOR2_X1 U808 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U809 ( .A(n762), .B(n761), .Z(G69) );
  XNOR2_X1 U810 ( .A(n763), .B(n764), .ZN(n767) );
  XNOR2_X1 U811 ( .A(n765), .B(n767), .ZN(n766) );
  NOR2_X1 U812 ( .A1(G953), .A2(n766), .ZN(n772) );
  XOR2_X1 U813 ( .A(n767), .B(G227), .Z(n768) );
  NAND2_X1 U814 ( .A1(n768), .A2(G900), .ZN(n769) );
  NAND2_X1 U815 ( .A1(G953), .A2(n769), .ZN(n770) );
  XOR2_X1 U816 ( .A(KEYINPUT126), .B(n770), .Z(n771) );
  NOR2_X1 U817 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U818 ( .A(KEYINPUT127), .B(n773), .ZN(G72) );
  XNOR2_X1 U819 ( .A(n774), .B(G131), .ZN(G33) );
  XNOR2_X1 U820 ( .A(n775), .B(G137), .ZN(G39) );
  XNOR2_X1 U821 ( .A(G140), .B(n776), .ZN(G42) );
  XOR2_X1 U822 ( .A(G119), .B(n777), .Z(G21) );
endmodule

