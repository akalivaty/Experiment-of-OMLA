//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(G58), .A2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n211), .B1(new_n214), .B2(new_n217), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G58), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G226), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G1698), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(G223), .B2(G1698), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G87), .ZN(new_n253));
  OAI22_X1  g0053(.A1(new_n248), .A2(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n255), .B1(new_n257), .B2(new_n212), .ZN(new_n258));
  INV_X1    g0058(.A(new_n212), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(KEYINPUT67), .A3(new_n256), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n212), .B1(KEYINPUT66), .B2(new_n256), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT66), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G33), .A3(G41), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n264), .B2(new_n266), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G232), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n262), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G200), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G190), .B2(new_n274), .ZN(new_n277));
  INV_X1    g0077(.A(G13), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n278), .A2(new_n206), .A3(G1), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n206), .A2(G1), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n284), .A2(KEYINPUT68), .A3(new_n212), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT68), .B1(new_n284), .B2(new_n212), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n285), .A2(new_n286), .A3(new_n279), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n283), .B1(new_n287), .B2(new_n281), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT75), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n252), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(new_n206), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT7), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n293), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT74), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT74), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n294), .B2(new_n295), .ZN(new_n300));
  OAI21_X1  g0100(.A(G68), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G58), .ZN(new_n302));
  INV_X1    g0102(.A(G68), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(G20), .B1(new_n304), .B2(new_n215), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G159), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT16), .B1(new_n301), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n296), .A2(new_n297), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G68), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(KEYINPUT16), .A3(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n284), .A2(new_n212), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n277), .B(new_n290), .C1(new_n310), .C2(new_n315), .ZN(new_n316));
  XOR2_X1   g0116(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n310), .A2(new_n315), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT17), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(KEYINPUT77), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n319), .A2(new_n290), .A3(new_n277), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n274), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n262), .A2(new_n271), .A3(new_n273), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT76), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n326), .A2(new_n331), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n290), .B1(new_n310), .B2(new_n315), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT18), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT18), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(new_n337), .A3(new_n334), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n324), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n279), .A2(new_n314), .ZN(new_n340));
  INV_X1    g0140(.A(new_n282), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(G77), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G77), .B2(new_n280), .ZN(new_n343));
  INV_X1    g0143(.A(new_n281), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n306), .B1(G20), .B2(G77), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n206), .A2(G33), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n343), .B1(new_n348), .B2(new_n314), .ZN(new_n349));
  AOI21_X1  g0149(.A(G1698), .B1(new_n292), .B2(new_n293), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G232), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n292), .A2(new_n293), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(G238), .A3(G1698), .ZN(new_n353));
  INV_X1    g0153(.A(G107), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n351), .B(new_n353), .C1(new_n354), .C2(new_n352), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n261), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n272), .A2(G244), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n271), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n349), .B1(new_n358), .B2(new_n325), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n358), .A2(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n356), .A2(G190), .A3(new_n271), .A4(new_n357), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n362), .A2(new_n349), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(G200), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n350), .A2(G222), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n352), .A2(G223), .A3(G1698), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n367), .B(new_n368), .C1(new_n202), .C2(new_n352), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n261), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n272), .A2(G226), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n271), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n327), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n285), .A2(new_n286), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n306), .A2(G150), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n377), .B1(new_n201), .B2(new_n206), .C1(new_n281), .C2(new_n346), .ZN(new_n378));
  INV_X1    g0178(.A(G50), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n376), .A2(new_n378), .B1(new_n379), .B2(new_n279), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n287), .A2(G50), .A3(new_n341), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n372), .A2(new_n325), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n374), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n382), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n373), .A2(G190), .B1(new_n385), .B2(KEYINPUT9), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT10), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT9), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n372), .A2(G200), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n387), .B1(new_n386), .B2(new_n389), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n366), .B(new_n384), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n306), .A2(G50), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n393), .B1(new_n206), .B2(G68), .C1(new_n202), .C2(new_n346), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n376), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT11), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n376), .A2(KEYINPUT11), .A3(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT70), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT71), .B1(new_n279), .B2(new_n303), .ZN(new_n401));
  XOR2_X1   g0201(.A(new_n401), .B(KEYINPUT12), .Z(new_n402));
  NOR2_X1   g0202(.A1(new_n282), .A2(new_n303), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(new_n340), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT70), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n397), .A2(new_n405), .A3(new_n398), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n400), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT73), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT73), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n400), .A2(new_n404), .A3(new_n409), .A4(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT72), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT14), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(new_n266), .A3(new_n259), .ZN(new_n415));
  INV_X1    g0215(.A(new_n270), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT69), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT69), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n419), .A3(new_n416), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(G238), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT13), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G97), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n230), .A2(G1698), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(G226), .B2(G1698), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n423), .B1(new_n425), .B2(new_n251), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n261), .B1(new_n267), .B2(new_n270), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n421), .A2(new_n422), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n422), .B1(new_n421), .B2(new_n427), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n413), .B(G169), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n415), .A2(new_n419), .A3(new_n416), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n419), .B1(new_n415), .B2(new_n416), .ZN(new_n432));
  INV_X1    g0232(.A(G238), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n426), .A2(new_n261), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n271), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n421), .A2(new_n422), .A3(new_n427), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(G179), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n413), .B1(new_n441), .B2(G169), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n412), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(G169), .B1(new_n428), .B2(new_n429), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT14), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n445), .A2(KEYINPUT72), .A3(new_n439), .A4(new_n430), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n411), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n407), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n441), .A2(G200), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n437), .A2(G190), .A3(new_n438), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NOR4_X1   g0251(.A1(new_n339), .A2(new_n392), .A3(new_n447), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n352), .A2(G257), .A3(G1698), .ZN(new_n453));
  INV_X1    g0253(.A(G1698), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n352), .A2(G250), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G294), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n261), .ZN(new_n458));
  NOR2_X1   g0258(.A1(KEYINPUT80), .A2(G41), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT5), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(KEYINPUT80), .B2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n269), .A2(G1), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G264), .A3(new_n415), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n458), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n205), .A2(G45), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(KEYINPUT5), .B2(new_n459), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n468), .A2(new_n415), .A3(G274), .A4(new_n462), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n327), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n458), .A2(new_n469), .A3(new_n465), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n325), .ZN(new_n472));
  INV_X1    g0272(.A(new_n314), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G116), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G20), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT23), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n206), .B2(G107), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n354), .A2(KEYINPUT23), .A3(G20), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n206), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n480), .A2(KEYINPUT22), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(KEYINPUT22), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT24), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(new_n479), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n473), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OR3_X1    g0287(.A1(new_n252), .A2(KEYINPUT78), .A3(G1), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT78), .B1(new_n252), .B2(G1), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n287), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n354), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n279), .A2(new_n354), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n493), .B(KEYINPUT25), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n470), .B(new_n472), .C1(new_n487), .C2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  OAI211_X1 g0297(.A(G264), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n498));
  OAI211_X1 g0298(.A(G257), .B(new_n454), .C1(new_n249), .C2(new_n250), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n292), .A2(G303), .A3(new_n293), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n261), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n464), .A2(new_n415), .A3(G270), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n469), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G169), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n340), .A2(new_n490), .A3(G116), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n278), .A2(G1), .ZN(new_n507));
  INV_X1    g0307(.A(G116), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(G20), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n284), .A2(new_n212), .B1(G20), .B2(new_n508), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  INV_X1    g0312(.A(G97), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n206), .C1(G33), .C2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n511), .A2(KEYINPUT20), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT20), .B1(new_n511), .B2(new_n514), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n497), .B1(new_n505), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n504), .A2(KEYINPUT21), .A3(G169), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n502), .A2(G179), .A3(new_n469), .A4(new_n503), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n518), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT85), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT85), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n525), .B(new_n518), .C1(new_n520), .C2(new_n521), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n496), .B(new_n519), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n487), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n466), .A2(G190), .A3(new_n469), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n492), .A2(new_n494), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n471), .A2(G200), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n504), .A2(G200), .ZN(new_n533));
  INV_X1    g0333(.A(G190), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n518), .C1(new_n534), .C2(new_n504), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n527), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT84), .ZN(new_n538));
  INV_X1    g0338(.A(new_n512), .ZN(new_n539));
  AND2_X1   g0339(.A1(KEYINPUT4), .A2(G244), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n350), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G244), .B(new_n454), .C1(new_n249), .C2(new_n250), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT4), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G250), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT79), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n352), .A2(KEYINPUT79), .A3(G250), .A4(G1698), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n541), .A2(new_n544), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n261), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n464), .A2(new_n415), .A3(G257), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n469), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AND4_X1   g0353(.A1(KEYINPUT81), .A2(new_n550), .A3(G190), .A4(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n552), .B1(new_n549), .B2(new_n261), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT81), .B1(new_n555), .B2(G190), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n275), .B1(new_n550), .B2(new_n553), .ZN(new_n558));
  OAI21_X1  g0358(.A(G107), .B1(new_n298), .B2(new_n300), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n354), .A2(KEYINPUT6), .A3(G97), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n513), .A2(new_n354), .ZN(new_n561));
  NOR2_X1   g0361(.A1(G97), .A2(G107), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n560), .B1(new_n563), .B2(KEYINPUT6), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(G20), .B1(G77), .B2(new_n306), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n473), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n280), .A2(G97), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n491), .B2(new_n513), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n558), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  AOI211_X1 g0370(.A(G179), .B(new_n552), .C1(new_n261), .C2(new_n549), .ZN(new_n571));
  AOI21_X1  g0371(.A(G169), .B1(new_n550), .B2(new_n553), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n569), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n559), .A2(new_n565), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(new_n473), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n557), .A2(new_n570), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G244), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n578));
  OAI211_X1 g0378(.A(G238), .B(new_n454), .C1(new_n249), .C2(new_n250), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n579), .A3(new_n474), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n261), .ZN(new_n581));
  AOI21_X1  g0381(.A(G250), .B1(new_n205), .B2(G45), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n263), .B2(new_n463), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n415), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n206), .B1(new_n423), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n562), .A2(new_n253), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n206), .B(G68), .C1(new_n249), .C2(new_n250), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n586), .B1(new_n346), .B2(new_n513), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n314), .B1(new_n279), .B2(new_n347), .ZN(new_n593));
  INV_X1    g0393(.A(new_n347), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n287), .A2(new_n594), .A3(new_n490), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n585), .A2(new_n325), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n580), .A2(new_n261), .B1(new_n415), .B2(new_n583), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n327), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT82), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT82), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n597), .A2(new_n600), .A3(new_n327), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT83), .B1(new_n585), .B2(new_n534), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT83), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n597), .A2(new_n604), .A3(G190), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n375), .A2(G87), .A3(new_n280), .A4(new_n490), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n592), .A2(new_n314), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n347), .A2(new_n279), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(G200), .B2(new_n585), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n596), .A2(new_n602), .B1(new_n606), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n538), .B1(new_n577), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n566), .A2(new_n569), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n550), .A2(G190), .A3(new_n553), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT81), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n550), .A2(new_n553), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G200), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n555), .A2(KEYINPUT81), .A3(G190), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n614), .A2(new_n617), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n555), .A2(new_n327), .ZN(new_n622));
  OAI221_X1 g0422(.A(new_n622), .B1(G169), .B2(new_n555), .C1(new_n566), .C2(new_n569), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n538), .A2(new_n612), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n452), .B(new_n537), .C1(new_n613), .C2(new_n624), .ZN(new_n625));
  XOR2_X1   g0425(.A(new_n625), .B(KEYINPUT86), .Z(G372));
  INV_X1    g0426(.A(new_n384), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n451), .A2(new_n361), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n324), .B1(new_n628), .B2(new_n447), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(new_n336), .A3(new_n338), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n390), .A2(new_n391), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n596), .A2(new_n598), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT88), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n610), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n593), .A2(KEYINPUT88), .A3(new_n607), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT87), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n585), .A2(new_n639), .A3(G200), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT87), .B1(new_n597), .B2(new_n275), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n638), .A2(new_n642), .A3(KEYINPUT89), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n606), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT89), .B1(new_n638), .B2(new_n642), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n633), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n621), .A2(new_n532), .A3(new_n623), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n522), .A2(new_n523), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n496), .A2(new_n519), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n634), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n602), .A2(new_n596), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n606), .A2(new_n611), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n654), .A2(new_n623), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n614), .A2(new_n572), .A3(new_n571), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n658), .B(new_n633), .C1(new_n644), .C2(new_n645), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n657), .B1(new_n660), .B2(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n651), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n452), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n632), .A2(new_n663), .ZN(G369));
  NAND2_X1  g0464(.A1(new_n507), .A2(new_n206), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(G213), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n496), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n519), .B1(new_n524), .B2(new_n526), .ZN(new_n672));
  INV_X1    g0472(.A(new_n670), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT91), .Z(new_n675));
  AOI21_X1  g0475(.A(new_n673), .B1(new_n528), .B2(new_n530), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT90), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n532), .B1(new_n676), .B2(new_n677), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n496), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n671), .B1(new_n675), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n649), .A2(new_n519), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n523), .A2(new_n670), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n535), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n672), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  INV_X1    g0486(.A(new_n671), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n680), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n681), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT92), .Z(G399));
  INV_X1    g0492(.A(new_n209), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n588), .A2(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n217), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n655), .B1(new_n654), .B2(new_n623), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n659), .B2(new_n655), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n621), .A2(new_n532), .A3(new_n623), .ZN(new_n702));
  INV_X1    g0502(.A(new_n645), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n606), .A3(new_n643), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n702), .A2(new_n527), .A3(new_n633), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n701), .A2(new_n705), .A3(new_n633), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT29), .A3(new_n673), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n670), .B1(new_n651), .B2(new_n661), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(KEYINPUT29), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n537), .B(new_n673), .C1(new_n613), .C2(new_n624), .ZN(new_n711));
  INV_X1    g0511(.A(new_n521), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n466), .A3(new_n555), .A4(new_n597), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(KEYINPUT30), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n458), .A2(new_n465), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n717), .A2(new_n521), .A3(new_n585), .ZN(new_n718));
  INV_X1    g0518(.A(new_n715), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n555), .A3(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n504), .A2(new_n327), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n618), .A3(new_n585), .A4(new_n471), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n716), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT31), .B1(new_n723), .B2(new_n670), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n710), .B1(new_n711), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n709), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n699), .B1(new_n731), .B2(G1), .ZN(G364));
  NOR2_X1   g0532(.A1(new_n278), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n205), .B1(new_n733), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n694), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n686), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n685), .A2(G330), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n685), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n212), .B1(G20), .B2(new_n325), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n693), .A2(new_n251), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n748), .A2(G355), .B1(new_n508), .B2(new_n693), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n693), .A2(new_n352), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G45), .B2(new_n217), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n244), .A2(new_n269), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n747), .B1(new_n753), .B2(KEYINPUT95), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(KEYINPUT95), .B2(new_n753), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n206), .A2(G179), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G190), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT32), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n206), .A2(new_n327), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n534), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n762), .A2(G190), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n760), .B1(new_n764), .B2(new_n379), .C1(new_n303), .C2(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n534), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n206), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n758), .A2(KEYINPUT32), .A3(new_n759), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G87), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n756), .A2(new_n534), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G107), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n771), .A2(new_n772), .A3(new_n775), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n761), .A2(new_n757), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n761), .A2(G190), .A3(new_n275), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n352), .B1(new_n780), .B2(new_n202), .C1(new_n302), .C2(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n767), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n781), .ZN(new_n784));
  INV_X1    g0584(.A(new_n758), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n784), .A2(G322), .B1(new_n785), .B2(G329), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n786), .B(new_n251), .C1(new_n787), .C2(new_n780), .ZN(new_n788));
  INV_X1    g0588(.A(G317), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(KEYINPUT33), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(KEYINPUT33), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n765), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n763), .A2(G326), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n769), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  INV_X1    g0596(.A(G303), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n796), .A2(new_n776), .B1(new_n773), .B2(new_n797), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n788), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n745), .B1(new_n783), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n736), .B(KEYINPUT94), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n755), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n738), .A2(new_n739), .B1(new_n744), .B2(new_n802), .ZN(G396));
  OAI21_X1  g0603(.A(new_n365), .B1(new_n349), .B2(new_n673), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n361), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n359), .A2(new_n360), .A3(new_n673), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n708), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n702), .A2(new_n633), .A3(new_n704), .A4(new_n650), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n633), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n656), .B1(new_n659), .B2(new_n655), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n673), .B(new_n809), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n736), .B1(new_n815), .B2(new_n729), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n729), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n745), .A2(new_n740), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n801), .B1(G77), .B2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT96), .Z(new_n821));
  OAI22_X1  g0621(.A1(new_n764), .A2(new_n797), .B1(new_n773), .B2(new_n354), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G87), .B2(new_n777), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n352), .B1(new_n784), .B2(G294), .ZN(new_n824));
  INV_X1    g0624(.A(new_n780), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G116), .A2(new_n825), .B1(new_n785), .B2(G311), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G97), .A2(new_n770), .B1(new_n765), .B2(G283), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n823), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n784), .A2(G143), .B1(new_n825), .B2(G159), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  INV_X1    g0630(.A(G150), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n764), .B2(new_n830), .C1(new_n831), .C2(new_n766), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n777), .A2(G68), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n251), .B1(new_n785), .B2(G132), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n770), .A2(G58), .B1(new_n774), .B2(G50), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n832), .A2(new_n833), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n828), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n821), .B1(new_n745), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n809), .B2(new_n741), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n817), .A2(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n733), .A2(new_n205), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n443), .A2(new_n446), .ZN(new_n845));
  INV_X1    g0645(.A(new_n411), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n451), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n670), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n846), .B(new_n670), .C1(new_n845), .C2(new_n451), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n711), .A2(new_n727), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n852), .A2(new_n853), .A3(new_n809), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT99), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT16), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n303), .B1(new_n296), .B2(new_n297), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n308), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n313), .A2(new_n376), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n288), .B(KEYINPUT75), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT98), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT98), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n290), .A2(new_n863), .A3(new_n859), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n333), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n668), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n862), .A2(new_n866), .A3(new_n864), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n867), .A3(new_n316), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n334), .A2(new_n866), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n335), .A2(new_n870), .A3(new_n871), .A4(new_n316), .ZN(new_n872));
  INV_X1    g0672(.A(new_n867), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n869), .A2(new_n872), .B1(new_n339), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n855), .B1(new_n874), .B2(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n869), .A2(new_n872), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n339), .A2(new_n873), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n855), .A4(KEYINPUT38), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(KEYINPUT38), .B2(new_n874), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n854), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n335), .A2(new_n316), .A3(new_n871), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(KEYINPUT100), .A3(new_n872), .ZN(new_n886));
  INV_X1    g0686(.A(new_n871), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n339), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT100), .B1(new_n885), .B2(new_n872), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n874), .A2(KEYINPUT38), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n882), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n880), .A2(new_n881), .B1(new_n854), .B2(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT102), .Z(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n452), .A2(new_n853), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT103), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n710), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n898), .B2(new_n896), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT39), .B1(new_n879), .B2(new_n875), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n891), .A2(new_n902), .A3(new_n892), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n447), .A2(new_n673), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n866), .B1(new_n336), .B2(new_n338), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n879), .A2(new_n875), .ZN(new_n909));
  INV_X1    g0709(.A(new_n852), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n807), .B2(new_n814), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n452), .B(new_n707), .C1(new_n708), .C2(KEYINPUT29), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n632), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n844), .B1(new_n900), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n916), .B2(new_n900), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n217), .A2(new_n202), .A3(new_n304), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n303), .A2(G50), .ZN(new_n920));
  OAI211_X1 g0720(.A(G1), .B(new_n278), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n508), .B(new_n214), .C1(new_n564), .C2(KEYINPUT35), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(KEYINPUT35), .B2(new_n564), .ZN(new_n923));
  XNOR2_X1  g0723(.A(KEYINPUT97), .B(KEYINPUT36), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n918), .A2(new_n921), .A3(new_n925), .ZN(G367));
  NAND3_X1  g0726(.A1(new_n636), .A2(new_n637), .A3(new_n670), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n704), .A2(new_n633), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n633), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n577), .B1(new_n614), .B2(new_n673), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n623), .B2(new_n673), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT104), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT105), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(new_n496), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n673), .B1(new_n936), .B2(new_n658), .ZN(new_n937));
  INV_X1    g0737(.A(new_n934), .ZN(new_n938));
  INV_X1    g0738(.A(new_n688), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n675), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT42), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT106), .Z(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n931), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n935), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n943), .A2(new_n931), .A3(new_n946), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n948), .A2(new_n689), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n950), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n952), .A2(new_n947), .B1(new_n690), .B2(new_n935), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n694), .B(KEYINPUT41), .Z(new_n954));
  OR2_X1    g0754(.A1(new_n675), .A2(new_n939), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT108), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n686), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n957), .A3(new_n940), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n686), .A2(new_n956), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n958), .B(new_n959), .Z(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(new_n730), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n681), .A2(new_n934), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n681), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n966), .A2(KEYINPUT44), .A3(new_n938), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT44), .B1(new_n966), .B2(new_n938), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n689), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n964), .B(new_n690), .C1(new_n968), .C2(new_n967), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n961), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n954), .B1(new_n972), .B2(new_n731), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n951), .B(new_n953), .C1(new_n735), .C2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n750), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n746), .B1(new_n209), .B2(new_n347), .C1(new_n975), .C2(new_n236), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n801), .A2(new_n976), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n780), .A2(new_n379), .B1(new_n758), .B2(new_n830), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n251), .B(new_n978), .C1(G150), .C2(new_n784), .ZN(new_n979));
  INV_X1    g0779(.A(G143), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n979), .B1(new_n980), .B2(new_n764), .C1(new_n759), .C2(new_n766), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n770), .A2(G68), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n302), .B2(new_n773), .C1(new_n202), .C2(new_n776), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n765), .A2(G294), .B1(new_n777), .B2(G97), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n354), .B2(new_n769), .C1(new_n787), .C2(new_n764), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n784), .A2(G303), .B1(new_n785), .B2(G317), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT46), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n773), .B2(new_n508), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n774), .A2(KEYINPUT46), .A3(G116), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n352), .B1(new_n825), .B2(G283), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n986), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n981), .A2(new_n983), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT47), .Z(new_n993));
  INV_X1    g0793(.A(new_n745), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n977), .B1(new_n993), .B2(new_n994), .C1(new_n929), .C2(new_n743), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n974), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT109), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n974), .A2(KEYINPUT109), .A3(new_n995), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(G387));
  INV_X1    g0800(.A(new_n961), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n960), .A2(new_n730), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1001), .A2(new_n694), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n696), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n748), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(G107), .B2(new_n209), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n233), .A2(new_n269), .ZN(new_n1007));
  AOI211_X1 g0807(.A(G45), .B(new_n1004), .C1(G68), .C2(G77), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n281), .A2(G50), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT50), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n975), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1006), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n801), .B1(new_n1012), .B2(new_n747), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n774), .A2(G77), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n347), .B2(new_n769), .C1(new_n766), .C2(new_n281), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G68), .A2(new_n825), .B1(new_n785), .B2(G150), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1016), .B(new_n352), .C1(new_n379), .C2(new_n781), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n764), .A2(new_n759), .B1(new_n776), .B2(new_n513), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT110), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n352), .B1(new_n785), .B2(G326), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n769), .A2(new_n796), .B1(new_n773), .B2(new_n794), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n784), .A2(G317), .B1(new_n825), .B2(G303), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n763), .A2(G322), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(new_n787), .C2(new_n766), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n1026), .B2(new_n1025), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1021), .B1(new_n508), .B2(new_n776), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1020), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT111), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n994), .B1(new_n1032), .B2(KEYINPUT111), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1013), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n939), .B2(new_n743), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1003), .B(new_n1036), .C1(new_n734), .C2(new_n960), .ZN(G393));
  INV_X1    g0837(.A(KEYINPUT112), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n970), .A2(new_n971), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n1001), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1040), .A2(new_n694), .A3(new_n972), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n970), .A2(new_n735), .A3(new_n971), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n241), .A2(new_n975), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n746), .B1(new_n513), .B2(new_n209), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n801), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G150), .A2(new_n763), .B1(new_n784), .B2(G159), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT51), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n352), .B1(new_n758), .B2(new_n980), .C1(new_n281), .C2(new_n780), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n766), .A2(new_n379), .B1(new_n776), .B2(new_n253), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n769), .A2(new_n202), .B1(new_n773), .B2(new_n303), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G317), .A2(new_n763), .B1(new_n784), .B2(G311), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT52), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n352), .B1(new_n785), .B2(G322), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n794), .B2(new_n780), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n778), .B1(new_n796), .B2(new_n773), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n766), .A2(new_n797), .B1(new_n508), .B2(new_n769), .ZN(new_n1057));
  NOR4_X1   g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1051), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1045), .B1(new_n1059), .B2(new_n745), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n949), .B2(new_n743), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1042), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1038), .B1(new_n1041), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1041), .A2(new_n1063), .A3(new_n1038), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(G390));
  NAND3_X1  g0867(.A1(new_n728), .A2(new_n852), .A3(new_n809), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT114), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n901), .B(new_n903), .C1(new_n906), .C2(new_n911), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n706), .A2(new_n673), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n807), .B1(new_n1072), .B2(new_n806), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n852), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n905), .A2(KEYINPUT113), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT113), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n447), .A2(new_n1076), .A3(new_n673), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n891), .B2(new_n892), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n728), .A2(new_n852), .A3(new_n809), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1074), .A2(new_n1079), .B1(new_n1080), .B2(KEYINPUT114), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1070), .B1(new_n1071), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1071), .A2(new_n1070), .A3(new_n1081), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n452), .A2(new_n728), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n914), .A2(new_n632), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n853), .A2(G330), .A3(new_n809), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n910), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n634), .B1(new_n648), .B2(new_n527), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n670), .B1(new_n1089), .B2(new_n701), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n808), .B1(new_n1090), .B2(new_n805), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1088), .A2(new_n1068), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n808), .B1(new_n708), .B2(new_n809), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1088), .B2(new_n1068), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1086), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1083), .A2(new_n1084), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n914), .A2(new_n632), .A3(new_n1085), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n814), .A2(new_n807), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n852), .B1(new_n728), .B2(new_n809), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n1080), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1088), .A2(new_n1091), .A3(new_n1068), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1071), .A2(new_n1070), .A3(new_n1081), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n1082), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1096), .A2(new_n1104), .A3(new_n694), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n801), .B1(new_n344), .B2(new_n819), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n765), .A2(G107), .B1(new_n825), .B2(G97), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT117), .Z(new_n1108));
  OAI21_X1  g0908(.A(new_n251), .B1(new_n781), .B2(new_n508), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G294), .B2(new_n785), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G77), .A2(new_n770), .B1(new_n763), .B2(G283), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1110), .A2(new_n1111), .A3(new_n775), .A4(new_n835), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n773), .A2(new_n831), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1114));
  XNOR2_X1  g0914(.A(new_n1113), .B(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G159), .A2(new_n770), .B1(new_n763), .B2(G128), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n251), .B1(new_n785), .B2(G125), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n784), .A2(G132), .B1(new_n825), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n765), .A2(G137), .B1(new_n777), .B2(G50), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1116), .A2(new_n1117), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1108), .A2(new_n1112), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1106), .B1(new_n1123), .B2(new_n745), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n904), .B2(new_n741), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT115), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n735), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1126), .B(new_n735), .C1(new_n1103), .C2(new_n1082), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1105), .B(new_n1125), .C1(new_n1128), .C2(new_n1130), .ZN(G378));
  NAND2_X1  g0931(.A1(new_n880), .A2(new_n881), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n893), .A2(new_n854), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(G330), .A3(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n384), .B1(new_n390), .B2(new_n391), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n385), .A2(new_n668), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n1135), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1134), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1145), .B(KEYINPUT119), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n894), .A2(G330), .A3(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1147), .A2(new_n913), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n913), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n735), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1148), .A2(new_n740), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n776), .A2(new_n302), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n766), .A2(new_n513), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(G116), .C2(new_n763), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n251), .A2(new_n268), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n781), .A2(new_n354), .B1(new_n758), .B2(new_n796), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n594), .C2(new_n825), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1156), .A2(new_n982), .A3(new_n1014), .A4(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT58), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1157), .B(new_n379), .C1(G33), .C2(G41), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n763), .A2(G125), .ZN(new_n1163));
  INV_X1    g0963(.A(G132), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n766), .B2(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n784), .A2(G128), .B1(new_n825), .B2(G137), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n773), .B2(new_n1118), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(G150), .C2(new_n770), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n777), .A2(G159), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1161), .B(new_n1162), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT118), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n994), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n1176), .B2(new_n1175), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n737), .B1(new_n379), .B2(new_n818), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1153), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1152), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n913), .ZN(new_n1182));
  AND4_X1   g0982(.A1(G330), .A2(new_n1148), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1145), .B1(new_n894), .B2(G330), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1147), .A2(new_n913), .A3(new_n1149), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1104), .A2(new_n1086), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(KEYINPUT57), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n694), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT57), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1181), .B1(new_n1190), .B2(new_n1191), .ZN(G375));
  OAI21_X1  g0992(.A(new_n735), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n251), .B1(new_n785), .B2(G128), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n830), .B2(new_n781), .C1(new_n831), .C2(new_n780), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1154), .B(new_n1195), .C1(new_n765), .C2(new_n1119), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n769), .A2(new_n379), .B1(new_n773), .B2(new_n759), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G132), .B2(new_n763), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n766), .A2(new_n508), .B1(new_n764), .B2(new_n794), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G97), .B2(new_n774), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n769), .A2(new_n347), .B1(new_n776), .B2(new_n202), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n781), .A2(new_n796), .B1(new_n780), .B2(new_n354), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n251), .B1(new_n758), .B2(new_n797), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1196), .A2(new_n1198), .B1(new_n1200), .B2(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n801), .B1(G68), .B2(new_n819), .C1(new_n1205), .C2(new_n994), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT120), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n852), .B2(new_n741), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1193), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n954), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1100), .A2(new_n1097), .A3(new_n1101), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1095), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(G381));
  OR3_X1    g1014(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1215));
  OR3_X1    g1015(.A1(G390), .A2(G381), .A3(new_n1215), .ZN(new_n1216));
  OR4_X1    g1016(.A1(G387), .A2(new_n1216), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1017(.A(G213), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(G375), .A2(new_n1218), .A3(G343), .A4(G378), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT121), .Z(new_n1220));
  NAND3_X1  g1020(.A1(G407), .A2(G213), .A3(new_n1220), .ZN(G409));
  NAND2_X1  g1021(.A1(G390), .A2(KEYINPUT125), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT125), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1065), .A2(new_n1223), .A3(new_n1066), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1222), .A2(new_n998), .A3(new_n999), .A4(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(G393), .B(G396), .Z(new_n1226));
  INV_X1    g1026(.A(new_n996), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(G390), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1227), .A2(G390), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n996), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1226), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT127), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT62), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1218), .A2(G343), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G378), .B(new_n1181), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1105), .A2(new_n1125), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1187), .A2(new_n1188), .A3(new_n1211), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1152), .A2(new_n1180), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1238), .B(new_n1239), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1236), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT122), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1100), .A2(new_n1097), .A3(new_n1101), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n694), .B1(new_n1246), .B2(KEYINPUT60), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1095), .B2(new_n1212), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1245), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT60), .B1(new_n1246), .B2(new_n1102), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n695), .B1(new_n1212), .B2(new_n1248), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(KEYINPUT122), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G384), .B1(new_n1254), .B2(new_n1210), .ZN(new_n1255));
  INV_X1    g1055(.A(G384), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1256), .B(new_n1209), .C1(new_n1250), .C2(new_n1253), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1244), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1251), .A2(KEYINPUT122), .A3(new_n1252), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT122), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1210), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1256), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1254), .A2(G384), .A3(new_n1210), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(KEYINPUT123), .A3(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1258), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1235), .B1(new_n1243), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1243), .A2(new_n1265), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1266), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1236), .A2(G2897), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1258), .A2(new_n1264), .A3(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G2897), .B(new_n1236), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT124), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1243), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1272), .A2(KEYINPUT124), .A3(new_n1273), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1270), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AOI211_X1 g1080(.A(KEYINPUT126), .B(KEYINPUT61), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1233), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1229), .A2(new_n1232), .B1(KEYINPUT63), .B2(new_n1268), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1283), .B(new_n1278), .C1(new_n1268), .C2(KEYINPUT63), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(G405));
  XNOR2_X1  g1085(.A(G375), .B(G378), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1265), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1288), .B2(new_n1286), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1233), .B(new_n1289), .ZN(G402));
endmodule


