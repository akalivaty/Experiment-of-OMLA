

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746;

  XNOR2_X1 U378 ( .A(n372), .B(n358), .ZN(n532) );
  XNOR2_X1 U379 ( .A(n373), .B(G146), .ZN(n493) );
  XNOR2_X1 U380 ( .A(n498), .B(n719), .ZN(n627) );
  INV_X1 U381 ( .A(G953), .ZN(n739) );
  OR2_X1 U382 ( .A1(n404), .A2(n512), .ZN(n356) );
  XNOR2_X2 U383 ( .A(KEYINPUT4), .B(KEYINPUT65), .ZN(n728) );
  NAND2_X1 U384 ( .A1(n401), .A2(n399), .ZN(n398) );
  NOR2_X2 U385 ( .A1(n684), .A2(n682), .ZN(n689) );
  NAND2_X1 U386 ( .A1(n375), .A2(n386), .ZN(n374) );
  XNOR2_X2 U387 ( .A(n374), .B(n588), .ZN(n712) );
  NOR2_X1 U388 ( .A1(n400), .A2(n688), .ZN(n399) );
  XOR2_X1 U389 ( .A(G131), .B(KEYINPUT67), .Z(n476) );
  XNOR2_X1 U390 ( .A(n493), .B(n435), .ZN(n477) );
  AND2_X2 U391 ( .A1(n365), .A2(n546), .ZN(n657) );
  XNOR2_X1 U392 ( .A(n366), .B(n363), .ZN(n365) );
  NOR2_X1 U393 ( .A1(n561), .A2(n505), .ZN(n407) );
  NAND2_X1 U394 ( .A1(n395), .A2(n393), .ZN(n392) );
  NOR2_X1 U395 ( .A1(n394), .A2(KEYINPUT86), .ZN(n393) );
  INV_X1 U396 ( .A(G469), .ZN(n455) );
  XNOR2_X1 U397 ( .A(n429), .B(n428), .ZN(n430) );
  INV_X1 U398 ( .A(KEYINPUT94), .ZN(n428) );
  XNOR2_X1 U399 ( .A(G110), .B(G119), .ZN(n429) );
  XOR2_X1 U400 ( .A(G113), .B(G104), .Z(n487) );
  NOR2_X1 U401 ( .A1(n542), .A2(n522), .ZN(n370) );
  OR2_X1 U402 ( .A1(n621), .A2(G902), .ZN(n372) );
  XNOR2_X1 U403 ( .A(n384), .B(KEYINPUT22), .ZN(n585) );
  NOR2_X1 U404 ( .A1(n645), .A2(n683), .ZN(n515) );
  XNOR2_X1 U405 ( .A(n468), .B(n406), .ZN(n727) );
  INV_X1 U406 ( .A(n476), .ZN(n406) );
  XNOR2_X1 U407 ( .A(G107), .B(G116), .ZN(n465) );
  XNOR2_X1 U408 ( .A(n377), .B(G134), .ZN(n468) );
  INV_X1 U409 ( .A(n607), .ZN(n390) );
  XNOR2_X1 U410 ( .A(n727), .B(G146), .ZN(n454) );
  XNOR2_X1 U411 ( .A(n728), .B(G101), .ZN(n448) );
  INV_X1 U412 ( .A(G125), .ZN(n373) );
  OR2_X1 U413 ( .A1(G902), .A2(G237), .ZN(n409) );
  XNOR2_X1 U414 ( .A(n565), .B(n564), .ZN(n575) );
  NOR2_X1 U415 ( .A1(n669), .A2(n668), .ZN(n565) );
  NAND2_X1 U416 ( .A1(n503), .A2(n590), .ZN(n403) );
  OR2_X1 U417 ( .A1(n627), .A2(n402), .ZN(n401) );
  NAND2_X1 U418 ( .A1(G234), .A2(G237), .ZN(n457) );
  XNOR2_X1 U419 ( .A(n447), .B(n383), .ZN(n718) );
  INV_X1 U420 ( .A(G110), .ZN(n383) );
  XNOR2_X1 U421 ( .A(G107), .B(G104), .ZN(n447) );
  XNOR2_X1 U422 ( .A(n448), .B(n718), .ZN(n495) );
  XNOR2_X1 U423 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n494) );
  NAND2_X1 U424 ( .A1(n589), .A2(n658), .ZN(n661) );
  XNOR2_X1 U425 ( .A(n537), .B(KEYINPUT41), .ZN(n679) );
  AND2_X1 U426 ( .A1(n577), .A2(n407), .ZN(n462) );
  XNOR2_X1 U427 ( .A(n436), .B(n726), .ZN(n614) );
  XNOR2_X1 U428 ( .A(n434), .B(n411), .ZN(n436) );
  XNOR2_X1 U429 ( .A(n431), .B(n430), .ZN(n434) );
  XNOR2_X1 U430 ( .A(n491), .B(n490), .ZN(n621) );
  AND2_X1 U431 ( .A1(n598), .A2(G953), .ZN(n711) );
  XNOR2_X1 U432 ( .A(n368), .B(KEYINPUT108), .ZN(n742) );
  NOR2_X1 U433 ( .A1(n369), .A2(n669), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n370), .B(n523), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n560), .B(n559), .ZN(n606) );
  AND2_X1 U436 ( .A1(n585), .A2(n410), .ZN(n560) );
  NAND2_X1 U437 ( .A1(n532), .A2(n371), .ZN(n644) );
  INV_X1 U438 ( .A(n533), .ZN(n371) );
  INV_X1 U439 ( .A(n532), .ZN(n513) );
  NOR2_X1 U440 ( .A1(n566), .A2(n580), .ZN(n357) );
  INV_X1 U441 ( .A(n666), .ZN(n408) );
  XOR2_X1 U442 ( .A(KEYINPUT13), .B(G475), .Z(n358) );
  AND2_X1 U443 ( .A1(n606), .A2(n605), .ZN(n359) );
  AND2_X1 U444 ( .A1(n526), .A2(n525), .ZN(n360) );
  AND2_X1 U445 ( .A1(n401), .A2(n403), .ZN(n361) );
  INV_X1 U446 ( .A(KEYINPUT86), .ZN(n512) );
  XOR2_X1 U447 ( .A(KEYINPUT87), .B(KEYINPUT33), .Z(n362) );
  XOR2_X1 U448 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n363) );
  XOR2_X1 U449 ( .A(KEYINPUT82), .B(KEYINPUT46), .Z(n364) );
  NAND2_X1 U450 ( .A1(n360), .A2(n367), .ZN(n366) );
  XNOR2_X1 U451 ( .A(n405), .B(n364), .ZN(n367) );
  XNOR2_X1 U452 ( .A(n376), .B(KEYINPUT85), .ZN(n375) );
  NAND2_X1 U453 ( .A1(n391), .A2(n587), .ZN(n376) );
  XNOR2_X1 U454 ( .A(n377), .B(n494), .ZN(n380) );
  XNOR2_X2 U455 ( .A(G143), .B(G128), .ZN(n377) );
  INV_X1 U456 ( .A(n568), .ZN(n692) );
  XNOR2_X2 U457 ( .A(n378), .B(n362), .ZN(n568) );
  NAND2_X1 U458 ( .A1(n575), .A2(n583), .ZN(n378) );
  XOR2_X2 U459 ( .A(G137), .B(G140), .Z(n449) );
  XNOR2_X1 U460 ( .A(n495), .B(n379), .ZN(n498) );
  XNOR2_X1 U461 ( .A(n381), .B(n380), .ZN(n379) );
  XNOR2_X1 U462 ( .A(n382), .B(n493), .ZN(n381) );
  NAND2_X1 U463 ( .A1(n739), .A2(G224), .ZN(n382) );
  NOR2_X2 U464 ( .A1(n566), .A2(n556), .ZN(n384) );
  XNOR2_X2 U465 ( .A(n385), .B(KEYINPUT0), .ZN(n566) );
  NAND2_X1 U466 ( .A1(n555), .A2(n554), .ZN(n385) );
  NAND2_X1 U467 ( .A1(n574), .A2(n387), .ZN(n386) );
  NAND2_X1 U468 ( .A1(n389), .A2(n388), .ZN(n387) );
  INV_X1 U469 ( .A(KEYINPUT44), .ZN(n388) );
  NAND2_X1 U470 ( .A1(n359), .A2(n390), .ZN(n389) );
  NAND2_X1 U471 ( .A1(n607), .A2(KEYINPUT44), .ZN(n391) );
  NAND2_X2 U472 ( .A1(n396), .A2(n392), .ZN(n522) );
  INV_X1 U473 ( .A(n404), .ZN(n394) );
  INV_X1 U474 ( .A(n398), .ZN(n395) );
  AND2_X2 U475 ( .A1(n397), .A2(n356), .ZN(n396) );
  NAND2_X1 U476 ( .A1(n398), .A2(KEYINPUT86), .ZN(n397) );
  NAND2_X1 U477 ( .A1(n404), .A2(n361), .ZN(n511) );
  INV_X1 U478 ( .A(n403), .ZN(n400) );
  OR2_X1 U479 ( .A1(n503), .A2(n590), .ZN(n402) );
  NAND2_X1 U480 ( .A1(n627), .A2(n503), .ZN(n404) );
  NAND2_X1 U481 ( .A1(n745), .A2(n744), .ZN(n405) );
  NOR2_X1 U482 ( .A1(n524), .A2(n408), .ZN(n577) );
  XNOR2_X1 U483 ( .A(n597), .B(n596), .ZN(n600) );
  NAND2_X1 U484 ( .A1(n661), .A2(n590), .ZN(n595) );
  NAND2_X1 U485 ( .A1(n704), .A2(G478), .ZN(n597) );
  XOR2_X2 U486 ( .A(KEYINPUT40), .B(n530), .Z(n745) );
  XNOR2_X2 U487 ( .A(n421), .B(G472), .ZN(n675) );
  AND2_X1 U488 ( .A1(n558), .A2(n557), .ZN(n410) );
  NAND2_X1 U489 ( .A1(G221), .A2(n469), .ZN(n411) );
  INV_X1 U490 ( .A(KEYINPUT47), .ZN(n514) );
  XNOR2_X1 U491 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U492 ( .A(KEYINPUT10), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U494 ( .A(KEYINPUT71), .ZN(n564) );
  XNOR2_X1 U495 ( .A(n489), .B(n488), .ZN(n490) );
  INV_X1 U496 ( .A(n566), .ZN(n567) );
  INV_X1 U497 ( .A(KEYINPUT45), .ZN(n588) );
  BUF_X1 U498 ( .A(n657), .Z(n736) );
  INV_X1 U499 ( .A(n711), .ZN(n599) );
  INV_X1 U500 ( .A(KEYINPUT30), .ZN(n425) );
  NOR2_X2 U501 ( .A1(G953), .A2(G237), .ZN(n481) );
  NAND2_X1 U502 ( .A1(n481), .A2(G210), .ZN(n412) );
  XNOR2_X1 U503 ( .A(n412), .B(G137), .ZN(n414) );
  XOR2_X1 U504 ( .A(KEYINPUT73), .B(KEYINPUT5), .Z(n413) );
  XNOR2_X1 U505 ( .A(n414), .B(n413), .ZN(n418) );
  XNOR2_X2 U506 ( .A(G119), .B(G116), .ZN(n415) );
  XNOR2_X1 U507 ( .A(n415), .B(KEYINPUT3), .ZN(n417) );
  XNOR2_X1 U508 ( .A(G113), .B(KEYINPUT69), .ZN(n416) );
  XNOR2_X1 U509 ( .A(n417), .B(n416), .ZN(n497) );
  XNOR2_X1 U510 ( .A(n418), .B(n497), .ZN(n419) );
  XNOR2_X1 U511 ( .A(n448), .B(n419), .ZN(n420) );
  XNOR2_X1 U512 ( .A(n454), .B(n420), .ZN(n608) );
  INV_X1 U513 ( .A(G902), .ZN(n474) );
  NAND2_X1 U514 ( .A1(n608), .A2(n474), .ZN(n421) );
  INV_X1 U515 ( .A(n675), .ZN(n507) );
  XNOR2_X1 U516 ( .A(KEYINPUT72), .B(n409), .ZN(n500) );
  NAND2_X1 U517 ( .A1(n500), .A2(G214), .ZN(n423) );
  INV_X1 U518 ( .A(KEYINPUT92), .ZN(n422) );
  XNOR2_X1 U519 ( .A(n423), .B(n422), .ZN(n688) );
  NOR2_X1 U520 ( .A1(n507), .A2(n688), .ZN(n424) );
  XNOR2_X1 U521 ( .A(n425), .B(n424), .ZN(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n427) );
  XNOR2_X1 U523 ( .A(G128), .B(KEYINPUT77), .ZN(n426) );
  XNOR2_X1 U524 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U525 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n433) );
  NAND2_X1 U526 ( .A1(G234), .A2(n739), .ZN(n432) );
  XNOR2_X1 U527 ( .A(n433), .B(n432), .ZN(n469) );
  XOR2_X1 U528 ( .A(n449), .B(n477), .Z(n726) );
  NAND2_X1 U529 ( .A1(n614), .A2(n474), .ZN(n443) );
  XOR2_X1 U530 ( .A(KEYINPUT25), .B(KEYINPUT95), .Z(n439) );
  XNOR2_X1 U531 ( .A(KEYINPUT15), .B(G902), .ZN(n499) );
  NAND2_X1 U532 ( .A1(G234), .A2(n499), .ZN(n437) );
  XNOR2_X1 U533 ( .A(KEYINPUT20), .B(n437), .ZN(n444) );
  NAND2_X1 U534 ( .A1(n444), .A2(G217), .ZN(n438) );
  XNOR2_X1 U535 ( .A(n439), .B(n438), .ZN(n441) );
  INV_X1 U536 ( .A(KEYINPUT76), .ZN(n440) );
  XNOR2_X1 U537 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X2 U538 ( .A(n443), .B(n442), .ZN(n578) );
  INV_X1 U539 ( .A(n578), .ZN(n561) );
  AND2_X1 U540 ( .A1(n444), .A2(G221), .ZN(n446) );
  XNOR2_X1 U541 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n445) );
  XNOR2_X1 U542 ( .A(n446), .B(n445), .ZN(n666) );
  XOR2_X1 U543 ( .A(n449), .B(KEYINPUT78), .Z(n451) );
  NAND2_X1 U544 ( .A1(G227), .A2(n739), .ZN(n450) );
  XNOR2_X1 U545 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U546 ( .A(n495), .B(n452), .ZN(n453) );
  XNOR2_X1 U547 ( .A(n454), .B(n453), .ZN(n705) );
  OR2_X2 U548 ( .A1(n705), .A2(G902), .ZN(n456) );
  XNOR2_X2 U549 ( .A(n456), .B(n455), .ZN(n524) );
  XNOR2_X1 U550 ( .A(n457), .B(KEYINPUT14), .ZN(n552) );
  NAND2_X1 U551 ( .A1(G953), .A2(G902), .ZN(n548) );
  NOR2_X1 U552 ( .A1(G900), .A2(n548), .ZN(n458) );
  NAND2_X1 U553 ( .A1(n552), .A2(n458), .ZN(n459) );
  XNOR2_X1 U554 ( .A(n459), .B(KEYINPUT105), .ZN(n461) );
  INV_X1 U555 ( .A(n552), .ZN(n697) );
  NAND2_X1 U556 ( .A1(n739), .A2(G952), .ZN(n550) );
  NOR2_X1 U557 ( .A1(n697), .A2(n550), .ZN(n460) );
  NOR2_X1 U558 ( .A1(n461), .A2(n460), .ZN(n505) );
  XNOR2_X1 U559 ( .A(n462), .B(KEYINPUT75), .ZN(n463) );
  NOR2_X2 U560 ( .A1(n464), .A2(n463), .ZN(n527) );
  BUF_X1 U561 ( .A(n527), .Z(n492) );
  XOR2_X1 U562 ( .A(KEYINPUT7), .B(G122), .Z(n466) );
  XNOR2_X1 U563 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U564 ( .A(n468), .B(n467), .ZN(n473) );
  NAND2_X1 U565 ( .A1(G217), .A2(n469), .ZN(n471) );
  XOR2_X1 U566 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n470) );
  XNOR2_X1 U567 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U568 ( .A(n473), .B(n472), .ZN(n596) );
  NAND2_X1 U569 ( .A1(n596), .A2(n474), .ZN(n475) );
  XNOR2_X1 U570 ( .A(n475), .B(G478), .ZN(n533) );
  XNOR2_X1 U571 ( .A(n478), .B(KEYINPUT98), .ZN(n491) );
  XOR2_X1 U572 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n480) );
  XNOR2_X1 U573 ( .A(G140), .B(KEYINPUT12), .ZN(n479) );
  XNOR2_X1 U574 ( .A(n480), .B(n479), .ZN(n485) );
  XOR2_X1 U575 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n483) );
  NAND2_X1 U576 ( .A1(G214), .A2(n481), .ZN(n482) );
  XNOR2_X1 U577 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U578 ( .A(n485), .B(n484), .ZN(n489) );
  XNOR2_X1 U579 ( .A(G143), .B(G122), .ZN(n486) );
  XNOR2_X1 U580 ( .A(n487), .B(n486), .ZN(n488) );
  AND2_X1 U581 ( .A1(n533), .A2(n532), .ZN(n571) );
  NAND2_X1 U582 ( .A1(n492), .A2(n571), .ZN(n504) );
  XNOR2_X1 U583 ( .A(KEYINPUT16), .B(G122), .ZN(n496) );
  XNOR2_X1 U584 ( .A(n497), .B(n496), .ZN(n719) );
  INV_X1 U585 ( .A(n499), .ZN(n590) );
  AND2_X1 U586 ( .A1(n500), .A2(G210), .ZN(n502) );
  XNOR2_X1 U587 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n501) );
  XNOR2_X1 U588 ( .A(n502), .B(n501), .ZN(n503) );
  NOR2_X1 U589 ( .A1(n504), .A2(n511), .ZN(n643) );
  NOR2_X1 U590 ( .A1(n578), .A2(n505), .ZN(n506) );
  NAND2_X1 U591 ( .A1(n666), .A2(n506), .ZN(n520) );
  NOR2_X1 U592 ( .A1(n507), .A2(n520), .ZN(n508) );
  XOR2_X1 U593 ( .A(KEYINPUT28), .B(n508), .Z(n510) );
  XNOR2_X1 U594 ( .A(n524), .B(KEYINPUT106), .ZN(n509) );
  NOR2_X1 U595 ( .A1(n510), .A2(n509), .ZN(n538) );
  XNOR2_X1 U596 ( .A(n522), .B(KEYINPUT19), .ZN(n555) );
  NAND2_X1 U597 ( .A1(n538), .A2(n555), .ZN(n645) );
  INV_X1 U598 ( .A(n644), .ZN(n648) );
  AND2_X1 U599 ( .A1(n533), .A2(n513), .ZN(n651) );
  NOR2_X1 U600 ( .A1(n648), .A2(n651), .ZN(n683) );
  NOR2_X1 U601 ( .A1(n643), .A2(n516), .ZN(n517) );
  XNOR2_X1 U602 ( .A(n517), .B(KEYINPUT70), .ZN(n526) );
  INV_X1 U603 ( .A(KEYINPUT102), .ZN(n518) );
  XNOR2_X1 U604 ( .A(n518), .B(KEYINPUT6), .ZN(n519) );
  XNOR2_X1 U605 ( .A(n675), .B(n519), .ZN(n583) );
  NOR2_X1 U606 ( .A1(n644), .A2(n520), .ZN(n521) );
  NAND2_X1 U607 ( .A1(n583), .A2(n521), .ZN(n542) );
  XNOR2_X1 U608 ( .A(KEYINPUT107), .B(KEYINPUT36), .ZN(n523) );
  XNOR2_X2 U609 ( .A(n524), .B(KEYINPUT1), .ZN(n669) );
  XNOR2_X1 U610 ( .A(n742), .B(KEYINPUT83), .ZN(n525) );
  XNOR2_X1 U611 ( .A(n511), .B(KEYINPUT38), .ZN(n531) );
  NAND2_X1 U612 ( .A1(n527), .A2(n531), .ZN(n529) );
  XOR2_X1 U613 ( .A(KEYINPUT84), .B(KEYINPUT39), .Z(n528) );
  XNOR2_X1 U614 ( .A(n529), .B(n528), .ZN(n540) );
  NOR2_X2 U615 ( .A1(n540), .A2(n644), .ZN(n530) );
  INV_X1 U616 ( .A(n531), .ZN(n684) );
  OR2_X2 U617 ( .A1(n533), .A2(n532), .ZN(n535) );
  INV_X1 U618 ( .A(KEYINPUT103), .ZN(n534) );
  XNOR2_X1 U619 ( .A(n535), .B(n534), .ZN(n682) );
  INV_X1 U620 ( .A(n688), .ZN(n536) );
  NAND2_X1 U621 ( .A1(n689), .A2(n536), .ZN(n537) );
  NAND2_X1 U622 ( .A1(n679), .A2(n538), .ZN(n539) );
  XNOR2_X1 U623 ( .A(KEYINPUT42), .B(n539), .ZN(n744) );
  BUF_X1 U624 ( .A(n540), .Z(n541) );
  INV_X1 U625 ( .A(n651), .ZN(n639) );
  NOR2_X1 U626 ( .A1(n541), .A2(n639), .ZN(n655) );
  NOR2_X1 U627 ( .A1(n688), .A2(n542), .ZN(n543) );
  NAND2_X1 U628 ( .A1(n669), .A2(n543), .ZN(n544) );
  XNOR2_X1 U629 ( .A(KEYINPUT43), .B(n544), .ZN(n545) );
  AND2_X1 U630 ( .A1(n545), .A2(n511), .ZN(n603) );
  NOR2_X1 U631 ( .A1(n655), .A2(n603), .ZN(n546) );
  NAND2_X1 U632 ( .A1(n657), .A2(KEYINPUT2), .ZN(n547) );
  XNOR2_X1 U633 ( .A(n547), .B(KEYINPUT81), .ZN(n589) );
  XNOR2_X1 U634 ( .A(G898), .B(KEYINPUT93), .ZN(n717) );
  INV_X1 U635 ( .A(n548), .ZN(n549) );
  NAND2_X1 U636 ( .A1(n717), .A2(n549), .ZN(n551) );
  NAND2_X1 U637 ( .A1(n551), .A2(n550), .ZN(n553) );
  AND2_X1 U638 ( .A1(n553), .A2(n552), .ZN(n554) );
  OR2_X1 U639 ( .A1(n682), .A2(n408), .ZN(n556) );
  INV_X1 U640 ( .A(n583), .ZN(n558) );
  XNOR2_X1 U641 ( .A(n578), .B(KEYINPUT104), .ZN(n665) );
  NOR2_X1 U642 ( .A1(n665), .A2(n669), .ZN(n557) );
  XOR2_X1 U643 ( .A(KEYINPUT80), .B(KEYINPUT32), .Z(n559) );
  NAND2_X1 U644 ( .A1(n669), .A2(n561), .ZN(n562) );
  NOR2_X1 U645 ( .A1(n562), .A2(n675), .ZN(n563) );
  NAND2_X1 U646 ( .A1(n585), .A2(n563), .ZN(n605) );
  NAND2_X1 U647 ( .A1(n578), .A2(n666), .ZN(n668) );
  NAND2_X1 U648 ( .A1(n568), .A2(n567), .ZN(n570) );
  XNOR2_X1 U649 ( .A(KEYINPUT79), .B(KEYINPUT34), .ZN(n569) );
  XNOR2_X1 U650 ( .A(n570), .B(n569), .ZN(n572) );
  NAND2_X1 U651 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X2 U652 ( .A(n573), .B(KEYINPUT35), .ZN(n607) );
  NAND2_X1 U653 ( .A1(n359), .A2(KEYINPUT44), .ZN(n574) );
  NAND2_X1 U654 ( .A1(n575), .A2(n675), .ZN(n664) );
  NOR2_X1 U655 ( .A1(n566), .A2(n664), .ZN(n576) );
  XOR2_X1 U656 ( .A(KEYINPUT31), .B(n576), .Z(n652) );
  NAND2_X1 U657 ( .A1(n578), .A2(n577), .ZN(n579) );
  OR2_X1 U658 ( .A1(n675), .A2(n579), .ZN(n580) );
  NOR2_X1 U659 ( .A1(n652), .A2(n357), .ZN(n581) );
  NOR2_X1 U660 ( .A1(n581), .A2(n683), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n665), .A2(n669), .ZN(n582) );
  NOR2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U663 ( .A1(n585), .A2(n584), .ZN(n632) );
  NOR2_X1 U664 ( .A1(n586), .A2(n632), .ZN(n587) );
  INV_X1 U665 ( .A(n712), .ZN(n658) );
  INV_X1 U666 ( .A(KEYINPUT74), .ZN(n591) );
  XNOR2_X1 U667 ( .A(n591), .B(n657), .ZN(n592) );
  NOR2_X1 U668 ( .A1(n712), .A2(n592), .ZN(n593) );
  NOR2_X1 U669 ( .A1(n593), .A2(KEYINPUT2), .ZN(n594) );
  NOR2_X4 U670 ( .A1(n595), .A2(n594), .ZN(n704) );
  INV_X1 U671 ( .A(G952), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n602) );
  INV_X1 U673 ( .A(KEYINPUT120), .ZN(n601) );
  XNOR2_X1 U674 ( .A(n602), .B(n601), .ZN(G63) );
  XOR2_X1 U675 ( .A(n603), .B(G140), .Z(G42) );
  XOR2_X1 U676 ( .A(G110), .B(KEYINPUT111), .Z(n604) );
  XNOR2_X1 U677 ( .A(n605), .B(n604), .ZN(G12) );
  XNOR2_X1 U678 ( .A(n606), .B(G119), .ZN(G21) );
  XOR2_X1 U679 ( .A(n607), .B(G122), .Z(G24) );
  NAND2_X1 U680 ( .A1(n704), .A2(G472), .ZN(n610) );
  XOR2_X1 U681 ( .A(KEYINPUT62), .B(n608), .Z(n609) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(n611) );
  NOR2_X2 U683 ( .A1(n611), .A2(n711), .ZN(n613) );
  XNOR2_X1 U684 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n613), .B(n612), .ZN(G57) );
  NAND2_X1 U686 ( .A1(n704), .A2(G217), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n614), .B(KEYINPUT121), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(n617) );
  NOR2_X2 U689 ( .A1(n617), .A2(n711), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n618), .B(KEYINPUT122), .ZN(G66) );
  NAND2_X1 U691 ( .A1(n704), .A2(G475), .ZN(n623) );
  XOR2_X1 U692 ( .A(KEYINPUT64), .B(KEYINPUT88), .Z(n619) );
  XNOR2_X1 U693 ( .A(n619), .B(KEYINPUT59), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X2 U696 ( .A1(n624), .A2(n711), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n625), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U698 ( .A1(n704), .A2(G210), .ZN(n629) );
  XOR2_X1 U699 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n626) );
  XNOR2_X1 U700 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(n630) );
  NOR2_X2 U702 ( .A1(n630), .A2(n711), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n631), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U704 ( .A(G101), .B(n632), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n633), .B(KEYINPUT109), .ZN(G3) );
  NAND2_X1 U706 ( .A1(n357), .A2(n648), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n634), .B(KEYINPUT110), .ZN(n635) );
  XNOR2_X1 U708 ( .A(G104), .B(n635), .ZN(G6) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n637) );
  NAND2_X1 U710 ( .A1(n357), .A2(n651), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U712 ( .A(G107), .B(n638), .ZN(G9) );
  NOR2_X1 U713 ( .A1(n645), .A2(n639), .ZN(n641) );
  XNOR2_X1 U714 ( .A(KEYINPUT112), .B(KEYINPUT29), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U716 ( .A(G128), .B(n642), .ZN(G30) );
  XOR2_X1 U717 ( .A(G143), .B(n643), .Z(G45) );
  NOR2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n647) );
  XNOR2_X1 U719 ( .A(G146), .B(KEYINPUT113), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(G48) );
  NAND2_X1 U721 ( .A1(n652), .A2(n648), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n649), .B(KEYINPUT114), .ZN(n650) );
  XNOR2_X1 U723 ( .A(G113), .B(n650), .ZN(G15) );
  XOR2_X1 U724 ( .A(G116), .B(KEYINPUT115), .Z(n654) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n654), .B(n653), .ZN(G18) );
  XOR2_X1 U727 ( .A(G134), .B(n655), .Z(n656) );
  XNOR2_X1 U728 ( .A(KEYINPUT116), .B(n656), .ZN(G36) );
  NAND2_X1 U729 ( .A1(n658), .A2(n736), .ZN(n660) );
  INV_X1 U730 ( .A(KEYINPUT2), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U733 ( .A1(n663), .A2(n739), .ZN(n702) );
  NAND2_X1 U734 ( .A1(n679), .A2(n568), .ZN(n700) );
  INV_X1 U735 ( .A(n664), .ZN(n677) );
  NOR2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U737 ( .A(KEYINPUT49), .B(n667), .ZN(n673) );
  XOR2_X1 U738 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n671) );
  NAND2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U744 ( .A(KEYINPUT51), .B(n678), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U746 ( .A(KEYINPUT118), .B(n681), .Z(n694) );
  INV_X1 U747 ( .A(n682), .ZN(n686) );
  NOR2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n690) );
  NOR2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U752 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U753 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U754 ( .A(n695), .B(KEYINPUT52), .ZN(n696) );
  NOR2_X1 U755 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U756 ( .A1(n698), .A2(G952), .ZN(n699) );
  NAND2_X1 U757 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U758 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U759 ( .A(n703), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U760 ( .A1(n704), .A2(G469), .ZN(n709) );
  XNOR2_X1 U761 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n705), .B(KEYINPUT57), .ZN(n706) );
  XNOR2_X1 U763 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n711), .A2(n710), .ZN(G54) );
  NOR2_X1 U766 ( .A1(n712), .A2(G953), .ZN(n716) );
  NAND2_X1 U767 ( .A1(G953), .A2(G224), .ZN(n713) );
  XOR2_X1 U768 ( .A(KEYINPUT61), .B(n713), .Z(n714) );
  NOR2_X1 U769 ( .A1(n717), .A2(n714), .ZN(n715) );
  NOR2_X1 U770 ( .A1(n716), .A2(n715), .ZN(n725) );
  NAND2_X1 U771 ( .A1(n717), .A2(G953), .ZN(n722) );
  XOR2_X1 U772 ( .A(n718), .B(G101), .Z(n720) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U774 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n723), .B(KEYINPUT123), .ZN(n724) );
  XOR2_X1 U776 ( .A(n725), .B(n724), .Z(G69) );
  XNOR2_X1 U777 ( .A(n726), .B(KEYINPUT124), .ZN(n730) );
  XNOR2_X1 U778 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(n735) );
  INV_X1 U780 ( .A(n735), .ZN(n731) );
  XNOR2_X1 U781 ( .A(G227), .B(n731), .ZN(n732) );
  NAND2_X1 U782 ( .A1(n732), .A2(G900), .ZN(n733) );
  XNOR2_X1 U783 ( .A(n733), .B(KEYINPUT126), .ZN(n734) );
  NAND2_X1 U784 ( .A1(n734), .A2(G953), .ZN(n741) );
  XNOR2_X1 U785 ( .A(n735), .B(KEYINPUT125), .ZN(n737) );
  XOR2_X1 U786 ( .A(n737), .B(n736), .Z(n738) );
  NAND2_X1 U787 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n741), .A2(n740), .ZN(G72) );
  XNOR2_X1 U789 ( .A(G125), .B(KEYINPUT37), .ZN(n743) );
  XNOR2_X1 U790 ( .A(n743), .B(n742), .ZN(G27) );
  XNOR2_X1 U791 ( .A(G137), .B(n744), .ZN(G39) );
  XOR2_X1 U792 ( .A(n745), .B(G131), .Z(n746) );
  XNOR2_X1 U793 ( .A(KEYINPUT127), .B(n746), .ZN(G33) );
endmodule

