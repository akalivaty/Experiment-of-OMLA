//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(new_n189), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G227), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G953), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n193), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(G137), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT11), .A3(G134), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n200), .A2(new_n203), .A3(new_n206), .A4(new_n201), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT10), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n215), .A2(KEYINPUT1), .A3(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT65), .A2(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT65), .A2(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n220), .A2(new_n221), .B1(new_n212), .B2(new_n214), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT73), .ZN(new_n225));
  INV_X1    g039(.A(G107), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G104), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT73), .A3(G107), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(G107), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT72), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT3), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n232), .A2(new_n226), .A3(KEYINPUT3), .A4(G104), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n224), .B(new_n230), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT75), .B1(new_n228), .B2(G107), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT75), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n226), .A3(G104), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n228), .A2(G107), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G101), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n236), .A2(KEYINPUT76), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT76), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n244), .A3(G101), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n210), .B(new_n223), .C1(new_n243), .C2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n230), .B1(new_n233), .B2(new_n235), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT74), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n232), .A2(new_n226), .A3(G104), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n234), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT74), .A3(new_n230), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(G101), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n252), .A2(new_n234), .B1(new_n227), .B2(new_n229), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(new_n224), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n249), .A2(KEYINPUT4), .A3(G101), .A4(new_n254), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n215), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n264), .ZN(new_n266));
  NOR2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n215), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n246), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n245), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n244), .B1(new_n257), .B2(new_n224), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(new_n242), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n221), .A2(G128), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n217), .B1(new_n215), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n210), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n209), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n269), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n260), .B2(new_n261), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n275), .B1(new_n243), .B2(new_n245), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(KEYINPUT10), .ZN(new_n281));
  NOR4_X1   g095(.A1(new_n279), .A2(new_n281), .A3(new_n246), .A4(new_n208), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n197), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n243), .A2(new_n245), .A3(new_n223), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n208), .B1(new_n284), .B2(new_n280), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT12), .B(new_n208), .C1(new_n284), .C2(new_n280), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n262), .A2(new_n269), .ZN(new_n290));
  INV_X1    g104(.A(new_n246), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n290), .A2(new_n209), .A3(new_n276), .A4(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n292), .A3(new_n196), .ZN(new_n293));
  AOI21_X1  g107(.A(G902), .B1(new_n283), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n192), .B1(new_n294), .B2(new_n191), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n296));
  INV_X1    g110(.A(new_n288), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n243), .A2(new_n245), .A3(new_n223), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n298), .B1(new_n273), .B2(new_n275), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT12), .B1(new_n299), .B2(new_n208), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n296), .B1(new_n301), .B2(new_n282), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n289), .A2(new_n292), .A3(KEYINPUT77), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(new_n197), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n277), .A2(new_n282), .A3(new_n197), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n306), .A3(G469), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n190), .B1(new_n295), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G214), .B1(G237), .B2(G902), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT67), .B(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n269), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(new_n310), .B2(new_n223), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT80), .B(G224), .ZN(new_n313));
  INV_X1    g127(.A(G953), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n312), .B(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT2), .B(G113), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G116), .B(G119), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n319), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n317), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI221_X4 g137(.A(new_n248), .B1(new_n227), .B2(new_n229), .C1(new_n252), .C2(new_n234), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT74), .B1(new_n253), .B2(new_n230), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n258), .B1(new_n326), .B2(G101), .ZN(new_n327));
  INV_X1    g141(.A(new_n261), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n331));
  INV_X1    g145(.A(G119), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G116), .ZN(new_n333));
  OAI211_X1 g147(.A(G113), .B(new_n333), .C1(new_n321), .C2(new_n331), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n320), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n273), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n329), .A2(new_n330), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n323), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n339), .B1(new_n260), .B2(new_n261), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT78), .B1(new_n340), .B2(new_n336), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(G110), .B(G122), .Z(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n343), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n329), .A2(new_n345), .A3(new_n337), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(KEYINPUT6), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n349));
  AND4_X1   g163(.A1(new_n348), .A2(new_n342), .A3(new_n349), .A4(new_n343), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n345), .B1(new_n338), .B2(new_n341), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n348), .B1(new_n351), .B2(new_n349), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n316), .B(new_n347), .C1(new_n350), .C2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(G210), .B1(G237), .B2(G902), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT81), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT7), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n315), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n316), .B(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n343), .B(KEYINPUT8), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n273), .A2(new_n335), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n337), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(G902), .B1(new_n363), .B2(new_n346), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n353), .A2(new_n356), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n356), .B1(new_n353), .B2(new_n364), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n308), .B(new_n309), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT16), .ZN(new_n368));
  INV_X1    g182(.A(G140), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n310), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G125), .A2(G140), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n310), .B2(G140), .ZN(new_n372));
  OAI211_X1 g186(.A(G146), .B(new_n370), .C1(new_n372), .C2(new_n368), .ZN(new_n373));
  XNOR2_X1  g187(.A(G125), .B(G140), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n211), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n332), .A2(KEYINPUT23), .A3(G128), .ZN(new_n376));
  MUX2_X1   g190(.A(new_n216), .B(new_n220), .S(G119), .Z(new_n377));
  AOI21_X1  g191(.A(new_n376), .B1(new_n377), .B2(KEYINPUT23), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(G110), .ZN(new_n379));
  XOR2_X1   g193(.A(KEYINPUT24), .B(G110), .Z(new_n380));
  NOR2_X1   g194(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n373), .B(new_n375), .C1(new_n379), .C2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT70), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n373), .B(KEYINPUT68), .ZN(new_n384));
  INV_X1    g198(.A(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT67), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT67), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G125), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n388), .A3(G140), .ZN(new_n389));
  INV_X1    g203(.A(new_n371), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n368), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND4_X1   g205(.A1(new_n368), .A2(new_n386), .A3(new_n388), .A4(new_n369), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n211), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT69), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(KEYINPUT69), .B(new_n211), .C1(new_n391), .C2(new_n392), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n384), .A2(new_n397), .B1(G110), .B2(new_n378), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n377), .A2(new_n380), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n383), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT68), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n373), .A2(new_n401), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n373), .A2(new_n401), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n397), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n378), .A2(G110), .ZN(new_n405));
  AND4_X1   g219(.A1(new_n383), .A2(new_n404), .A3(new_n399), .A4(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n382), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n314), .A2(G221), .A3(G234), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT22), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(G137), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n382), .B(new_n410), .C1(new_n400), .C2(new_n406), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n189), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT25), .ZN(new_n415));
  INV_X1    g229(.A(G217), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(G234), .B2(new_n189), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT25), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n412), .A2(new_n418), .A3(new_n189), .A4(new_n413), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n415), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n269), .A2(new_n208), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n202), .A2(G134), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n201), .A2(new_n422), .A3(KEYINPUT64), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(G131), .C1(KEYINPUT64), .C2(new_n422), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n424), .B(new_n207), .C1(new_n217), .C2(new_n222), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n427), .A2(KEYINPUT66), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(KEYINPUT66), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n421), .A2(new_n425), .A3(KEYINPUT66), .A4(new_n427), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n339), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n421), .A2(new_n425), .A3(new_n339), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT31), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(G101), .ZN(new_n437));
  INV_X1    g251(.A(G237), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n314), .A3(G210), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n437), .B(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n434), .A2(new_n435), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n339), .B1(new_n421), .B2(new_n425), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT28), .B1(new_n433), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n421), .A2(new_n425), .A3(new_n339), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT28), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n440), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT31), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n432), .A2(new_n433), .A3(new_n448), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n441), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT32), .ZN(new_n452));
  NOR2_X1   g266(.A1(G472), .A2(G902), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n451), .B2(new_n453), .ZN(new_n455));
  INV_X1    g269(.A(G472), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n443), .A2(KEYINPUT29), .A3(new_n440), .A4(new_n446), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n434), .A2(new_n440), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n447), .B2(new_n448), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n457), .B(new_n189), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  OAI22_X1  g276(.A1(new_n454), .A2(new_n455), .B1(new_n456), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n412), .A2(new_n413), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n417), .A2(G902), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT71), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n420), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n470));
  INV_X1    g284(.A(G116), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT14), .A3(G122), .ZN(new_n472));
  XNOR2_X1  g286(.A(G116), .B(G122), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(G107), .B(new_n472), .C1(new_n474), .C2(KEYINPUT14), .ZN(new_n475));
  OAI21_X1  g289(.A(G143), .B1(new_n218), .B2(new_n219), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n213), .A2(G128), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n199), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n473), .A2(new_n226), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(G134), .A3(new_n477), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n475), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n473), .B(new_n226), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT85), .B(KEYINPUT13), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n476), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n486), .A2(G134), .B1(new_n477), .B2(new_n476), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT85), .B(KEYINPUT13), .Z(new_n488));
  AND4_X1   g302(.A1(G134), .A2(new_n488), .A3(new_n476), .A4(new_n477), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n484), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(KEYINPUT86), .B(new_n484), .C1(new_n487), .C2(new_n489), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n483), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n188), .A2(G217), .A3(new_n314), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n470), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n496), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n500));
  INV_X1    g314(.A(G478), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(KEYINPUT15), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n499), .A2(new_n500), .A3(new_n189), .A4(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n492), .A2(new_n493), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n495), .B1(new_n505), .B2(new_n483), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n470), .A3(new_n498), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(KEYINPUT87), .A3(new_n496), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n500), .A4(new_n189), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n502), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(G234), .A2(G237), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n513), .A2(G952), .A3(new_n314), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(G902), .A3(G953), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n516), .B(KEYINPUT89), .Z(new_n517));
  XOR2_X1   g331(.A(KEYINPUT21), .B(G898), .Z(new_n518));
  OAI21_X1  g332(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n438), .A2(new_n314), .A3(G214), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n213), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n438), .A2(new_n314), .A3(G143), .A4(G214), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(KEYINPUT18), .A2(G131), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n372), .A2(G146), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n375), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT82), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n526), .A2(KEYINPUT82), .A3(new_n528), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(G113), .B(G122), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(G104), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT83), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n524), .A2(KEYINPUT17), .A3(G131), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n397), .A2(new_n402), .A3(new_n403), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n524), .A2(G131), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n522), .A2(new_n206), .A3(new_n523), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT84), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n533), .B(new_n536), .C1(new_n538), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n539), .A2(new_n541), .ZN(new_n546));
  MUX2_X1   g360(.A(new_n374), .B(new_n372), .S(KEYINPUT19), .Z(new_n547));
  OAI211_X1 g361(.A(new_n373), .B(new_n546), .C1(new_n547), .C2(G146), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n526), .A2(KEYINPUT82), .A3(new_n528), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT82), .B1(new_n526), .B2(new_n528), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n535), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(G475), .A2(G902), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n520), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  AOI211_X1 g370(.A(KEYINPUT20), .B(new_n556), .C1(new_n545), .C2(new_n552), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n533), .B1(new_n538), .B2(new_n544), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n535), .ZN(new_n559));
  AOI21_X1  g373(.A(G902), .B1(new_n559), .B2(new_n545), .ZN(new_n560));
  INV_X1    g374(.A(G475), .ZN(new_n561));
  OAI22_X1  g375(.A1(new_n555), .A2(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n512), .A2(new_n519), .A3(new_n563), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n367), .A2(new_n469), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(new_n224), .ZN(G3));
  AND2_X1   g380(.A1(new_n420), .A2(new_n468), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT90), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n456), .B1(new_n451), .B2(new_n189), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n451), .B2(new_n453), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n567), .A2(new_n568), .A3(new_n308), .A4(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n308), .A2(new_n468), .A3(new_n420), .A4(new_n570), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT90), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n309), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n353), .A2(new_n364), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n355), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n353), .A2(new_n356), .A3(new_n364), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n507), .A2(new_n580), .A3(new_n508), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n506), .A2(KEYINPUT33), .A3(new_n498), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n581), .A2(G478), .A3(new_n189), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n507), .A2(new_n189), .A3(new_n508), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n501), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n562), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n579), .A2(new_n519), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n574), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT34), .B(G104), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  XNOR2_X1  g406(.A(new_n572), .B(new_n568), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n519), .B(new_n309), .C1(new_n365), .C2(new_n366), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n560), .A2(new_n561), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n504), .B2(new_n510), .ZN(new_n597));
  AND4_X1   g411(.A1(KEYINPUT91), .A2(new_n553), .A3(new_n520), .A4(new_n554), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n555), .A2(new_n557), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n593), .A2(new_n595), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G107), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  INV_X1    g419(.A(new_n367), .ZN(new_n606));
  INV_X1    g420(.A(new_n564), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n411), .A2(KEYINPUT36), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n407), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n407), .A2(new_n609), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n467), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n420), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n606), .A2(new_n607), .A3(new_n570), .A4(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT37), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G110), .ZN(G12));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n617));
  INV_X1    g431(.A(new_n517), .ZN(new_n618));
  INV_X1    g432(.A(G900), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n514), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT92), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n597), .A2(new_n601), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT93), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT93), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n597), .A2(new_n601), .A3(new_n625), .A4(new_n622), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n309), .B1(new_n365), .B2(new_n366), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n617), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n613), .A2(new_n463), .A3(new_n308), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n579), .A2(KEYINPUT94), .A3(new_n626), .A4(new_n624), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G128), .ZN(G30));
  NOR4_X1   g448(.A1(new_n613), .A2(new_n512), .A3(new_n563), .A4(new_n575), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT97), .Z(new_n636));
  NAND2_X1  g450(.A1(new_n577), .A2(new_n578), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n621), .B(KEYINPUT39), .Z(new_n641));
  NAND2_X1  g455(.A1(new_n308), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT40), .ZN(new_n643));
  NOR4_X1   g457(.A1(new_n432), .A2(KEYINPUT31), .A3(new_n433), .A4(new_n448), .ZN(new_n644));
  INV_X1    g458(.A(new_n449), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n430), .A2(new_n431), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n323), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n444), .A3(new_n440), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n644), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n453), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT32), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT95), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n448), .B1(new_n433), .B2(new_n442), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n648), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n189), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n654), .B1(new_n648), .B2(new_n655), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT96), .B1(new_n653), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n659), .B(KEYINPUT96), .C1(new_n454), .C2(new_n455), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n643), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n636), .A2(new_n640), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  NAND3_X1  g480(.A1(new_n586), .A2(new_n562), .A3(new_n622), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n630), .A2(new_n628), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n211), .ZN(G48));
  NOR2_X1   g483(.A1(new_n594), .A2(new_n587), .ZN(new_n670));
  INV_X1    g484(.A(new_n190), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n290), .A2(new_n276), .A3(new_n291), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n208), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n196), .B1(new_n673), .B2(new_n292), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n289), .A2(new_n292), .A3(new_n196), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n191), .B(new_n189), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n294), .A2(new_n191), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n294), .A2(new_n677), .A3(new_n191), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n671), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n469), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n670), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT99), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n684), .B(new_n686), .ZN(G15));
  NAND3_X1  g501(.A1(new_n595), .A2(new_n683), .A3(new_n602), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT100), .B(G116), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G18));
  OAI21_X1  g504(.A(KEYINPUT101), .B1(new_n628), .B2(new_n682), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n189), .B1(new_n674), .B2(new_n675), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n677), .A3(new_n676), .ZN(new_n694));
  INV_X1    g508(.A(new_n681), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n190), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT101), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n637), .A2(new_n696), .A3(new_n697), .A4(new_n309), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n613), .A2(new_n463), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n699), .A2(new_n607), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  OAI21_X1  g517(.A(G472), .B1(new_n649), .B2(G902), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n645), .A2(KEYINPUT102), .A3(new_n648), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n705), .B(new_n453), .C1(new_n451), .C2(KEYINPUT102), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n420), .A2(new_n707), .A3(new_n468), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n594), .A2(new_n682), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n710), .B1(new_n512), .B2(new_n563), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n511), .A2(KEYINPUT103), .A3(new_n562), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  INV_X1    g530(.A(new_n667), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n613), .A2(new_n717), .A3(new_n707), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n628), .A2(new_n682), .A3(KEYINPUT101), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n697), .B1(new_n579), .B2(new_n696), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  NOR2_X1   g536(.A1(new_n190), .A2(new_n575), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n365), .A2(new_n366), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n420), .A2(new_n463), .A3(new_n468), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n307), .A2(KEYINPUT104), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n304), .A2(new_n306), .A3(new_n728), .A4(G469), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n295), .A3(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n725), .A2(new_n726), .A3(new_n717), .A4(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT106), .B1(new_n732), .B2(KEYINPUT105), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n577), .A2(new_n730), .A3(new_n578), .A4(new_n723), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n733), .B1(KEYINPUT106), .B2(new_n732), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n726), .A3(new_n717), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G131), .ZN(G33));
  NAND4_X1  g555(.A1(new_n736), .A2(new_n726), .A3(new_n626), .A4(new_n624), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NOR2_X1   g557(.A1(new_n637), .A2(new_n575), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT107), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n562), .B1(new_n585), .B2(new_n583), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n746), .A2(KEYINPUT43), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(KEYINPUT43), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n570), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n613), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n745), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n289), .A2(new_n292), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n196), .B1(new_n757), .B2(new_n296), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n305), .B1(new_n758), .B2(new_n303), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(KEYINPUT45), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(KEYINPUT45), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(G469), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n192), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n763), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n676), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(new_n671), .A3(new_n641), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n745), .A2(new_n753), .A3(new_n770), .A4(new_n754), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n756), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  INV_X1    g587(.A(new_n567), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n463), .A2(new_n667), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n744), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT109), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n768), .A2(new_n671), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT47), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n768), .A2(KEYINPUT47), .A3(new_n671), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n777), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  NAND2_X1  g599(.A1(new_n694), .A2(new_n695), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n190), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n780), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n515), .B(new_n708), .C1(new_n747), .C2(new_n748), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n788), .A2(new_n745), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n637), .A2(new_n638), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT38), .B1(new_n577), .B2(new_n578), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n575), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n682), .A2(new_n708), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n515), .B1(new_n747), .B2(new_n748), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT50), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n725), .A2(new_n786), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n613), .A3(new_n707), .A4(new_n795), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n793), .A2(new_n796), .A3(KEYINPUT50), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n725), .A2(new_n567), .A3(new_n786), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n663), .A2(new_n514), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT112), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT112), .B1(new_n803), .B2(new_n804), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n586), .A2(new_n562), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n790), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(G952), .B(new_n314), .C1(new_n810), .C2(KEYINPUT51), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n788), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n780), .A2(KEYINPUT114), .A3(new_n782), .A4(new_n787), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n745), .A3(new_n789), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n802), .A2(new_n816), .A3(new_n808), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n802), .B2(new_n808), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n815), .B(KEYINPUT51), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n809), .A2(KEYINPUT113), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n802), .A2(new_n816), .A3(new_n808), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT51), .A4(new_n815), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n811), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n798), .A2(new_n726), .A3(new_n795), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT48), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n699), .A2(new_n789), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n597), .B1(new_n555), .B2(new_n557), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n571), .A2(new_n595), .A3(new_n573), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n614), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(KEYINPUT110), .A3(new_n614), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n565), .B1(new_n593), .B2(new_n670), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n709), .A2(new_n714), .B1(new_n670), .B2(new_n683), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n702), .A3(new_n688), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n718), .A2(new_n736), .A3(KEYINPUT111), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n613), .A2(new_n717), .A3(new_n707), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n730), .A2(new_n577), .A3(new_n578), .A4(new_n723), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n622), .B1(new_n560), .B2(new_n561), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n630), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n512), .A3(new_n601), .A4(new_n744), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n740), .A2(new_n847), .A3(new_n742), .A4(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n838), .A2(new_n841), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n668), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n730), .A2(new_n420), .A3(new_n612), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n663), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n628), .A2(new_n713), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n856), .A3(new_n671), .A4(new_n622), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n721), .A2(new_n633), .A3(new_n853), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT52), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n668), .B1(new_n699), .B2(new_n718), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n861), .A3(new_n633), .A4(new_n857), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT53), .B1(new_n852), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n606), .A2(new_n726), .A3(new_n607), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n688), .B(new_n865), .C1(new_n574), .C2(new_n589), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n564), .B(new_n700), .C1(new_n691), .C2(new_n698), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n595), .A2(new_n794), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n726), .A2(new_n696), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n868), .A2(new_n713), .B1(new_n589), .B2(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n866), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n833), .A2(KEYINPUT110), .A3(new_n614), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT110), .B1(new_n833), .B2(new_n614), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n740), .A2(new_n742), .A3(new_n847), .A4(new_n850), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n859), .A2(new_n862), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n830), .B1(new_n864), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n852), .A2(new_n863), .A3(KEYINPUT53), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n878), .B1(new_n876), .B2(new_n877), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT54), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n826), .A2(new_n828), .A3(new_n829), .A4(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n805), .A2(new_n588), .A3(new_n806), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n885), .A2(new_n886), .B1(G952), .B2(G953), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT49), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n662), .B(new_n660), .C1(new_n888), .C2(new_n786), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n694), .A2(new_n695), .A3(KEYINPUT49), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n890), .A2(new_n723), .A3(new_n746), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n639), .A2(new_n889), .A3(new_n567), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n892), .ZN(G75));
  AOI21_X1  g707(.A(new_n189), .B1(new_n881), .B2(new_n882), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT56), .B1(new_n894), .B2(new_n355), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n347), .B1(new_n350), .B2(new_n352), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n316), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT55), .ZN(new_n898));
  OR3_X1    g712(.A1(new_n895), .A2(KEYINPUT116), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n314), .A2(G952), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n895), .B2(KEYINPUT116), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n898), .B1(new_n895), .B2(KEYINPUT116), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(G51));
  XNOR2_X1  g717(.A(new_n192), .B(KEYINPUT117), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT57), .Z(new_n905));
  NAND3_X1  g719(.A1(new_n880), .A2(new_n883), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n283), .A2(new_n293), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n894), .A2(G469), .A3(new_n760), .A4(new_n761), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n900), .B1(new_n911), .B2(new_n912), .ZN(G54));
  NAND3_X1  g727(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .ZN(new_n914));
  INV_X1    g728(.A(new_n553), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n917), .A3(new_n900), .ZN(G60));
  NAND2_X1  g732(.A1(new_n581), .A2(new_n582), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT119), .Z(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT59), .ZN(new_n922));
  OR3_X1    g736(.A1(new_n884), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n900), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n919), .B1(new_n884), .B2(new_n922), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G63));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n610), .A2(new_n611), .ZN(new_n928));
  XNOR2_X1  g742(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n416), .A2(new_n189), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n928), .B(new_n932), .C1(new_n881), .C2(new_n882), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n927), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n881), .A2(new_n882), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n931), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n900), .B1(new_n938), .B2(new_n464), .ZN(new_n939));
  INV_X1    g753(.A(new_n933), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n932), .B1(new_n881), .B2(new_n882), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n924), .B1(new_n942), .B2(new_n465), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n943), .A2(KEYINPUT122), .A3(new_n933), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n935), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n939), .A2(new_n936), .A3(new_n940), .ZN(new_n946));
  INV_X1    g760(.A(new_n935), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT122), .B1(new_n943), .B2(new_n933), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n945), .A2(new_n949), .ZN(G66));
  AOI21_X1  g764(.A(new_n314), .B1(new_n518), .B2(new_n313), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n871), .A2(new_n874), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n314), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n896), .B1(G898), .B2(new_n314), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n953), .B(new_n954), .Z(G69));
  XNOR2_X1  g769(.A(new_n547), .B(KEYINPUT123), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n646), .B(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT124), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n772), .A2(new_n784), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n469), .B1(new_n587), .B2(new_n831), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n308), .A3(new_n744), .A4(new_n641), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n860), .A2(new_n633), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT62), .B1(new_n665), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n665), .A2(new_n962), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n959), .B(new_n961), .C1(new_n963), .C2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n958), .B1(new_n967), .B2(new_n314), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n769), .A2(new_n726), .A3(new_n856), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n969), .A2(new_n740), .A3(new_n742), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n959), .A2(new_n962), .A3(new_n970), .ZN(new_n971));
  MUX2_X1   g785(.A(new_n619), .B(new_n971), .S(new_n314), .Z(new_n972));
  AOI21_X1  g786(.A(new_n968), .B1(new_n972), .B2(new_n957), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n194), .B2(new_n619), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT125), .Z(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n967), .B2(new_n952), .ZN(new_n979));
  INV_X1    g793(.A(new_n434), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n980), .A3(new_n440), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n978), .B1(new_n971), .B2(new_n952), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n982), .A2(new_n434), .A3(new_n448), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n977), .B1(new_n458), .B2(new_n450), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT126), .Z(new_n985));
  AOI21_X1  g799(.A(new_n900), .B1(new_n937), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n981), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n981), .A2(new_n983), .A3(KEYINPUT127), .A4(new_n986), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G57));
endmodule


