//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G97), .A2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G68), .A2(G238), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n214), .B(new_n218), .C1(G58), .C2(G232), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G1), .B2(G20), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n207), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n210), .B(new_n221), .C1(new_n223), .C2(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G244), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT64), .B(KEYINPUT2), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT65), .B(G238), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n217), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G97), .B(G107), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G87), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n216), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(KEYINPUT13), .ZN(new_n244));
  INV_X1    g0044(.A(G1698), .ZN(new_n245));
  AND2_X1   g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  OAI211_X1 g0047(.A(G226), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  OAI211_X1 g0048(.A(G232), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G97), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G238), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AND4_X1   g0061(.A1(new_n244), .A2(new_n255), .A3(new_n258), .A4(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n251), .B2(new_n254), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n244), .B1(new_n263), .B2(new_n258), .ZN(new_n264));
  OAI21_X1  g0064(.A(G169), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT14), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n262), .A2(new_n264), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G179), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT14), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n269), .B(G169), .C1(new_n262), .C2(new_n264), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT75), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT75), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n266), .A2(new_n268), .A3(new_n273), .A4(new_n270), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT70), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT70), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(new_n206), .A3(G13), .A4(G20), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n206), .A2(G20), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n222), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n280), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G68), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT12), .B1(new_n280), .B2(G68), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT74), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(G20), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  OR4_X1    g0091(.A1(KEYINPUT12), .A2(new_n290), .A3(G1), .A4(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n287), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n207), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G77), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n290), .B1(new_n294), .B2(new_n295), .C1(new_n297), .C2(new_n202), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n283), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n299), .B(KEYINPUT11), .Z(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n275), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n267), .A2(G190), .ZN(new_n305));
  OAI21_X1  g0105(.A(G200), .B1(new_n262), .B2(new_n264), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT68), .ZN(new_n309));
  OAI21_X1  g0109(.A(G1698), .B1(new_n246), .B2(new_n247), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT66), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(KEYINPUT66), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(G238), .A3(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n246), .A2(new_n247), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G232), .ZN(new_n317));
  AND2_X1   g0117(.A1(KEYINPUT67), .A2(G107), .ZN(new_n318));
  NOR2_X1   g0118(.A1(KEYINPUT67), .A2(G107), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n315), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n314), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n254), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n260), .B1(new_n257), .B2(G244), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n309), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n324), .ZN(new_n326));
  AOI211_X1 g0126(.A(KEYINPUT68), .B(new_n326), .C1(new_n322), .C2(new_n254), .ZN(new_n327));
  OAI21_X1  g0127(.A(G190), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT69), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g0130(.A(KEYINPUT69), .B(G190), .C1(new_n325), .C2(new_n327), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n285), .A2(new_n295), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT8), .B(G58), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n335), .A2(new_n296), .B1(G20), .B2(G77), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT15), .B(G87), .Z(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n336), .B1(new_n294), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n333), .B1(new_n283), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n277), .A2(new_n279), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n295), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n325), .A2(new_n327), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n332), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n325), .A2(new_n327), .A3(G169), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT71), .B1(new_n349), .B2(new_n344), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT71), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n323), .A2(new_n324), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT68), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n323), .A2(new_n309), .A3(new_n324), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n351), .B(new_n343), .C1(new_n355), .C2(G169), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n350), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT73), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT10), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n361), .A2(KEYINPUT10), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n312), .A2(G223), .A3(new_n313), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n316), .A2(G222), .ZN(new_n365));
  OR2_X1    g0165(.A1(KEYINPUT3), .A2(G33), .ZN(new_n366));
  NAND2_X1  g0166(.A1(KEYINPUT3), .A2(G33), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n364), .B(new_n365), .C1(new_n295), .C2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n260), .B1(new_n369), .B2(new_n254), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n257), .A2(G226), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(G190), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n276), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n202), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n283), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(G50), .A3(new_n281), .ZN(new_n376));
  INV_X1    g0176(.A(G150), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n334), .A2(new_n294), .B1(new_n377), .B2(new_n297), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(G20), .B2(new_n203), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n374), .B(new_n376), .C1(new_n379), .C2(new_n284), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT9), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n370), .A2(new_n371), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n372), .B(new_n382), .C1(new_n383), .C2(new_n345), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n381), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT72), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n362), .B(new_n363), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n372), .A2(new_n382), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n345), .B1(new_n370), .B2(new_n371), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT72), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n385), .B(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n390), .A2(new_n392), .A3(new_n361), .A4(KEYINPUT10), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n383), .A2(new_n357), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(new_n380), .C1(G169), .C2(new_n383), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n387), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT18), .ZN(new_n397));
  OAI211_X1 g0197(.A(G226), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n398));
  OAI211_X1 g0198(.A(G223), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n254), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n253), .A2(G232), .A3(new_n256), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n402), .A2(new_n357), .A3(new_n261), .A4(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT79), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n260), .B(new_n403), .C1(new_n401), .C2(new_n254), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n405), .B(new_n406), .C1(new_n407), .C2(G169), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n402), .A2(new_n261), .A3(new_n404), .ZN(new_n410));
  INV_X1    g0210(.A(G169), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n406), .B1(new_n412), .B2(new_n405), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n334), .B1(new_n206), .B2(G20), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(new_n375), .B1(new_n373), .B2(new_n334), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n246), .A2(new_n247), .A3(G20), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT76), .B(KEYINPUT7), .Z(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT78), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(KEYINPUT7), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n366), .A2(new_n207), .A3(new_n367), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT78), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n420), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G68), .ZN(new_n427));
  AND2_X1   g0227(.A1(G58), .A2(G68), .ZN(new_n428));
  OAI21_X1  g0228(.A(G20), .B1(new_n428), .B2(new_n201), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT77), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n296), .A2(G159), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT77), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(G20), .C1(new_n428), .C2(new_n201), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n427), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT16), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n422), .A2(KEYINPUT7), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(G68), .C1(new_n422), .C2(new_n419), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n440), .A3(KEYINPUT16), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n441), .A2(new_n283), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n417), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n397), .B1(new_n414), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT16), .B1(new_n427), .B2(new_n435), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n441), .A2(new_n283), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n416), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(KEYINPUT18), .C1(new_n413), .C2(new_n409), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G190), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n402), .A2(new_n450), .A3(new_n261), .A4(new_n404), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT80), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n410), .A2(new_n345), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n260), .B1(new_n401), .B2(new_n254), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT80), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n454), .A2(new_n455), .A3(new_n450), .A4(new_n404), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT81), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT81), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n452), .A2(new_n453), .A3(new_n459), .A4(new_n456), .ZN(new_n460));
  AOI211_X1 g0260(.A(KEYINPUT17), .B(new_n447), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT17), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n460), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(new_n443), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n449), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NOR4_X1   g0265(.A1(new_n308), .A2(new_n360), .A3(new_n396), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n206), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n276), .A2(new_n467), .A3(new_n222), .A4(new_n282), .ZN(new_n468));
  INV_X1    g0268(.A(G107), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n276), .A2(G107), .ZN(new_n471));
  XOR2_X1   g0271(.A(new_n471), .B(KEYINPUT25), .Z(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n474));
  OAI21_X1  g0274(.A(G20), .B1(new_n318), .B2(new_n319), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(KEYINPUT23), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n207), .B(G87), .C1(new_n246), .C2(new_n247), .ZN(new_n477));
  XNOR2_X1  g0277(.A(KEYINPUT91), .B(KEYINPUT22), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT22), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(KEYINPUT91), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n368), .A2(new_n207), .A3(G87), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n476), .A2(new_n479), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n484), .B(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n470), .B(new_n473), .C1(new_n486), .C2(new_n284), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT93), .ZN(new_n489));
  OAI211_X1 g0289(.A(G257), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n490));
  OAI211_X1 g0290(.A(G250), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G294), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT92), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT92), .A4(new_n492), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n254), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n206), .A2(G45), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT5), .A2(G41), .ZN(new_n500));
  AND2_X1   g0300(.A1(KEYINPUT5), .A2(G41), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n499), .B(G274), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n499), .B1(new_n501), .B2(new_n500), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(G264), .A3(new_n253), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n497), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n489), .B1(new_n505), .B2(new_n345), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n489), .A3(new_n345), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n505), .A2(G190), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n488), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT88), .ZN(new_n512));
  OAI211_X1 g0312(.A(G238), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  INV_X1    g0314(.A(G244), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n514), .C1(new_n310), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n254), .ZN(new_n517));
  INV_X1    g0317(.A(G45), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT86), .B1(new_n518), .B2(G1), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT86), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(new_n206), .A3(G45), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n253), .A2(new_n519), .A3(new_n521), .A4(G250), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT87), .ZN(new_n523));
  INV_X1    g0323(.A(G250), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n498), .B2(KEYINPUT86), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT87), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n525), .A2(new_n526), .A3(new_n253), .A4(new_n521), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n499), .A2(G274), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n517), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n512), .B1(new_n530), .B2(new_n450), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(G200), .ZN(new_n532));
  INV_X1    g0332(.A(G87), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n468), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n337), .B1(new_n277), .B2(new_n279), .ZN(new_n535));
  INV_X1    g0335(.A(G97), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n533), .B(new_n536), .C1(new_n318), .C2(new_n319), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n207), .B1(new_n250), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n368), .A2(new_n207), .A3(G68), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n538), .B1(new_n250), .B2(G20), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n534), .B(new_n535), .C1(new_n543), .C2(new_n283), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n516), .A2(new_n254), .B1(G274), .B2(new_n499), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n545), .A2(KEYINPUT88), .A3(G190), .A4(new_n528), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n531), .A2(new_n532), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n535), .B1(new_n543), .B2(new_n283), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n338), .B2(new_n468), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n530), .A2(new_n411), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n357), .A3(new_n528), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n505), .A2(new_n411), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n497), .A2(new_n504), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(new_n357), .A3(new_n502), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n487), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G264), .ZN(new_n559));
  INV_X1    g0359(.A(G303), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n310), .A2(new_n559), .B1(new_n368), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G257), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n254), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n503), .A2(G270), .A3(new_n253), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n502), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n216), .B1(new_n206), .B2(G33), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n280), .A2(new_n284), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(G33), .ZN(new_n569));
  AOI21_X1  g0369(.A(G20), .B1(new_n569), .B2(G97), .ZN(new_n570));
  NAND3_X1  g0370(.A1(KEYINPUT84), .A2(G33), .A3(G283), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT84), .B1(G33), .B2(G283), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n282), .A2(new_n222), .B1(G20), .B2(new_n216), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT20), .B1(new_n574), .B2(new_n575), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n568), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT89), .B1(new_n341), .B2(new_n216), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT89), .ZN(new_n581));
  AOI211_X1 g0381(.A(new_n581), .B(G116), .C1(new_n277), .C2(new_n279), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n579), .A2(new_n583), .A3(KEYINPUT90), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT90), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n284), .A2(new_n277), .A3(new_n279), .A4(new_n567), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT20), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n207), .B1(new_n536), .B2(G33), .ZN(new_n588));
  INV_X1    g0388(.A(new_n573), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(new_n571), .ZN(new_n590));
  INV_X1    g0390(.A(new_n575), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n586), .B1(new_n592), .B2(new_n576), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n341), .A2(new_n216), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n581), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n341), .A2(KEYINPUT89), .A3(new_n216), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n585), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G169), .B(new_n566), .C1(new_n584), .C2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT90), .B1(new_n579), .B2(new_n583), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n593), .A2(new_n597), .A3(new_n585), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n564), .A2(new_n502), .A3(new_n565), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(G179), .A3(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(KEYINPUT21), .A3(G169), .A4(new_n566), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(G190), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n566), .A2(G200), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n603), .A4(new_n602), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n601), .A2(new_n606), .A3(new_n607), .A4(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n245), .B1(new_n366), .B2(new_n367), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(G250), .B1(new_n589), .B2(new_n571), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  OAI211_X1 g0414(.A(G244), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(KEYINPUT82), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT4), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n615), .B2(new_n614), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n613), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n616), .A2(KEYINPUT4), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n254), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n503), .A2(G257), .A3(new_n253), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n502), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT85), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT85), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n625), .A3(new_n502), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n411), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n373), .A2(new_n536), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n468), .B2(new_n536), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT6), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n240), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n469), .A2(KEYINPUT6), .A3(G97), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n207), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n297), .A2(new_n295), .ZN(new_n637));
  AOI211_X1 g0437(.A(new_n636), .B(new_n637), .C1(new_n426), .C2(new_n320), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n632), .B1(new_n638), .B2(new_n284), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n621), .A2(new_n627), .A3(new_n357), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n629), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n628), .A2(G200), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n426), .A2(new_n320), .ZN(new_n643));
  INV_X1    g0443(.A(new_n636), .ZN(new_n644));
  INV_X1    g0444(.A(new_n637), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n631), .B1(new_n646), .B2(new_n283), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n621), .A2(new_n627), .A3(G190), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n642), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n611), .A2(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n466), .A2(new_n511), .A3(new_n558), .A4(new_n651), .ZN(G372));
  NAND2_X1  g0452(.A1(new_n547), .A2(new_n552), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT26), .B1(new_n641), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n545), .A2(G190), .A3(new_n528), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n532), .A2(new_n544), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n552), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n646), .A2(new_n283), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n616), .A2(KEYINPUT4), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n659), .B(new_n613), .C1(new_n616), .C2(new_n618), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n254), .B1(new_n624), .B2(new_n626), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n658), .A2(new_n632), .B1(new_n661), .B2(new_n357), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n657), .A2(new_n662), .A3(new_n663), .A4(new_n629), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n654), .A2(new_n664), .A3(new_n552), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n641), .A2(new_n649), .A3(new_n657), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n557), .A2(new_n601), .A3(new_n606), .A4(new_n607), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n511), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n466), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT94), .Z(new_n671));
  AOI21_X1  g0471(.A(new_n447), .B1(new_n458), .B2(new_n460), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(new_n462), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n307), .A2(new_n350), .A3(new_n358), .A4(new_n356), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n302), .B1(new_n272), .B2(new_n274), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT95), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(new_n449), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n461), .A2(new_n464), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n304), .B2(new_n674), .ZN(new_n681));
  INV_X1    g0481(.A(new_n449), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT95), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n387), .A2(new_n393), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n679), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(new_n395), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n671), .A2(new_n686), .ZN(G369));
  NAND3_X1  g0487(.A1(new_n601), .A2(new_n606), .A3(new_n607), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n291), .A2(G20), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n206), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n602), .B2(new_n603), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n688), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n611), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n557), .A2(new_n695), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n511), .B1(new_n488), .B2(new_n696), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(new_n557), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n688), .A2(new_n696), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n702), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n208), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n537), .A2(G116), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n224), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n669), .A2(new_n696), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n553), .A2(new_n663), .A3(new_n629), .A4(new_n662), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n552), .A2(new_n656), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT26), .B1(new_n641), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n668), .A2(new_n552), .A3(new_n720), .A4(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .A3(new_n696), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n695), .B1(new_n665), .B2(new_n668), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT96), .B1(new_n725), .B2(KEYINPUT29), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n719), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n651), .A2(new_n511), .A3(new_n558), .A4(new_n696), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n555), .A2(new_n621), .A3(new_n627), .ZN(new_n730));
  INV_X1    g0530(.A(new_n530), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n605), .A2(new_n731), .A3(G179), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n566), .A2(new_n530), .A3(new_n357), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(new_n661), .A3(KEYINPUT30), .A4(new_n555), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n731), .A2(G179), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n628), .A3(new_n505), .A4(new_n566), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n733), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n695), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n728), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n727), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n715), .B1(new_n745), .B2(G1), .ZN(G364));
  NOR3_X1   g0546(.A1(new_n207), .A2(new_n357), .A3(new_n345), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n450), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G326), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n315), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n207), .A2(new_n450), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n345), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n357), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G322), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n560), .A2(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n207), .A2(G190), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n759), .B1(G329), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G283), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n760), .A2(new_n754), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n207), .B1(new_n761), .B2(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n752), .B(new_n767), .C1(G294), .C2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n756), .A2(new_n760), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT99), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(new_n748), .B2(G190), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n747), .A2(KEYINPUT99), .A3(new_n450), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT33), .B(G317), .Z(new_n778));
  OAI221_X1 g0578(.A(new_n770), .B1(new_n771), .B2(new_n772), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G58), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n750), .A2(new_n202), .B1(new_n780), .B2(new_n757), .ZN(new_n781));
  INV_X1    g0581(.A(new_n772), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(G77), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n776), .A2(G68), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n768), .A2(new_n536), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G159), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n762), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT32), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n783), .A2(new_n784), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n755), .A2(new_n533), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n766), .A2(new_n469), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n791), .A2(new_n792), .A3(new_n315), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT98), .Z(new_n794));
  OAI21_X1  g0594(.A(new_n779), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n222), .B1(G20), .B2(new_n411), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n291), .A2(new_n569), .A3(KEYINPUT97), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT97), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G13), .B2(G33), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n796), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n239), .A2(G45), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n709), .A2(new_n368), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n804), .B(new_n805), .C1(G45), .C2(new_n224), .ZN(new_n806));
  INV_X1    g0606(.A(G355), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n368), .A2(new_n208), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(G116), .B2(new_n208), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n795), .A2(new_n796), .B1(new_n803), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n802), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n699), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n206), .B1(new_n689), .B2(G45), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n710), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n700), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n699), .A2(G330), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n812), .A2(new_n816), .B1(new_n817), .B2(new_n818), .ZN(G396));
  AOI22_X1  g0619(.A1(new_n749), .A2(G137), .B1(G159), .B2(new_n782), .ZN(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n821), .B2(new_n757), .C1(new_n777), .C2(new_n377), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT34), .ZN(new_n823));
  INV_X1    g0623(.A(new_n766), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G68), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n315), .B1(new_n763), .B2(G132), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n202), .B2(new_n755), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G58), .B2(new_n769), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n823), .A2(new_n825), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n766), .A2(new_n533), .ZN(new_n830));
  INV_X1    g0630(.A(G294), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n757), .A2(new_n831), .B1(new_n762), .B2(new_n771), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G116), .B2(new_n782), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n315), .B1(new_n755), .B2(new_n469), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n785), .B(new_n834), .C1(G303), .C2(new_n749), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n776), .A2(KEYINPUT100), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n776), .A2(KEYINPUT100), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n833), .B(new_n835), .C1(new_n838), .C2(new_n765), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n829), .B1(new_n830), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n800), .A2(new_n796), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n840), .A2(new_n796), .B1(new_n295), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n344), .A2(new_n696), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n348), .B2(new_n359), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n359), .A2(new_n843), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n815), .B(new_n842), .C1(new_n846), .C2(new_n801), .ZN(new_n847));
  INV_X1    g0647(.A(new_n846), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT101), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT101), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n851), .A3(new_n716), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n359), .A2(new_n843), .ZN(new_n853));
  INV_X1    g0653(.A(new_n843), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n350), .A2(new_n356), .A3(new_n358), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n343), .B(new_n346), .C1(new_n330), .C2(new_n331), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n725), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(new_n744), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n847), .B1(new_n860), .B2(new_n815), .ZN(G384));
  INV_X1    g0661(.A(new_n693), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n435), .A2(new_n440), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n437), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n417), .B1(new_n442), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n465), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n412), .A2(new_n405), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT79), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n434), .B1(new_n426), .B2(G68), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n283), .B(new_n441), .C1(new_n870), .C2(KEYINPUT16), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n869), .A2(new_n408), .B1(new_n871), .B2(new_n416), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n672), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n693), .B1(new_n871), .B2(new_n416), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n865), .B1(new_n414), .B2(new_n693), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n878), .B2(new_n672), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n867), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n304), .A2(new_n696), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT103), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n275), .B2(new_n303), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n302), .A2(new_n696), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n888), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NOR4_X1   g0693(.A1(new_n676), .A2(new_n889), .A3(KEYINPUT103), .A4(new_n891), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n887), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n508), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n896), .A2(new_n506), .A3(new_n510), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n553), .B(new_n557), .C1(new_n897), .C2(new_n487), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n898), .A2(new_n611), .A3(new_n650), .A4(new_n695), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n741), .A2(new_n742), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n857), .B(new_n853), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n885), .A2(new_n895), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n304), .A2(new_n307), .A3(new_n892), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT103), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n890), .A2(new_n888), .A3(new_n892), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n886), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n901), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n876), .B1(new_n673), .B2(new_n449), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n874), .B1(new_n873), .B2(new_n876), .ZN(new_n911));
  NOR4_X1   g0711(.A1(new_n672), .A2(new_n872), .A3(KEYINPUT37), .A4(new_n875), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n882), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n904), .B1(new_n914), .B2(new_n884), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n903), .A2(new_n904), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n466), .A2(new_n743), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(G330), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n449), .A2(new_n862), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n359), .A2(new_n695), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n858), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n895), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT38), .B1(new_n867), .B2(new_n880), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n921), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n304), .A2(new_n695), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT39), .B1(new_n926), .B2(new_n927), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n914), .A2(new_n933), .A3(new_n884), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n719), .A2(new_n466), .A3(new_n726), .A4(new_n724), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n686), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n919), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n206), .B2(new_n689), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n634), .A2(new_n635), .ZN(new_n942));
  OAI211_X1 g0742(.A(G116), .B(new_n223), .C1(new_n942), .C2(KEYINPUT35), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT102), .Z(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(KEYINPUT35), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  OAI21_X1  g0747(.A(G77), .B1(new_n780), .B2(new_n286), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n948), .A2(new_n224), .B1(G50), .B2(new_n286), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n291), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n941), .A2(new_n947), .A3(new_n950), .ZN(G367));
  NOR2_X1   g0751(.A1(new_n755), .A2(new_n216), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT46), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n315), .B1(new_n750), .B2(new_n771), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n766), .A2(new_n536), .ZN(new_n955));
  INV_X1    g0755(.A(G317), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n757), .A2(new_n560), .B1(new_n762), .B2(new_n956), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n953), .B(new_n958), .C1(new_n320), .C2(new_n769), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n959), .B1(new_n765), .B2(new_n772), .C1(new_n831), .C2(new_n838), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n766), .A2(new_n295), .ZN(new_n961));
  INV_X1    g0761(.A(new_n757), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(G150), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n202), .B2(new_n772), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n750), .A2(new_n821), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n368), .B1(new_n755), .B2(new_n780), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n768), .A2(new_n286), .ZN(new_n967));
  NOR4_X1   g0767(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(G137), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n968), .B1(new_n969), .B2(new_n762), .C1(new_n838), .C2(new_n787), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n960), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n816), .B1(new_n972), .B2(new_n796), .ZN(new_n973));
  INV_X1    g0773(.A(new_n805), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n803), .B1(new_n208), .B2(new_n338), .C1(new_n235), .C2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n544), .A2(new_n696), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n552), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n657), .B2(new_n976), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT104), .Z(new_n979));
  OAI211_X1 g0779(.A(new_n973), .B(new_n975), .C1(new_n811), .C2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n813), .B(KEYINPUT106), .Z(new_n981));
  XNOR2_X1  g0781(.A(new_n704), .B(new_n706), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n701), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n745), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT105), .Z(new_n985));
  OAI211_X1 g0785(.A(new_n641), .B(new_n649), .C1(new_n647), .C2(new_n696), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n641), .B2(new_n696), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n707), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT45), .Z(new_n989));
  NOR2_X1   g0789(.A1(new_n707), .A2(new_n987), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT44), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n705), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n705), .A3(new_n991), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n745), .B1(new_n985), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n710), .B(KEYINPUT41), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n981), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n704), .A2(new_n706), .A3(new_n987), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT42), .Z(new_n1001));
  OAI21_X1  g0801(.A(new_n641), .B1(new_n986), .B2(new_n557), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n696), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1001), .A2(new_n1003), .B1(KEYINPUT43), .B2(new_n979), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n993), .A2(new_n987), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1004), .B(new_n1005), .Z(new_n1006));
  NOR2_X1   g0806(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n980), .B1(new_n999), .B2(new_n1008), .ZN(G387));
  OR2_X1    g0809(.A1(new_n983), .A2(new_n745), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(new_n710), .A3(new_n984), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n983), .A2(new_n981), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n749), .A2(G322), .B1(G303), .B2(new_n782), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n956), .B2(new_n757), .C1(new_n838), .C2(new_n771), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT48), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n755), .A2(new_n831), .B1(new_n768), .B2(new_n765), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT110), .Z(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT49), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n368), .B1(new_n824), .B2(G116), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n751), .C2(new_n762), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n755), .A2(new_n295), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n757), .A2(new_n202), .B1(new_n772), .B2(new_n286), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G150), .C2(new_n763), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n315), .B(new_n955), .C1(new_n749), .C2(G159), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n776), .A2(new_n335), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n338), .A2(new_n768), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1021), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n796), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n712), .B(KEYINPUT107), .ZN(new_n1032));
  XOR2_X1   g0832(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n1033));
  AND3_X1   g0833(.A1(new_n335), .A2(new_n202), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1033), .B1(new_n335), .B2(new_n202), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1034), .A2(new_n1035), .A3(G45), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1032), .B(new_n1036), .C1(new_n286), .C2(new_n295), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n805), .B(new_n1037), .C1(new_n232), .C2(new_n518), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(G107), .B2(new_n208), .C1(new_n712), .C2(new_n808), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n816), .B1(new_n1039), .B2(new_n803), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT109), .Z(new_n1041));
  OAI211_X1 g0841(.A(new_n1031), .B(new_n1041), .C1(new_n704), .C2(new_n811), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1011), .A2(new_n1012), .A3(new_n1042), .ZN(G393));
  NOR2_X1   g0843(.A1(new_n985), .A2(new_n996), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n711), .B(new_n1044), .C1(new_n996), .C2(new_n984), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n749), .A2(G317), .B1(G311), .B2(new_n962), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT52), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n368), .B(new_n1047), .C1(G116), .C2(new_n769), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n755), .A2(new_n765), .B1(new_n772), .B2(new_n831), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n792), .B(new_n1049), .C1(G322), .C2(new_n763), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1048), .B(new_n1050), .C1(new_n560), .C2(new_n838), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n838), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(G50), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n749), .A2(G150), .B1(G159), .B2(new_n962), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT51), .Z(new_n1055));
  NOR2_X1   g0855(.A1(new_n768), .A2(new_n295), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n755), .A2(new_n286), .B1(new_n762), .B2(new_n821), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n335), .C2(new_n782), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1053), .A2(new_n368), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1051), .B1(new_n830), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n816), .B1(new_n1060), .B2(new_n796), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n803), .B1(new_n536), .B2(new_n208), .C1(new_n242), .C2(new_n974), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n811), .C2(new_n987), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n996), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT111), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n981), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1045), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(G390));
  AOI21_X1  g0869(.A(new_n930), .B1(new_n914), .B2(new_n884), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n720), .A2(new_n722), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n897), .A2(new_n487), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n641), .A2(new_n649), .A3(new_n657), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1071), .B1(new_n1074), .B2(new_n667), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n695), .B1(new_n1075), .B2(new_n552), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n922), .B1(new_n1076), .B2(new_n846), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1070), .B1(new_n1077), .B2(new_n908), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n932), .A2(new_n934), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n930), .B1(new_n924), .B2(new_n895), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n743), .A2(new_n846), .A3(G330), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT112), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n908), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1078), .B(new_n1084), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n981), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT54), .B(G143), .Z(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n838), .A2(new_n969), .B1(new_n772), .B2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT114), .ZN(new_n1093));
  INV_X1    g0893(.A(G125), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n368), .B1(new_n762), .B2(new_n1094), .C1(new_n202), .C2(new_n766), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT53), .B1(new_n755), .B2(new_n377), .ZN(new_n1096));
  OR3_X1    g0896(.A1(new_n755), .A2(KEYINPUT53), .A3(new_n377), .ZN(new_n1097));
  INV_X1    g0897(.A(G128), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1096), .B(new_n1097), .C1(new_n750), .C2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1095), .B(new_n1099), .C1(G132), .C2(new_n962), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1093), .B(new_n1100), .C1(new_n787), .C2(new_n768), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT115), .Z(new_n1102));
  OAI221_X1 g0902(.A(new_n825), .B1(new_n536), .B2(new_n772), .C1(new_n831), .C2(new_n762), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1056), .B(new_n1103), .C1(G116), .C2(new_n962), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n368), .B(new_n791), .C1(new_n749), .C2(G283), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n320), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1104), .B(new_n1105), .C1(new_n1106), .C2(new_n838), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n816), .B1(new_n1108), .B2(new_n796), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n841), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1109), .B1(new_n335), .B2(new_n1110), .C1(new_n1079), .C2(new_n801), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n466), .A2(G330), .A3(new_n743), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n937), .A2(new_n395), .A3(new_n685), .A4(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n902), .A2(new_n895), .A3(G330), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n744), .B1(new_n849), .B2(new_n851), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n1077), .C1(new_n1116), .C2(new_n895), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n908), .A2(new_n1082), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n924), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1114), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(new_n1088), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT113), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1113), .B(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1121), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1087), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n922), .B1(new_n846), .B2(new_n725), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n931), .B1(new_n908), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(new_n932), .A3(new_n934), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1084), .B1(new_n1131), .B2(new_n1078), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n710), .B1(new_n1127), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1089), .B(new_n1111), .C1(new_n1124), .C2(new_n1134), .ZN(G378));
  INV_X1    g0935(.A(KEYINPUT57), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n902), .A2(new_n895), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n904), .B1(new_n1137), .B2(new_n928), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n909), .A2(new_n915), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1138), .A2(new_n1139), .A3(G330), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT56), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n380), .A2(new_n862), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n396), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT55), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n387), .A2(new_n393), .A3(new_n395), .A4(new_n1142), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1141), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(KEYINPUT55), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(KEYINPUT56), .A3(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1149), .A2(new_n1153), .A3(KEYINPUT117), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n929), .B2(new_n935), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n933), .B1(new_n883), .B2(new_n884), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n914), .A2(new_n933), .A3(new_n884), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n930), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n906), .A2(new_n907), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1159), .A2(new_n887), .B1(new_n858), .B2(new_n923), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n920), .B1(new_n1160), .B2(new_n885), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1149), .A2(new_n1153), .A3(KEYINPUT117), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1158), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1140), .A2(new_n1155), .A3(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1155), .A2(new_n1163), .B1(G330), .B2(new_n916), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1114), .B1(new_n1088), .B2(new_n1121), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1136), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1126), .B1(new_n1133), .B2(new_n1122), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n916), .A2(G330), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n929), .A2(new_n1154), .A3(new_n935), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1162), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1140), .A2(new_n1155), .A3(new_n1163), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1169), .A2(new_n1175), .A3(KEYINPUT57), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1168), .A2(new_n710), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1149), .A2(new_n1153), .A3(new_n800), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n841), .A2(new_n202), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1091), .A2(new_n755), .B1(new_n772), .B2(new_n969), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n750), .A2(new_n1094), .B1(new_n377), .B2(new_n768), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G132), .C2(new_n776), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1098), .B2(new_n757), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT59), .Z(new_n1184));
  AOI21_X1  g0984(.A(G41), .B1(new_n824), .B2(G159), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT116), .ZN(new_n1186));
  INV_X1    g0986(.A(G124), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n762), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1184), .A2(new_n569), .A3(new_n1185), .A4(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n202), .B1(new_n246), .B2(G41), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n750), .A2(new_n216), .ZN(new_n1192));
  OR4_X1    g0992(.A1(G41), .A2(new_n1192), .A3(new_n368), .A4(new_n1022), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n777), .A2(new_n536), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n962), .A2(G107), .B1(new_n782), .B2(new_n337), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n780), .B2(new_n766), .C1(new_n765), .C2(new_n762), .ZN(new_n1196));
  NOR4_X1   g0996(.A1(new_n1193), .A2(new_n967), .A3(new_n1194), .A4(new_n1196), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT58), .Z(new_n1198));
  NAND3_X1  g0998(.A1(new_n1190), .A2(new_n1191), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n816), .B1(new_n1199), .B2(new_n796), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1178), .A2(new_n1179), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1166), .B2(new_n1066), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1177), .A2(new_n1203), .ZN(G375));
  NAND2_X1  g1004(.A1(new_n1114), .A2(new_n1122), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(new_n1127), .A3(new_n998), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1052), .A2(G116), .B1(new_n320), .B2(new_n782), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT118), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n536), .A2(new_n755), .B1(new_n757), .B2(new_n765), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1210), .B(new_n1027), .C1(G303), .C2(new_n763), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n368), .B(new_n961), .C1(new_n749), .C2(G294), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n766), .A2(new_n780), .B1(new_n768), .B2(new_n202), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n315), .B(new_n1215), .C1(G132), .C2(new_n749), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n772), .A2(new_n377), .B1(new_n762), .B2(new_n1098), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G137), .B2(new_n962), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n787), .B2(new_n755), .C1(new_n838), .C2(new_n1091), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1214), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n796), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(G68), .B2(new_n1110), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n816), .B(new_n1223), .C1(new_n908), .C2(new_n800), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1121), .B2(new_n981), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1206), .A2(new_n1225), .ZN(G381));
  XOR2_X1   g1026(.A(G375), .B(KEYINPUT119), .Z(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(G378), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(G390), .A2(G387), .A3(G396), .A4(G393), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(G381), .A2(G384), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(G407));
  INV_X1    g1031(.A(G213), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1228), .B2(new_n694), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(G407), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT120), .ZN(G409));
  NAND3_X1  g1035(.A1(new_n1177), .A2(G378), .A3(new_n1203), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1089), .A2(new_n1111), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n711), .B1(new_n1123), .B2(new_n1088), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1127), .A2(new_n1133), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1169), .A2(new_n1175), .A3(new_n998), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1240), .B1(new_n1241), .B2(new_n1202), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1236), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT60), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1126), .B2(new_n1121), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1114), .A2(new_n1122), .A3(KEYINPUT60), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1245), .A2(new_n1246), .A3(new_n710), .A4(new_n1127), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1225), .ZN(new_n1248));
  INV_X1    g1048(.A(G384), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1247), .A2(G384), .A3(new_n1225), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1232), .A2(G343), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1243), .A2(KEYINPUT62), .A3(new_n1253), .A4(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT125), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1254), .B1(new_n1236), .B2(new_n1242), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1259), .A2(KEYINPUT125), .A3(KEYINPUT62), .A4(new_n1253), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT124), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1253), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1262), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  AOI211_X1 g1065(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n1259), .C2(new_n1253), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1261), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT123), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1254), .A2(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1255), .A2(KEYINPUT121), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1253), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1250), .A2(new_n1251), .A3(new_n1272), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1269), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1259), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1268), .B1(new_n1276), .B2(KEYINPUT61), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1274), .B(new_n1270), .ZN(new_n1279));
  OAI211_X1 g1079(.A(KEYINPUT123), .B(new_n1278), .C1(new_n1279), .C2(new_n1259), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(KEYINPUT126), .B1(new_n1267), .B2(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1068), .A2(G387), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1068), .A2(G387), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  XOR2_X1   g1085(.A(G393), .B(G396), .Z(new_n1286));
  AND2_X1   g1086(.A1(new_n1068), .A2(G387), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1285), .A2(new_n1286), .B1(KEYINPUT122), .B2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1286), .A2(KEYINPUT122), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1283), .A2(new_n1284), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1243), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT124), .B1(new_n1293), .B2(KEYINPUT62), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1263), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1294), .A2(new_n1258), .A3(new_n1260), .A4(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1277), .A4(new_n1280), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1282), .A2(new_n1292), .A3(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1263), .B1(new_n1276), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1293), .A2(KEYINPUT63), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1291), .A2(new_n1278), .A3(new_n1301), .A4(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1299), .A2(new_n1303), .ZN(G405));
  NAND2_X1  g1104(.A1(G375), .A2(new_n1240), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1236), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1253), .A2(KEYINPUT127), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT127), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1252), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1307), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1310), .B2(new_n1307), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1291), .B(new_n1312), .ZN(G402));
endmodule


