//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  INV_X1    g0000(.A(KEYINPUT65), .ZN(new_n201));
  XNOR2_X1  g0001(.A(KEYINPUT64), .B(G50), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(G58), .A2(G68), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g0005(.A(new_n201), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  NAND3_X1  g0007(.A1(new_n202), .A2(KEYINPUT65), .A3(new_n204), .ZN(new_n208));
  AND3_X1   g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n205), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT66), .B(G238), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n221), .A2(G68), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G107), .A2(G264), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n217), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n218), .B1(new_n206), .B2(new_n208), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  OR2_X1    g0050(.A1(new_n250), .A2(KEYINPUT8), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(KEYINPUT8), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n218), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n218), .A2(new_n256), .A3(KEYINPUT68), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G20), .B2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n254), .A2(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n248), .B1(new_n249), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT69), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n265), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n268), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n248), .ZN(new_n274));
  INV_X1    g0074(.A(G50), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n268), .B2(G20), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n274), .A2(new_n276), .B1(new_n275), .B2(new_n273), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n266), .A2(new_n267), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G169), .ZN(new_n279));
  AND2_X1   g0079(.A1(G1), .A2(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT67), .B1(new_n290), .B2(G1698), .ZN(new_n291));
  OAI21_X1  g0091(.A(G223), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n286), .A2(G1698), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n293), .A2(G222), .B1(G77), .B2(new_n286), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n282), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n280), .B2(new_n281), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n282), .A2(new_n298), .ZN(new_n301));
  INV_X1    g0101(.A(G226), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n279), .B1(new_n295), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n278), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n295), .A2(new_n303), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n305), .A2(KEYINPUT71), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(KEYINPUT71), .B2(new_n305), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(new_n267), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n277), .B1(new_n264), .B2(new_n265), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT9), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT9), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n266), .A2(new_n314), .A3(new_n267), .A4(new_n277), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(G190), .B2(new_n307), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n310), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n316), .A2(new_n310), .A3(new_n319), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n309), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT17), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT7), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n290), .A2(new_n324), .A3(G20), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT7), .B1(new_n286), .B2(new_n218), .ZN(new_n326));
  OAI21_X1  g0126(.A(G68), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n260), .A2(G159), .ZN(new_n328));
  INV_X1    g0128(.A(G68), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n250), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(G20), .B1(new_n330), .B2(new_n204), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n327), .A2(new_n333), .A3(KEYINPUT16), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n324), .B1(new_n290), .B2(G20), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n329), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n338), .B2(new_n332), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n339), .A3(new_n248), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n268), .A2(G20), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n253), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n274), .A2(new_n342), .B1(new_n254), .B2(new_n273), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n300), .B1(new_n301), .B2(new_n232), .ZN(new_n344));
  OR2_X1    g0144(.A1(G223), .A2(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n302), .A2(G1698), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n283), .A2(new_n345), .A3(new_n285), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G87), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n282), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(KEYINPUT74), .A3(new_n348), .ZN(new_n352));
  AOI211_X1 g0152(.A(G190), .B(new_n344), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(new_n350), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(new_n352), .ZN(new_n356));
  INV_X1    g0156(.A(new_n344), .ZN(new_n357));
  AOI21_X1  g0157(.A(G200), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n340), .B(new_n343), .C1(new_n353), .C2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT76), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n356), .A2(new_n362), .A3(new_n357), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n344), .B1(new_n351), .B2(new_n352), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(G200), .B2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n365), .A2(KEYINPUT76), .A3(new_n340), .A4(new_n343), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n323), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT18), .ZN(new_n368));
  INV_X1    g0168(.A(new_n348), .ZN(new_n369));
  NOR2_X1   g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n302), .B2(G1698), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n369), .B1(new_n371), .B2(new_n290), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n355), .B1(new_n372), .B2(KEYINPUT74), .ZN(new_n373));
  INV_X1    g0173(.A(new_n352), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n357), .B(G179), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n364), .B2(new_n279), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n376), .A2(new_n377), .B1(new_n340), .B2(new_n343), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n375), .B(KEYINPUT75), .C1(new_n279), .C2(new_n364), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n368), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI211_X1 g0180(.A(new_n306), .B(new_n344), .C1(new_n351), .C2(new_n352), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n279), .B1(new_n356), .B2(new_n357), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n377), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n340), .A2(new_n343), .ZN(new_n384));
  AND4_X1   g0184(.A1(new_n368), .A2(new_n383), .A3(new_n384), .A4(new_n379), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n359), .A2(new_n323), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NOR4_X1   g0187(.A1(new_n367), .A2(new_n380), .A3(new_n385), .A4(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n286), .A2(new_n232), .A3(G1698), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(G107), .B2(new_n286), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n221), .B1(new_n289), .B2(new_n291), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n282), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G244), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n300), .B1(new_n301), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n279), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G20), .A2(G77), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT15), .B(G87), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n397), .B1(new_n255), .B2(new_n398), .C1(new_n254), .C2(new_n261), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n207), .B1(new_n268), .B2(G20), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n399), .A2(new_n248), .B1(new_n274), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n273), .A2(new_n207), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT72), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n396), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n395), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n391), .A2(new_n392), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n306), .B(new_n406), .C1(new_n407), .C2(new_n282), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(G190), .B(new_n406), .C1(new_n407), .C2(new_n282), .ZN(new_n410));
  OAI21_X1  g0210(.A(G200), .B1(new_n393), .B2(new_n395), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n410), .A2(new_n403), .A3(new_n411), .A4(new_n401), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT73), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n273), .A2(new_n329), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT12), .ZN(new_n417));
  INV_X1    g0217(.A(new_n248), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n255), .A2(new_n207), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(G20), .B2(new_n329), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n260), .A2(G50), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n422), .A2(KEYINPUT11), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n274), .A2(G68), .A3(new_n341), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(KEYINPUT11), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n417), .A2(new_n423), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT14), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n290), .A2(G232), .A3(G1698), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n290), .A2(G226), .A3(new_n288), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G97), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n355), .ZN(new_n432));
  INV_X1    g0232(.A(new_n301), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n433), .A2(G238), .B1(new_n297), .B2(new_n299), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n432), .B2(new_n434), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n427), .B(G169), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n432), .A2(new_n434), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT13), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(G179), .A3(new_n436), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n436), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n427), .B1(new_n444), .B2(G169), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n426), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(G200), .ZN(new_n447));
  INV_X1    g0247(.A(new_n426), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n447), .B(new_n448), .C1(new_n362), .C2(new_n444), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n409), .A2(KEYINPUT73), .A3(new_n412), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n415), .A2(new_n446), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n322), .A2(new_n389), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n283), .A2(new_n285), .A3(new_n218), .A4(G68), .ZN(new_n453));
  INV_X1    g0253(.A(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT79), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G97), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n255), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n453), .B1(new_n458), .B2(KEYINPUT19), .ZN(new_n459));
  NOR2_X1   g0259(.A1(G87), .A2(G107), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n455), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT19), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n218), .B1(new_n430), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n248), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n273), .A2(new_n398), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n271), .A2(new_n272), .ZN(new_n467));
  INV_X1    g0267(.A(new_n398), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n256), .A2(G1), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n467), .A2(new_n418), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n465), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  INV_X1    g0274(.A(G250), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n268), .B2(G45), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n297), .A2(new_n474), .B1(new_n282), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G238), .A2(G1698), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n394), .B2(G1698), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n481), .B2(new_n290), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n477), .B1(new_n482), .B2(new_n282), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n279), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n477), .B(new_n306), .C1(new_n482), .C2(new_n282), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n394), .A2(G1698), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(G238), .B2(G1698), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n478), .B1(new_n488), .B2(new_n286), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n355), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n490), .A2(new_n491), .A3(new_n306), .A4(new_n477), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n472), .A2(new_n484), .A3(new_n486), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n461), .A2(new_n463), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(new_n453), .C1(KEYINPUT19), .C2(new_n458), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(new_n248), .B1(new_n273), .B2(new_n398), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n483), .A2(G200), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n469), .B(new_n248), .C1(new_n271), .C2(new_n272), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G87), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n490), .A2(G190), .A3(new_n477), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n496), .A2(new_n497), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n493), .A2(KEYINPUT82), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT82), .B1(new_n493), .B2(new_n501), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n498), .A2(G97), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n273), .A2(new_n454), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  INV_X1    g0309(.A(G107), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n454), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n508), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n455), .A2(new_n457), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n510), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n514), .B2(new_n508), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G20), .ZN(new_n516));
  OAI21_X1  g0316(.A(G107), .B1(new_n325), .B2(new_n326), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT77), .B1(new_n260), .B2(G77), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT77), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n519), .B(new_n207), .C1(new_n257), .C2(new_n259), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n516), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n507), .B1(new_n522), .B2(new_n248), .ZN(new_n523));
  XNOR2_X1  g0323(.A(KEYINPUT5), .B(G41), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n297), .A2(new_n474), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(KEYINPUT5), .A2(G41), .ZN(new_n526));
  NOR2_X1   g0326(.A1(KEYINPUT5), .A2(G41), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n474), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n282), .ZN(new_n529));
  INV_X1    g0329(.A(G257), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n283), .A2(new_n285), .A3(G244), .A4(new_n288), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n290), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G283), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n290), .A2(G250), .A3(G1698), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n531), .B1(new_n538), .B2(new_n355), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G169), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n355), .ZN(new_n541));
  INV_X1    g0341(.A(new_n531), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n541), .A2(new_n542), .A3(new_n306), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n523), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n542), .A3(new_n362), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(G200), .B2(new_n539), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n523), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT80), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(KEYINPUT80), .A3(new_n523), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n467), .A2(G116), .A3(new_n418), .A4(new_n470), .ZN(new_n552));
  INV_X1    g0352(.A(G116), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n273), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g0354(.A(KEYINPUT79), .B(G97), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n218), .B(new_n536), .C1(new_n555), .C2(G33), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n247), .A2(new_n217), .B1(G20), .B2(new_n553), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT20), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(G33), .B1(new_n455), .B2(new_n457), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n536), .A2(new_n218), .ZN(new_n560));
  OAI211_X1 g0360(.A(KEYINPUT20), .B(new_n557), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n552), .B(new_n554), .C1(new_n558), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G169), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n528), .A2(G270), .A3(new_n282), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n525), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n286), .A2(G303), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n283), .A2(new_n285), .A3(G264), .A4(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n283), .A2(new_n285), .A3(G257), .A4(new_n288), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT83), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT83), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n567), .A2(new_n572), .A3(new_n568), .A4(new_n569), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n566), .B1(new_n574), .B2(new_n355), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT86), .B1(new_n564), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n554), .A2(new_n552), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT20), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n560), .B1(new_n513), .B2(new_n256), .ZN(new_n579));
  INV_X1    g0379(.A(new_n557), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n561), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n279), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT86), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n282), .B1(new_n571), .B2(new_n573), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n584), .C1(new_n566), .C2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n576), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT84), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n587), .A2(new_n279), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n563), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n589), .B1(new_n591), .B2(new_n575), .ZN(new_n592));
  INV_X1    g0392(.A(new_n590), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n577), .B2(new_n582), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n594), .B(KEYINPUT84), .C1(new_n566), .C2(new_n585), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n574), .A2(new_n355), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n565), .A2(new_n525), .A3(G179), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n563), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT85), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n597), .A2(new_n563), .A3(KEYINPUT85), .A4(new_n599), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n575), .A2(G190), .ZN(new_n605));
  INV_X1    g0405(.A(new_n563), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n605), .B(new_n606), .C1(new_n317), .C2(new_n575), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n588), .A2(new_n596), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n283), .A2(new_n285), .A3(G257), .A4(G1698), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n283), .A2(new_n285), .A3(G250), .A4(new_n288), .ZN(new_n610));
  INV_X1    g0410(.A(G294), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n609), .B(new_n610), .C1(new_n256), .C2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n612), .A2(new_n355), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n528), .A2(G264), .A3(new_n282), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n525), .ZN(new_n615));
  OAI21_X1  g0415(.A(G169), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT88), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n528), .A2(KEYINPUT88), .A3(G264), .A4(new_n282), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n612), .A2(new_n355), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n620), .A2(G179), .A3(new_n525), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n283), .A2(new_n285), .A3(new_n218), .A4(G87), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT22), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT22), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n290), .A2(new_n626), .A3(new_n218), .A4(G87), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(KEYINPUT87), .B(KEYINPUT23), .C1(new_n218), .C2(G107), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT23), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n510), .A3(G20), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n629), .B(new_n631), .C1(G20), .C2(new_n478), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n510), .A2(G20), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT87), .B1(new_n633), .B2(KEYINPUT23), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT24), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT24), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n628), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n418), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n467), .A2(G107), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT25), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n498), .A2(G107), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n623), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n628), .A2(new_n635), .A3(new_n638), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n638), .B1(new_n628), .B2(new_n635), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n248), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n641), .A2(KEYINPUT25), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n641), .A2(KEYINPUT25), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n649), .A2(new_n650), .B1(G107), .B2(new_n498), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n618), .A2(new_n619), .B1(new_n612), .B2(new_n355), .ZN(new_n652));
  AOI21_X1  g0452(.A(G200), .B1(new_n652), .B2(new_n525), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n613), .A2(G190), .A3(new_n615), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n648), .B(new_n651), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n645), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n608), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n452), .A2(new_n504), .A3(new_n551), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n659), .B(KEYINPUT89), .Z(G372));
  NAND2_X1  g0460(.A1(new_n384), .A2(new_n376), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(KEYINPUT18), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n368), .B1(new_n384), .B2(new_n376), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n449), .A2(new_n408), .A3(new_n405), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n446), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n361), .A2(new_n366), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n387), .B1(new_n668), .B2(KEYINPUT17), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n665), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n321), .A2(new_n320), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n309), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(KEYINPUT91), .B(new_n309), .C1(new_n670), .C2(new_n671), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT90), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n504), .B2(new_n544), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n472), .A2(new_n484), .A3(new_n485), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n501), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n544), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n679), .B1(new_n682), .B2(KEYINPUT26), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n676), .B1(new_n678), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n588), .A2(new_n596), .A3(new_n604), .A4(new_n645), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n681), .A2(new_n655), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n551), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n493), .A2(new_n501), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT82), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n493), .A2(new_n501), .A3(KEYINPUT82), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(new_n544), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT26), .ZN(new_n693));
  INV_X1    g0493(.A(new_n679), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n541), .A2(new_n542), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n279), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n539), .A2(new_n306), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n258), .A2(G20), .A3(G33), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT68), .B1(new_n218), .B2(new_n256), .ZN(new_n699));
  OAI21_X1  g0499(.A(G77), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n519), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n260), .A2(KEYINPUT77), .A3(G77), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n510), .B1(new_n336), .B2(new_n337), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n418), .B1(new_n705), .B2(new_n516), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n696), .B(new_n697), .C1(new_n706), .C2(new_n507), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n680), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n694), .B1(new_n708), .B2(new_n677), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n693), .A2(new_n709), .A3(KEYINPUT90), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n684), .A2(new_n687), .A3(new_n710), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n674), .A2(new_n675), .B1(new_n452), .B2(new_n711), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT92), .Z(G369));
  INV_X1    g0513(.A(G330), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n268), .A2(new_n218), .A3(G13), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n715), .A2(KEYINPUT27), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(KEYINPUT27), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G213), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  XNOR2_X1  g0519(.A(KEYINPUT93), .B(G343), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n606), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n608), .A2(new_n722), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n592), .A2(new_n595), .B1(new_n602), .B2(new_n603), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n588), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n722), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n714), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n721), .B1(new_n648), .B2(new_n651), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n657), .A2(new_n728), .B1(new_n645), .B2(new_n721), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n721), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n724), .B2(new_n588), .ZN(new_n732));
  INV_X1    g0532(.A(new_n645), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n732), .A2(new_n656), .B1(new_n733), .B2(new_n721), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(G399));
  INV_X1    g0535(.A(new_n212), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G41), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n268), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n555), .A2(new_n553), .A3(new_n460), .ZN(new_n740));
  INV_X1    g0540(.A(new_n737), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n739), .A2(new_n740), .B1(new_n215), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n483), .A2(new_n598), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n597), .A2(new_n539), .A3(new_n652), .A4(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT94), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n539), .A2(new_n652), .A3(new_n744), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT94), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT30), .A4(new_n597), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n745), .A2(new_n746), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n483), .A2(new_n306), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n539), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n652), .A2(new_n525), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n753), .B(new_n754), .C1(new_n566), .C2(new_n585), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n747), .A2(new_n750), .A3(new_n751), .A4(new_n755), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n756), .A2(KEYINPUT31), .A3(new_n731), .ZN(new_n757));
  AOI21_X1  g0557(.A(KEYINPUT31), .B1(new_n756), .B2(new_n731), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n546), .A2(KEYINPUT80), .A3(new_n523), .ZN(new_n760));
  AOI21_X1  g0560(.A(KEYINPUT80), .B1(new_n546), .B2(new_n523), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n707), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n690), .A2(new_n691), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n762), .A2(new_n763), .A3(new_n731), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n658), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n714), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n710), .A2(new_n687), .ZN(new_n767));
  AOI21_X1  g0567(.A(KEYINPUT90), .B1(new_n693), .B2(new_n709), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n721), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT29), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT95), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g0573(.A(KEYINPUT95), .B(new_n707), .C1(new_n760), .C2(new_n761), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n773), .A2(new_n685), .A3(new_n686), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n692), .A2(KEYINPUT26), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n679), .B1(new_n708), .B2(new_n677), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(KEYINPUT29), .A3(new_n721), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n766), .B1(new_n771), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n743), .B1(new_n781), .B2(G1), .ZN(G364));
  INV_X1    g0582(.A(new_n727), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n218), .A2(G13), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G45), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT96), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n739), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n723), .A2(new_n714), .A3(new_n726), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n783), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n723), .A2(new_n726), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n736), .A2(new_n286), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G355), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G116), .B2(new_n212), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n242), .A2(G45), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n736), .A2(new_n290), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n473), .B2(new_n216), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n797), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n217), .B1(G20), .B2(new_n279), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n793), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n787), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n362), .A2(G179), .A3(G200), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n218), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n454), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n362), .A2(new_n317), .ZN(new_n810));
  NAND2_X1  g0610(.A1(G20), .A2(G179), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n286), .B(new_n809), .C1(G50), .C2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n218), .A2(G179), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n811), .A2(new_n362), .A3(G200), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(G87), .B1(G58), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G190), .A2(G200), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n812), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n815), .B(new_n820), .C1(new_n207), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n317), .A2(G190), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n816), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT98), .Z(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G107), .ZN(new_n827));
  XOR2_X1   g0627(.A(KEYINPUT97), .B(G159), .Z(new_n828));
  NAND2_X1  g0628(.A1(new_n816), .A2(new_n821), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT32), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n824), .A2(new_n812), .A3(KEYINPUT99), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT99), .B1(new_n824), .B2(new_n812), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n827), .B(new_n831), .C1(new_n329), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n826), .A2(G283), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n290), .B1(G322), .B2(new_n819), .ZN(new_n837));
  INV_X1    g0637(.A(G303), .ZN(new_n838));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n817), .A2(new_n838), .B1(new_n822), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n829), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(G329), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n834), .ZN(new_n843));
  XNOR2_X1  g0643(.A(KEYINPUT33), .B(G317), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n836), .A2(new_n837), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n808), .ZN(new_n847));
  XNOR2_X1  g0647(.A(KEYINPUT100), .B(G326), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n847), .A2(G294), .B1(new_n814), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT101), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n823), .A2(new_n835), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n806), .B1(new_n851), .B2(new_n803), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n794), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n790), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  NOR2_X1   g0655(.A1(new_n409), .A2(new_n731), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n404), .A2(new_n731), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n412), .A2(new_n857), .B1(new_n405), .B2(new_n408), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n791), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n803), .A2(new_n791), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n787), .B1(G77), .B2(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT102), .Z(new_n863));
  AOI211_X1 g0663(.A(new_n290), .B(new_n809), .C1(G303), .C2(new_n814), .ZN(new_n864));
  INV_X1    g0664(.A(new_n819), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n865), .A2(new_n611), .B1(new_n817), .B2(new_n510), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n829), .A2(new_n839), .B1(new_n822), .B2(new_n553), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n826), .A2(G87), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n843), .A2(G283), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n864), .A2(new_n868), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n822), .ZN(new_n872));
  INV_X1    g0672(.A(new_n828), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n872), .A2(new_n873), .B1(new_n814), .B2(G137), .ZN(new_n874));
  INV_X1    g0674(.A(G143), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n874), .B1(new_n875), .B2(new_n865), .C1(new_n262), .C2(new_n834), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT34), .Z(new_n877));
  NAND2_X1  g0677(.A1(new_n826), .A2(G68), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n290), .B1(new_n817), .B2(new_n275), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(G132), .B2(new_n841), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n878), .B(new_n880), .C1(new_n250), .C2(new_n808), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n871), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n863), .B1(new_n882), .B2(new_n803), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n859), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n856), .A2(new_n858), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n711), .B2(new_n721), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n413), .A2(new_n731), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n711), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n787), .B1(new_n888), .B2(new_n766), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT103), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n888), .A2(new_n766), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n889), .A2(new_n890), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n884), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(G384));
  OR2_X1    g0696(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(G116), .A3(new_n219), .A4(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT36), .Z(new_n900));
  OR3_X1    g0700(.A1(new_n215), .A2(new_n207), .A3(new_n330), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n202), .A2(G68), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n268), .B(G13), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n383), .A2(new_n384), .A3(new_n379), .ZN(new_n906));
  XOR2_X1   g0706(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n384), .B2(new_n719), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n361), .A2(new_n906), .A3(new_n908), .A4(new_n366), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n384), .A2(new_n719), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT105), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n384), .A2(new_n913), .A3(new_n719), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n915), .A2(new_n361), .A3(new_n366), .A4(new_n661), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n910), .B1(new_n916), .B2(KEYINPUT37), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n380), .A2(new_n385), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n915), .B1(new_n669), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n905), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n361), .A2(new_n366), .A3(new_n661), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n913), .B1(new_n384), .B2(new_n719), .ZN(new_n922));
  AOI211_X1 g0722(.A(KEYINPUT105), .B(new_n718), .C1(new_n340), .C2(new_n343), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT37), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n909), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(KEYINPUT38), .C1(new_n388), .C2(new_n915), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n920), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n756), .A2(new_n731), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT31), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n756), .A2(KEYINPUT31), .A3(new_n731), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n724), .A2(new_n656), .A3(new_n588), .A4(new_n607), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n549), .A2(new_n550), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n934), .A2(new_n504), .A3(new_n707), .A4(new_n721), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n931), .B(new_n932), .C1(new_n933), .C2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n426), .A2(new_n731), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT104), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n446), .A2(new_n938), .A3(new_n449), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n446), .A2(KEYINPUT104), .A3(new_n449), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n443), .A2(new_n445), .A3(new_n937), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n937), .A2(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n936), .A2(new_n885), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT40), .B1(new_n928), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n911), .B1(new_n669), .B2(new_n664), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n661), .A2(new_n911), .A3(new_n359), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n907), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n909), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n905), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n927), .A2(new_n950), .A3(KEYINPUT107), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT107), .B1(new_n927), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND4_X1   g0753(.A1(KEYINPUT40), .A2(new_n936), .A3(new_n885), .A4(new_n942), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n944), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n452), .A2(new_n936), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n957), .A2(new_n958), .A3(new_n714), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n664), .A2(new_n719), .ZN(new_n960));
  INV_X1    g0760(.A(new_n942), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n887), .B1(new_n767), .B2(new_n768), .ZN(new_n962));
  INV_X1    g0762(.A(new_n856), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n960), .B1(new_n964), .B2(new_n928), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT39), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n917), .A2(new_n919), .A3(new_n905), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(new_n664), .A3(new_n386), .ZN(new_n969));
  INV_X1    g0769(.A(new_n911), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT38), .B1(new_n971), .B2(new_n948), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n966), .B1(new_n967), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n446), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n721), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n920), .A2(new_n927), .A3(KEYINPUT39), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n965), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n771), .A2(new_n452), .A3(new_n780), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n674), .A2(new_n675), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n979), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n959), .A2(new_n984), .B1(new_n268), .B2(new_n784), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n959), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n904), .B1(new_n985), .B2(new_n986), .ZN(G367));
  INV_X1    g0787(.A(KEYINPUT110), .ZN(new_n988));
  INV_X1    g0788(.A(new_n730), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n773), .B(new_n774), .C1(new_n523), .C2(new_n721), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n544), .A2(new_n731), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n988), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n992), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n730), .A2(new_n994), .A3(KEYINPUT110), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n721), .B1(new_n496), .B2(new_n499), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n694), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n680), .B2(new_n997), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(KEYINPUT109), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n993), .A2(new_n995), .B1(KEYINPUT109), .B2(new_n1000), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT108), .Z(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT109), .B2(new_n1000), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n992), .A2(new_n656), .A3(new_n732), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT42), .Z(new_n1010));
  OR2_X1    g0810(.A1(new_n990), .A2(new_n645), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n707), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n721), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1008), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1004), .B(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n737), .B(KEYINPUT41), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n992), .A2(new_n734), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT45), .Z(new_n1018));
  NOR2_X1   g0818(.A1(new_n992), .A2(new_n734), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT44), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n989), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n732), .A2(new_n656), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n729), .B2(new_n732), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n727), .B(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1018), .A2(new_n730), .A3(new_n1020), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n781), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1016), .B1(new_n1027), .B2(new_n781), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n786), .A2(new_n268), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1015), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n238), .A2(new_n799), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n805), .B1(new_n736), .B2(new_n468), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n788), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n793), .ZN(new_n1035));
  INV_X1    g0835(.A(G317), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n813), .A2(new_n839), .B1(new_n829), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n286), .B1(new_n865), .B2(new_n838), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n825), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1037), .B(new_n1038), .C1(new_n513), .C2(new_n1039), .ZN(new_n1040));
  OR3_X1    g0840(.A1(new_n817), .A2(KEYINPUT46), .A3(new_n553), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT46), .B1(new_n817), .B2(new_n553), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n843), .A2(G294), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(G283), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n808), .A2(new_n510), .B1(new_n822), .B2(new_n1044), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT111), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(KEYINPUT111), .ZN(new_n1047));
  AND4_X1   g0847(.A1(new_n1040), .A2(new_n1043), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n834), .A2(new_n828), .B1(new_n202), .B2(new_n822), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT113), .Z(new_n1050));
  INV_X1    g0850(.A(G137), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n813), .A2(new_n875), .B1(new_n829), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G58), .B2(new_n818), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n808), .A2(new_n329), .B1(new_n865), .B2(new_n262), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(KEYINPUT112), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n286), .B1(new_n1039), .B2(G77), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1054), .A2(KEYINPUT112), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1048), .B1(new_n1050), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT47), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n803), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1034), .B1(new_n1035), .B2(new_n999), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1031), .A2(new_n1063), .ZN(G387));
  NAND2_X1  g0864(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n235), .A2(new_n473), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1066), .A2(new_n799), .B1(new_n740), .B2(new_n795), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n253), .A2(new_n275), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT50), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n473), .B1(new_n329), .B2(new_n207), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1069), .A2(new_n740), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n510), .B2(new_n736), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n787), .B1(new_n1073), .B2(new_n805), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n808), .A2(new_n398), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n286), .B(new_n1075), .C1(G159), .C2(new_n814), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n865), .A2(new_n275), .B1(new_n829), .B2(new_n262), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n817), .A2(new_n207), .B1(new_n822), .B2(new_n329), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n843), .A2(new_n253), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n826), .A2(G97), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1076), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n814), .A2(G322), .B1(new_n872), .B2(G303), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n1036), .B2(new_n865), .C1(new_n839), .C2(new_n834), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT114), .Z(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1086), .A2(KEYINPUT48), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(KEYINPUT48), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n808), .A2(new_n1044), .B1(new_n817), .B2(new_n611), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT49), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n286), .B1(new_n825), .B2(new_n553), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n841), .B2(new_n848), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1090), .A2(KEYINPUT49), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1082), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1074), .B1(new_n1096), .B2(new_n803), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n729), .B2(new_n1035), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n781), .A2(new_n1025), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n737), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n781), .A2(new_n1025), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1065), .B(new_n1098), .C1(new_n1100), .C2(new_n1101), .ZN(G393));
  INV_X1    g0902(.A(new_n1026), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n730), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1103), .A2(new_n1104), .A3(new_n1029), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n994), .A2(new_n793), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n804), .B1(new_n212), .B2(new_n555), .C1(new_n245), .C2(new_n800), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n787), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G283), .A2(new_n818), .B1(new_n841), .B2(G322), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1109), .B(new_n286), .C1(new_n611), .C2(new_n822), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G116), .B2(new_n847), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1111), .B(new_n827), .C1(new_n838), .C2(new_n834), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n814), .A2(G317), .B1(G311), .B2(new_n819), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT52), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n1115), .A2(KEYINPUT115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(KEYINPUT115), .ZN(new_n1117));
  INV_X1    g0917(.A(G159), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n865), .A2(new_n1118), .B1(new_n813), .B2(new_n262), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT51), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n254), .A2(new_n822), .B1(new_n829), .B2(new_n875), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n808), .A2(new_n207), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n290), .B1(new_n817), .B2(new_n329), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n843), .A2(new_n203), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1120), .A2(new_n1124), .A3(new_n869), .A4(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1116), .A2(new_n1117), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1108), .B1(new_n1127), .B2(new_n803), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1105), .B1(new_n1106), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1099), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(new_n1027), .A3(new_n737), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(G390));
  AND3_X1   g0932(.A1(new_n920), .A2(new_n927), .A3(KEYINPUT39), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT39), .B1(new_n927), .B2(new_n950), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n791), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n808), .A2(new_n1118), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n286), .B(new_n1136), .C1(G125), .C2(new_n841), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n822), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G132), .B2(new_n819), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n814), .A2(G128), .B1(new_n1039), .B2(new_n203), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT53), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n817), .B2(new_n262), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n818), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n843), .A2(G137), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1137), .A2(new_n1140), .A3(new_n1141), .A4(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n290), .B(new_n1122), .C1(G87), .C2(new_n818), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n865), .A2(new_n553), .B1(new_n822), .B2(new_n555), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n813), .A2(new_n1044), .B1(new_n829), .B2(new_n611), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n843), .A2(G107), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1147), .A2(new_n878), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1062), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n788), .B(new_n1153), .C1(new_n254), .C2(new_n860), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1135), .A2(new_n1154), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n731), .B(new_n858), .C1(new_n775), .C2(new_n778), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n942), .B1(new_n1156), .B2(new_n856), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT107), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n967), .B2(new_n972), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n927), .A2(new_n950), .A3(KEYINPUT107), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1157), .A2(new_n1159), .A3(new_n975), .A4(new_n1160), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1133), .A2(new_n1134), .B1(new_n964), .B2(new_n976), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n936), .A2(new_n942), .A3(G330), .A4(new_n885), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1161), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1155), .B1(new_n1168), .B2(new_n1029), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n452), .A2(new_n766), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n980), .A2(new_n981), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n856), .B1(new_n711), .B2(new_n887), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n931), .A2(new_n932), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n935), .A2(new_n933), .ZN(new_n1175));
  OAI211_X1 g0975(.A(G330), .B(new_n885), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n961), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1173), .B1(new_n1177), .B2(new_n1164), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT116), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1156), .A2(new_n856), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n1164), .A3(new_n1177), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1172), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n741), .B1(new_n1168), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1173), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n942), .B1(new_n766), .B2(new_n885), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n1165), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT116), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n1182), .A3(new_n1180), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1166), .A2(new_n1167), .A3(new_n1191), .A4(new_n1172), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1169), .B1(new_n1186), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(G378));
  OAI22_X1  g0994(.A1(new_n825), .A2(new_n250), .B1(new_n829), .B2(new_n1044), .ZN(new_n1195));
  INV_X1    g0995(.A(G41), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n286), .C1(new_n817), .C2(new_n207), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(G68), .C2(new_n847), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n814), .A2(G116), .B1(new_n872), .B2(new_n468), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n510), .B2(new_n865), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1198), .B(new_n1201), .C1(new_n454), .C2(new_n834), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT58), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(G50), .B1(new_n256), .B2(new_n1196), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n290), .B2(G41), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1202), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1207), .B2(KEYINPUT58), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n256), .B(new_n1196), .C1(new_n828), .C2(new_n825), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n872), .A2(G137), .B1(G128), .B2(new_n819), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n817), .B2(new_n1138), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n847), .A2(G150), .B1(new_n814), .B2(G125), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT117), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(G132), .C2(new_n843), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT118), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1209), .B(new_n1216), .C1(G124), .C2(new_n841), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1204), .B(new_n1208), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n787), .B1(new_n203), .B2(new_n861), .C1(new_n1219), .C2(new_n1062), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n278), .A2(new_n719), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT55), .Z(new_n1222));
  XNOR2_X1  g1022(.A(new_n322), .B(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1224));
  XNOR2_X1  g1024(.A(new_n1223), .B(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1220), .B1(new_n1225), .B2(new_n791), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1225), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n979), .B1(new_n955), .B2(G330), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n965), .A2(new_n978), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n928), .A2(new_n943), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT40), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1159), .A2(new_n1160), .A3(new_n954), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1233), .A3(G330), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1229), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1227), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1229), .A2(new_n1234), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n955), .A2(new_n979), .A3(G330), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1225), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1226), .B1(new_n1240), .B2(new_n1030), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1236), .A2(new_n1239), .B1(new_n1192), .B2(new_n1172), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n737), .B1(new_n1242), .B2(KEYINPUT57), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1237), .A2(new_n1238), .A3(new_n1225), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1225), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT57), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1161), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1164), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1171), .B1(new_n1250), .B2(new_n1191), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1246), .A2(new_n1247), .A3(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1241), .B1(new_n1243), .B2(new_n1252), .ZN(G375));
  NAND2_X1  g1053(.A1(new_n1191), .A2(new_n1030), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n788), .B1(new_n329), .B2(new_n860), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n814), .A2(G132), .ZN(new_n1256));
  XOR2_X1   g1056(.A(new_n1256), .B(KEYINPUT122), .Z(new_n1257));
  OAI221_X1 g1057(.A(new_n1257), .B1(new_n1051), .B2(new_n865), .C1(new_n834), .C2(new_n1138), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT123), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n290), .B1(new_n825), .B2(new_n250), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(G128), .A2(new_n841), .B1(new_n872), .B2(G150), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1118), .B2(new_n817), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1260), .B(new_n1262), .C1(G50), .C2(new_n847), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n813), .A2(new_n611), .B1(new_n822), .B2(new_n510), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n843), .B2(G116), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT121), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n290), .B1(G283), .B2(new_n819), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1267), .B1(new_n454), .B2(new_n817), .C1(new_n838), .C2(new_n829), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1075), .B(new_n1268), .C1(G77), .C2(new_n826), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1259), .A2(new_n1263), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1255), .B1(new_n1062), .B2(new_n1270), .C1(new_n942), .C2(new_n792), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1254), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1190), .A2(new_n1171), .A3(new_n1182), .A4(new_n1180), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1016), .B(KEYINPUT120), .Z(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1185), .A2(new_n1274), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1277), .ZN(G381));
  NOR2_X1   g1078(.A1(G375), .A2(G378), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OR4_X1    g1080(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1281));
  OR4_X1    g1081(.A1(G387), .A2(new_n1280), .A3(G381), .A4(new_n1281), .ZN(G407));
  INV_X1    g1082(.A(G213), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n720), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G407), .B(G213), .C1(new_n1280), .C2(new_n1285), .ZN(G409));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  OAI211_X1 g1087(.A(G378), .B(new_n1241), .C1(new_n1243), .C2(new_n1252), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1246), .A2(new_n1251), .A3(new_n1275), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1226), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1246), .B2(new_n1029), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1193), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT60), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1274), .A2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1188), .A2(new_n1165), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1181), .A2(new_n1296), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1297), .A2(KEYINPUT60), .A3(new_n1171), .A4(new_n1190), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1295), .A2(new_n737), .A3(new_n1298), .A4(new_n1185), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT124), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n741), .B1(new_n1191), .B2(new_n1172), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT124), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1301), .A2(new_n1295), .A3(new_n1302), .A4(new_n1298), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G384), .B1(new_n1304), .B2(new_n1273), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1272), .B(new_n895), .C1(new_n1300), .C2(new_n1303), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  AND4_X1   g1107(.A1(new_n1287), .A2(new_n1293), .A3(new_n1285), .A4(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1284), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1287), .B1(new_n1309), .B2(new_n1307), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  XOR2_X1   g1111(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1312));
  NAND2_X1  g1112(.A1(new_n1304), .A2(new_n1273), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n895), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1304), .A2(G384), .A3(new_n1273), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1284), .A2(G2897), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1316), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1318), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1312), .B1(new_n1320), .B2(new_n1309), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  OAI211_X1 g1123(.A(KEYINPUT127), .B(new_n1312), .C1(new_n1320), .C2(new_n1309), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1311), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1031), .A2(G390), .A3(new_n1063), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT125), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(G393), .B(new_n854), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(G387), .A2(new_n1131), .A3(new_n1129), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1326), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1331), .A2(KEYINPUT125), .A3(new_n1326), .A4(new_n1329), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1325), .A2(new_n1335), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(KEYINPUT61), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1309), .A2(KEYINPUT63), .A3(new_n1307), .ZN(new_n1338));
  OR2_X1    g1138(.A1(new_n1320), .A2(new_n1309), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1309), .A2(new_n1307), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT63), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1337), .A2(new_n1338), .A3(new_n1339), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1336), .A2(new_n1343), .ZN(G405));
  NAND2_X1  g1144(.A1(G375), .A2(new_n1193), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1335), .A2(new_n1288), .A3(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1288), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1333), .A2(new_n1347), .A3(new_n1334), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1346), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1349), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1346), .A2(new_n1307), .A3(new_n1348), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(G402));
endmodule


