

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n876) );
  OR2_X1 U556 ( .A1(n700), .A2(n699), .ZN(n705) );
  BUF_X1 U557 ( .A(n689), .Z(n730) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  NAND2_X1 U559 ( .A1(n760), .A2(n522), .ZN(n770) );
  NAND2_X1 U560 ( .A1(n583), .A2(n582), .ZN(n924) );
  NOR2_X2 U561 ( .A1(n538), .A2(n537), .ZN(G160) );
  AND2_X1 U562 ( .A1(n525), .A2(n929), .ZN(n522) );
  XOR2_X1 U563 ( .A(KEYINPUT14), .B(n580), .Z(n523) );
  OR2_X1 U564 ( .A1(n768), .A2(n767), .ZN(n524) );
  OR2_X1 U565 ( .A1(n758), .A2(n768), .ZN(n525) );
  NOR2_X1 U566 ( .A1(n751), .A2(n768), .ZN(n526) );
  AND2_X1 U567 ( .A1(n769), .A2(n524), .ZN(n527) );
  NOR2_X1 U568 ( .A1(n689), .A2(n688), .ZN(n691) );
  NOR2_X1 U569 ( .A1(n694), .A2(n924), .ZN(n698) );
  XNOR2_X1 U570 ( .A(n719), .B(KEYINPUT30), .ZN(n720) );
  XNOR2_X1 U571 ( .A(n721), .B(n720), .ZN(n722) );
  INV_X1 U572 ( .A(KEYINPUT31), .ZN(n726) );
  XNOR2_X1 U573 ( .A(n749), .B(KEYINPUT100), .ZN(n763) );
  NAND2_X1 U574 ( .A1(G8), .A2(n730), .ZN(n768) );
  AND2_X2 U575 ( .A1(n535), .A2(G2105), .ZN(n875) );
  NOR2_X2 U576 ( .A1(G2105), .A2(n535), .ZN(n872) );
  NOR2_X1 U577 ( .A1(G651), .A2(n624), .ZN(n653) );
  NOR2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n534) );
  AND2_X1 U579 ( .A1(G113), .A2(n876), .ZN(n528) );
  XNOR2_X1 U580 ( .A(n528), .B(KEYINPUT66), .ZN(n531) );
  NAND2_X1 U581 ( .A1(G125), .A2(n875), .ZN(n529) );
  XNOR2_X1 U582 ( .A(n529), .B(KEYINPUT65), .ZN(n530) );
  XOR2_X2 U583 ( .A(KEYINPUT17), .B(n532), .Z(n871) );
  NAND2_X1 U584 ( .A1(n871), .A2(G137), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n538) );
  INV_X1 U586 ( .A(G2104), .ZN(n535) );
  NAND2_X1 U587 ( .A1(G101), .A2(n872), .ZN(n536) );
  XNOR2_X1 U588 ( .A(KEYINPUT23), .B(n536), .ZN(n537) );
  NOR2_X2 U589 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U590 ( .A1(G89), .A2(n645), .ZN(n539) );
  XNOR2_X1 U591 ( .A(n539), .B(KEYINPUT70), .ZN(n540) );
  XNOR2_X1 U592 ( .A(n540), .B(KEYINPUT4), .ZN(n542) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n624) );
  INV_X1 U594 ( .A(G651), .ZN(n544) );
  NOR2_X1 U595 ( .A1(n624), .A2(n544), .ZN(n649) );
  NAND2_X1 U596 ( .A1(G76), .A2(n649), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U598 ( .A(n543), .B(KEYINPUT5), .ZN(n550) );
  NOR2_X1 U599 ( .A1(G543), .A2(n544), .ZN(n545) );
  XOR2_X2 U600 ( .A(KEYINPUT1), .B(n545), .Z(n646) );
  NAND2_X1 U601 ( .A1(G63), .A2(n646), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G51), .A2(n653), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U604 ( .A(KEYINPUT6), .B(n548), .Z(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U606 ( .A(n551), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U607 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U608 ( .A1(n875), .A2(G126), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n552), .B(KEYINPUT84), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G138), .A2(n871), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U612 ( .A1(G102), .A2(n872), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G114), .A2(n876), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U615 ( .A1(n558), .A2(n557), .ZN(G164) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U617 ( .A1(G64), .A2(n646), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G52), .A2(n653), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G90), .A2(n645), .ZN(n562) );
  NAND2_X1 U621 ( .A1(G77), .A2(n649), .ZN(n561) );
  NAND2_X1 U622 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U624 ( .A1(n565), .A2(n564), .ZN(G171) );
  INV_X1 U625 ( .A(G171), .ZN(G301) );
  NAND2_X1 U626 ( .A1(G65), .A2(n646), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G53), .A2(n653), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U629 ( .A1(G91), .A2(n645), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G78), .A2(n649), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n921) );
  INV_X1 U633 ( .A(n921), .ZN(G299) );
  INV_X1 U634 ( .A(G57), .ZN(G237) );
  INV_X1 U635 ( .A(G132), .ZN(G219) );
  INV_X1 U636 ( .A(G82), .ZN(G220) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U639 ( .A(G223), .ZN(n822) );
  NAND2_X1 U640 ( .A1(n822), .A2(G567), .ZN(n573) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  XNOR2_X1 U642 ( .A(KEYINPUT13), .B(KEYINPUT69), .ZN(n579) );
  NAND2_X1 U643 ( .A1(G81), .A2(n645), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT68), .ZN(n575) );
  XNOR2_X1 U645 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U646 ( .A1(G68), .A2(n649), .ZN(n576) );
  NAND2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U648 ( .A(n579), .B(n578), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n646), .A2(G56), .ZN(n580) );
  NOR2_X1 U650 ( .A1(n581), .A2(n523), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n653), .A2(G43), .ZN(n582) );
  INV_X1 U652 ( .A(G860), .ZN(n614) );
  OR2_X1 U653 ( .A1(n924), .A2(n614), .ZN(G153) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n592) );
  NAND2_X1 U655 ( .A1(G92), .A2(n645), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G79), .A2(n649), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G66), .A2(n646), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G54), .A2(n653), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U662 ( .A(KEYINPUT15), .B(n590), .Z(n896) );
  INV_X1 U663 ( .A(n896), .ZN(n917) );
  INV_X1 U664 ( .A(G868), .ZN(n665) );
  NAND2_X1 U665 ( .A1(n917), .A2(n665), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(G284) );
  NOR2_X1 U667 ( .A1(G286), .A2(n665), .ZN(n593) );
  XOR2_X1 U668 ( .A(KEYINPUT71), .B(n593), .Z(n595) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U670 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U671 ( .A1(n614), .A2(G559), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n596), .A2(n896), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(n917), .A2(n665), .ZN(n598) );
  XOR2_X1 U675 ( .A(KEYINPUT72), .B(n598), .Z(n599) );
  NOR2_X1 U676 ( .A1(G559), .A2(n599), .ZN(n601) );
  NOR2_X1 U677 ( .A1(G868), .A2(n924), .ZN(n600) );
  NOR2_X1 U678 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U679 ( .A1(G123), .A2(n875), .ZN(n602) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(n602), .Z(n603) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT73), .ZN(n605) );
  NAND2_X1 U682 ( .A1(G135), .A2(n871), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U684 ( .A(KEYINPUT74), .B(n606), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G99), .A2(n872), .ZN(n608) );
  NAND2_X1 U686 ( .A1(G111), .A2(n876), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n1002) );
  XNOR2_X1 U689 ( .A(G2096), .B(n1002), .ZN(n612) );
  INV_X1 U690 ( .A(G2100), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(G156) );
  NAND2_X1 U692 ( .A1(G559), .A2(n896), .ZN(n613) );
  XOR2_X1 U693 ( .A(n924), .B(n613), .Z(n662) );
  NAND2_X1 U694 ( .A1(n614), .A2(n662), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n653), .A2(G55), .ZN(n615) );
  XOR2_X1 U696 ( .A(KEYINPUT75), .B(n615), .Z(n617) );
  NAND2_X1 U697 ( .A1(n646), .A2(G67), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U699 ( .A(KEYINPUT76), .B(n618), .Z(n622) );
  NAND2_X1 U700 ( .A1(G93), .A2(n645), .ZN(n620) );
  NAND2_X1 U701 ( .A1(G80), .A2(n649), .ZN(n619) );
  AND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n664) );
  XNOR2_X1 U704 ( .A(n623), .B(n664), .ZN(G145) );
  NAND2_X1 U705 ( .A1(G49), .A2(n653), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G87), .A2(n624), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U708 ( .A1(n646), .A2(n627), .ZN(n630) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n628) );
  XOR2_X1 U710 ( .A(KEYINPUT77), .B(n628), .Z(n629) );
  NAND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U712 ( .A1(G60), .A2(n646), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G47), .A2(n653), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G85), .A2(n645), .ZN(n634) );
  NAND2_X1 U716 ( .A1(G72), .A2(n649), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U719 ( .A(n637), .B(KEYINPUT67), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G62), .A2(n646), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G50), .A2(n653), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U723 ( .A(KEYINPUT78), .B(n640), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G88), .A2(n645), .ZN(n642) );
  NAND2_X1 U725 ( .A1(G75), .A2(n649), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U727 ( .A1(n644), .A2(n643), .ZN(G166) );
  NAND2_X1 U728 ( .A1(G86), .A2(n645), .ZN(n648) );
  NAND2_X1 U729 ( .A1(G61), .A2(n646), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n649), .A2(G73), .ZN(n650) );
  XOR2_X1 U732 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n653), .A2(G48), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(G305) );
  XOR2_X1 U736 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n656) );
  XNOR2_X1 U737 ( .A(G288), .B(n656), .ZN(n657) );
  XOR2_X1 U738 ( .A(n664), .B(n657), .Z(n659) );
  XNOR2_X1 U739 ( .A(G290), .B(G166), .ZN(n658) );
  XNOR2_X1 U740 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n660), .B(G299), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n661), .B(G305), .ZN(n893) );
  XNOR2_X1 U743 ( .A(n662), .B(n893), .ZN(n663) );
  NAND2_X1 U744 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U748 ( .A(KEYINPUT80), .B(KEYINPUT20), .Z(n668) );
  XNOR2_X1 U749 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n670), .A2(G2090), .ZN(n671) );
  XOR2_X1 U751 ( .A(KEYINPUT21), .B(n671), .Z(n672) );
  XNOR2_X1 U752 ( .A(KEYINPUT81), .B(n672), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n674) );
  XNOR2_X1 U756 ( .A(KEYINPUT22), .B(n674), .ZN(n675) );
  NAND2_X1 U757 ( .A1(n675), .A2(G96), .ZN(n676) );
  NOR2_X1 U758 ( .A1(G218), .A2(n676), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT82), .B(n677), .Z(n829) );
  NAND2_X1 U760 ( .A1(n829), .A2(G2106), .ZN(n681) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n678) );
  NOR2_X1 U762 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U763 ( .A1(G108), .A2(n679), .ZN(n828) );
  NAND2_X1 U764 ( .A1(G567), .A2(n828), .ZN(n680) );
  NAND2_X1 U765 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U766 ( .A(KEYINPUT83), .B(n682), .ZN(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n684) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n683) );
  NOR2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n827) );
  NAND2_X1 U770 ( .A1(n827), .A2(G36), .ZN(G176) );
  XNOR2_X1 U771 ( .A(KEYINPUT85), .B(G166), .ZN(G303) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n771) );
  INV_X1 U773 ( .A(n771), .ZN(n685) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n772) );
  NAND2_X1 U775 ( .A1(n685), .A2(n772), .ZN(n689) );
  INV_X1 U776 ( .A(n730), .ZN(n712) );
  NOR2_X1 U777 ( .A1(n712), .A2(G1348), .ZN(n687) );
  NOR2_X1 U778 ( .A1(G2067), .A2(n730), .ZN(n686) );
  NOR2_X1 U779 ( .A1(n687), .A2(n686), .ZN(n696) );
  INV_X1 U780 ( .A(G1996), .ZN(n688) );
  XOR2_X1 U781 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n690) );
  XNOR2_X1 U782 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n730), .A2(G1341), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n698), .A2(n896), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U787 ( .A(KEYINPUT95), .B(n697), .ZN(n700) );
  NOR2_X1 U788 ( .A1(n896), .A2(n698), .ZN(n699) );
  NAND2_X1 U789 ( .A1(n712), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U790 ( .A(n701), .B(KEYINPUT27), .ZN(n703) );
  INV_X1 U791 ( .A(G1956), .ZN(n922) );
  NOR2_X1 U792 ( .A1(n922), .A2(n712), .ZN(n702) );
  NOR2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n921), .A2(n706), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n710) );
  NOR2_X1 U796 ( .A1(n921), .A2(n706), .ZN(n708) );
  XNOR2_X1 U797 ( .A(KEYINPUT28), .B(KEYINPUT93), .ZN(n707) );
  XNOR2_X1 U798 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U800 ( .A(KEYINPUT29), .B(n711), .Z(n716) );
  OR2_X1 U801 ( .A1(n712), .A2(G1961), .ZN(n714) );
  XNOR2_X1 U802 ( .A(KEYINPUT25), .B(G2078), .ZN(n971) );
  NAND2_X1 U803 ( .A1(n712), .A2(n971), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n723) );
  NAND2_X1 U805 ( .A1(n723), .A2(G171), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n729) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n768), .ZN(n743) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n730), .ZN(n740) );
  NOR2_X1 U809 ( .A1(n743), .A2(n740), .ZN(n717) );
  XNOR2_X1 U810 ( .A(n717), .B(KEYINPUT96), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n718), .A2(G8), .ZN(n721) );
  INV_X1 U812 ( .A(KEYINPUT97), .ZN(n719) );
  NOR2_X1 U813 ( .A1(n722), .A2(G168), .ZN(n725) );
  NOR2_X1 U814 ( .A1(G171), .A2(n723), .ZN(n724) );
  NOR2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n727) );
  XNOR2_X1 U816 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U817 ( .A1(n729), .A2(n728), .ZN(n742) );
  NAND2_X1 U818 ( .A1(n742), .A2(G286), .ZN(n737) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n730), .ZN(n731) );
  XOR2_X1 U820 ( .A(KEYINPUT98), .B(n731), .Z(n732) );
  NAND2_X1 U821 ( .A1(n732), .A2(G303), .ZN(n734) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n768), .ZN(n733) );
  NOR2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U824 ( .A(n735), .B(KEYINPUT99), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n738), .A2(G8), .ZN(n739) );
  XNOR2_X1 U827 ( .A(n739), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U828 ( .A1(G8), .A2(n740), .ZN(n741) );
  XNOR2_X1 U829 ( .A(KEYINPUT92), .B(n741), .ZN(n746) );
  INV_X1 U830 ( .A(n742), .ZN(n744) );
  NOR2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U832 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U833 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n757) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U836 ( .A1(n757), .A2(n750), .ZN(n933) );
  NAND2_X1 U837 ( .A1(n763), .A2(n933), .ZN(n752) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n932) );
  INV_X1 U839 ( .A(n932), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n526), .ZN(n754) );
  INV_X1 U841 ( .A(KEYINPUT64), .ZN(n753) );
  XNOR2_X1 U842 ( .A(n754), .B(n753), .ZN(n755) );
  NOR2_X1 U843 ( .A1(KEYINPUT33), .A2(n755), .ZN(n756) );
  XNOR2_X1 U844 ( .A(n756), .B(KEYINPUT101), .ZN(n760) );
  NAND2_X1 U845 ( .A1(n757), .A2(KEYINPUT33), .ZN(n758) );
  XOR2_X1 U846 ( .A(G1981), .B(KEYINPUT102), .Z(n759) );
  XNOR2_X1 U847 ( .A(G305), .B(n759), .ZN(n929) );
  NOR2_X1 U848 ( .A1(G2090), .A2(G303), .ZN(n761) );
  NAND2_X1 U849 ( .A1(G8), .A2(n761), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U851 ( .A(KEYINPUT103), .B(n764), .Z(n765) );
  NAND2_X1 U852 ( .A1(n768), .A2(n765), .ZN(n769) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XOR2_X1 U854 ( .A(n766), .B(KEYINPUT24), .Z(n767) );
  NAND2_X1 U855 ( .A1(n770), .A2(n527), .ZN(n806) );
  XNOR2_X1 U856 ( .A(G1986), .B(G290), .ZN(n926) );
  NOR2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n817) );
  NAND2_X1 U858 ( .A1(n926), .A2(n817), .ZN(n804) );
  XNOR2_X1 U859 ( .A(KEYINPUT87), .B(KEYINPUT36), .ZN(n783) );
  NAND2_X1 U860 ( .A1(G128), .A2(n875), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G116), .A2(n876), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U863 ( .A(KEYINPUT35), .B(n775), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G140), .A2(n871), .ZN(n777) );
  NAND2_X1 U865 ( .A1(G104), .A2(n872), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n779) );
  XOR2_X1 U867 ( .A(KEYINPUT86), .B(KEYINPUT34), .Z(n778) );
  XNOR2_X1 U868 ( .A(n779), .B(n778), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U870 ( .A(n783), .B(n782), .ZN(n889) );
  XNOR2_X1 U871 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NOR2_X1 U872 ( .A1(n889), .A2(n815), .ZN(n994) );
  NAND2_X1 U873 ( .A1(n817), .A2(n994), .ZN(n784) );
  XNOR2_X1 U874 ( .A(KEYINPUT88), .B(n784), .ZN(n813) );
  XNOR2_X1 U875 ( .A(KEYINPUT89), .B(G1991), .ZN(n970) );
  NAND2_X1 U876 ( .A1(G119), .A2(n875), .ZN(n786) );
  NAND2_X1 U877 ( .A1(G131), .A2(n871), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G95), .A2(n872), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G107), .A2(n876), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n868) );
  OR2_X1 U883 ( .A1(n970), .A2(n868), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G117), .A2(n876), .ZN(n797) );
  NAND2_X1 U885 ( .A1(G129), .A2(n875), .ZN(n792) );
  NAND2_X1 U886 ( .A1(G141), .A2(n871), .ZN(n791) );
  NAND2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n872), .A2(G105), .ZN(n793) );
  XOR2_X1 U889 ( .A(KEYINPUT38), .B(n793), .Z(n794) );
  NOR2_X1 U890 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U892 ( .A(n798), .B(KEYINPUT90), .ZN(n884) );
  NAND2_X1 U893 ( .A1(G1996), .A2(n884), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n993) );
  NAND2_X1 U895 ( .A1(n993), .A2(n817), .ZN(n801) );
  XNOR2_X1 U896 ( .A(n801), .B(KEYINPUT91), .ZN(n810) );
  INV_X1 U897 ( .A(n810), .ZN(n802) );
  AND2_X1 U898 ( .A1(n813), .A2(n802), .ZN(n803) );
  AND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n820) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n884), .ZN(n998) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n970), .A2(n868), .ZN(n807) );
  XOR2_X1 U904 ( .A(KEYINPUT104), .B(n807), .Z(n1001) );
  NOR2_X1 U905 ( .A1(n808), .A2(n1001), .ZN(n809) );
  NOR2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n998), .A2(n811), .ZN(n812) );
  XNOR2_X1 U908 ( .A(KEYINPUT39), .B(n812), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n889), .A2(n815), .ZN(n996) );
  NAND2_X1 U911 ( .A1(n816), .A2(n996), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U914 ( .A(KEYINPUT40), .B(n821), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n822), .ZN(G217) );
  NAND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n824) );
  INV_X1 U917 ( .A(G661), .ZN(n823) );
  NOR2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n825), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n829), .A2(n828), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XOR2_X1 U928 ( .A(G2096), .B(KEYINPUT106), .Z(n831) );
  XNOR2_X1 U929 ( .A(G2090), .B(KEYINPUT43), .ZN(n830) );
  XNOR2_X1 U930 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U931 ( .A(n832), .B(KEYINPUT42), .Z(n834) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2072), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U934 ( .A(G2678), .B(G2100), .Z(n836) );
  XNOR2_X1 U935 ( .A(G2078), .B(G2084), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U938 ( .A(G1976), .B(G1956), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1996), .B(G1961), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U941 ( .A(G1981), .B(G1971), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1966), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U944 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U945 ( .A(G2474), .B(KEYINPUT107), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n848) );
  XOR2_X1 U947 ( .A(G1991), .B(KEYINPUT41), .Z(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U949 ( .A1(n875), .A2(G124), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U951 ( .A1(G136), .A2(n871), .ZN(n850) );
  NAND2_X1 U952 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U953 ( .A(KEYINPUT108), .B(n852), .ZN(n856) );
  NAND2_X1 U954 ( .A1(G100), .A2(n872), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G112), .A2(n876), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U957 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U958 ( .A1(G142), .A2(n871), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G106), .A2(n872), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n859), .B(KEYINPUT45), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G130), .A2(n875), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G118), .A2(n876), .ZN(n862) );
  XNOR2_X1 U965 ( .A(KEYINPUT109), .B(n862), .ZN(n863) );
  NOR2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n888) );
  XOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT110), .Z(n866) );
  XNOR2_X1 U968 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U970 ( .A(n867), .B(G162), .Z(n870) );
  XNOR2_X1 U971 ( .A(G160), .B(n868), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n883) );
  NAND2_X1 U973 ( .A1(G139), .A2(n871), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G103), .A2(n872), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n882) );
  NAND2_X1 U976 ( .A1(G127), .A2(n875), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G115), .A2(n876), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U979 ( .A(KEYINPUT47), .B(n879), .ZN(n880) );
  XNOR2_X1 U980 ( .A(KEYINPUT111), .B(n880), .ZN(n881) );
  NOR2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n1004) );
  XOR2_X1 U982 ( .A(n883), .B(n1004), .Z(n886) );
  XNOR2_X1 U983 ( .A(G164), .B(n884), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n891) );
  XNOR2_X1 U986 ( .A(n889), .B(n1002), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U988 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U989 ( .A(n893), .B(G301), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n894), .B(n924), .ZN(n895) );
  XOR2_X1 U991 ( .A(n895), .B(KEYINPUT114), .Z(n898) );
  XNOR2_X1 U992 ( .A(n896), .B(KEYINPUT113), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U994 ( .A(G286), .B(n899), .Z(n900) );
  NOR2_X1 U995 ( .A1(G37), .A2(n900), .ZN(G397) );
  XOR2_X1 U996 ( .A(G2451), .B(G2430), .Z(n902) );
  XNOR2_X1 U997 ( .A(G2438), .B(G2443), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n908) );
  XOR2_X1 U999 ( .A(G2435), .B(G2454), .Z(n904) );
  XNOR2_X1 U1000 ( .A(G1341), .B(G1348), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1002 ( .A(G2446), .B(G2427), .Z(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1004 ( .A(n908), .B(n907), .Z(n909) );
  NAND2_X1 U1005 ( .A1(G14), .A2(n909), .ZN(n916) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n916), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n910) );
  XOR2_X1 U1008 ( .A(KEYINPUT115), .B(n910), .Z(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(KEYINPUT49), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(n916), .ZN(G401) );
  XNOR2_X1 U1016 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1026) );
  XNOR2_X1 U1017 ( .A(KEYINPUT56), .B(G16), .ZN(n944) );
  XNOR2_X1 U1018 ( .A(G301), .B(G1961), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n917), .B(G1348), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(KEYINPUT122), .B(n920), .ZN(n942) );
  XNOR2_X1 U1022 ( .A(n922), .B(n921), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(n923), .B(KEYINPUT123), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(G1341), .B(n924), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n940) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G168), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n931), .B(KEYINPUT57), .ZN(n938) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n935) );
  AND2_X1 U1031 ( .A1(G303), .A2(G1971), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(n936), .B(KEYINPUT124), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n1024) );
  XOR2_X1 U1038 ( .A(G1976), .B(G23), .Z(n946) );
  XOR2_X1 U1039 ( .A(G1971), .B(G22), .Z(n945) );
  NAND2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G24), .B(G1986), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1043 ( .A(KEYINPUT58), .B(n949), .Z(n965) );
  XNOR2_X1 U1044 ( .A(G1348), .B(KEYINPUT59), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(n950), .B(G4), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G1956), .B(G20), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G6), .B(G1981), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1050 ( .A(KEYINPUT125), .B(G1341), .Z(n955) );
  XNOR2_X1 U1051 ( .A(G19), .B(n955), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(KEYINPUT60), .B(n958), .ZN(n960) );
  XOR2_X1 U1054 ( .A(G1961), .B(G5), .Z(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(G21), .B(G1966), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1058 ( .A(KEYINPUT126), .B(n963), .Z(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT61), .B(n966), .ZN(n968) );
  INV_X1 U1061 ( .A(G16), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n969), .A2(G11), .ZN(n1022) );
  XOR2_X1 U1064 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n983) );
  XOR2_X1 U1065 ( .A(n970), .B(G25), .Z(n980) );
  XNOR2_X1 U1066 ( .A(G27), .B(n971), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(G2067), .B(G26), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(G1996), .B(G32), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(G33), .B(G2072), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(KEYINPUT119), .B(n978), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n981), .A2(G28), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(n983), .B(n982), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(G35), .B(G2090), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1079 ( .A(G2084), .B(KEYINPUT54), .Z(n986) );
  XNOR2_X1 U1080 ( .A(G34), .B(n986), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT121), .B(n989), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(G29), .A2(n990), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(n991), .B(KEYINPUT55), .ZN(n1020) );
  XOR2_X1 U1085 ( .A(G160), .B(G2084), .Z(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n1016) );
  INV_X1 U1087 ( .A(n994), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n1014) );
  XOR2_X1 U1089 ( .A(G2090), .B(G162), .Z(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(KEYINPUT117), .B(n999), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(n1000), .B(KEYINPUT51), .ZN(n1012) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1094 ( .A(KEYINPUT116), .B(n1003), .Z(n1010) );
  XOR2_X1 U1095 ( .A(G164), .B(G2078), .Z(n1007) );
  XOR2_X1 U1096 ( .A(n1004), .B(KEYINPUT118), .Z(n1005) );
  XNOR2_X1 U1097 ( .A(G2072), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(KEYINPUT50), .B(n1008), .Z(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT52), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(G29), .A2(n1018), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(n1026), .B(n1025), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

