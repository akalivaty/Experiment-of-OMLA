//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G78gat), .B(G106gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT31), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(G141gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT79), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT2), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G155gat), .ZN(new_n219));
  INV_X1    g018(.A(G162gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n221), .A2(new_n216), .ZN(new_n222));
  OR3_X1    g021(.A1(new_n210), .A2(KEYINPUT80), .A3(G148gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n214), .A2(KEYINPUT80), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(new_n213), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n216), .B1(new_n221), .B2(KEYINPUT2), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n218), .A2(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G197gat), .B(G204gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT22), .ZN(new_n229));
  INV_X1    g028(.A(G211gat), .ZN(new_n230));
  INV_X1    g029(.A(G218gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n228), .A3(new_n232), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n227), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n238), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT29), .B1(new_n227), .B2(new_n241), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(KEYINPUT84), .ZN(new_n246));
  XNOR2_X1  g045(.A(G141gat), .B(G148gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n217), .B1(new_n247), .B2(KEYINPUT79), .ZN(new_n248));
  INV_X1    g047(.A(new_n215), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n222), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n225), .A2(new_n226), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n241), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n239), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT84), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n243), .B1(new_n246), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G228gat), .ZN(new_n257));
  INV_X1    g056(.A(G233gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n238), .B1(new_n252), .B2(new_n239), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n261), .A2(new_n242), .A3(new_n259), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n206), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  AOI211_X1 g063(.A(new_n205), .B(new_n262), .C1(new_n256), .C2(new_n259), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n203), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n238), .B1(new_n253), .B2(new_n254), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n245), .A2(KEYINPUT84), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n242), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n259), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n263), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n205), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n260), .A2(new_n263), .A3(new_n206), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n202), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT78), .ZN(new_n276));
  NAND2_X1  g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT26), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT27), .B(G183gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(G190gat), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n288));
  AOI21_X1  g087(.A(G190gat), .B1(new_n288), .B2(KEYINPUT27), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT27), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT28), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n277), .B(new_n283), .C1(new_n287), .C2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT23), .B1(new_n278), .B2(KEYINPUT65), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n295), .B(new_n296), .C1(G169gat), .C2(G176gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n297), .A3(new_n281), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT25), .ZN(new_n300));
  NAND3_X1  g099(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  AND2_X1   g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(KEYINPUT24), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n299), .B(new_n300), .C1(new_n305), .C2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n306), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(KEYINPUT24), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT24), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT66), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n277), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n310), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(KEYINPUT66), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n311), .A2(KEYINPUT24), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n307), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(KEYINPUT68), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n320), .A2(KEYINPUT67), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n298), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n293), .B(new_n309), .C1(new_n325), .C2(new_n300), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n326), .A2(new_n239), .B1(G226gat), .B2(G233gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT66), .B(KEYINPUT24), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n316), .B1(new_n328), .B2(new_n307), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n322), .A2(new_n323), .ZN(new_n330));
  OAI211_X1 g129(.A(KEYINPUT67), .B(new_n277), .C1(new_n312), .C2(new_n314), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .A4(new_n306), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n300), .B1(new_n332), .B2(new_n299), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n289), .A2(new_n291), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n334), .A2(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n283), .A2(new_n277), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n308), .B1(new_n304), .B2(new_n303), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n294), .A2(new_n300), .A3(new_n297), .A4(new_n281), .ZN(new_n338));
  OAI22_X1  g137(.A1(new_n335), .A2(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G226gat), .A2(G233gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n327), .A2(new_n342), .A3(new_n244), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n340), .B2(KEYINPUT29), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n326), .A2(G226gat), .A3(G233gat), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n238), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n276), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n244), .B1(new_n327), .B2(new_n342), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n345), .A3(new_n238), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT78), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G8gat), .B(G36gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(G64gat), .ZN(new_n352));
  INV_X1    g151(.A(G92gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n348), .A2(new_n349), .A3(new_n354), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT30), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n348), .A2(KEYINPUT30), .A3(new_n349), .A4(new_n354), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n275), .A2(new_n361), .A3(KEYINPUT35), .ZN(new_n362));
  INV_X1    g161(.A(G127gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G134gat), .ZN(new_n364));
  INV_X1    g163(.A(G134gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G127gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n366), .A3(KEYINPUT70), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(KEYINPUT70), .B2(new_n364), .ZN(new_n368));
  INV_X1    g167(.A(G113gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G120gat), .ZN(new_n370));
  INV_X1    g169(.A(G120gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G113gat), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT1), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n365), .A2(G127gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n363), .A2(G134gat), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT72), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT72), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n364), .A2(new_n366), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT71), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n371), .ZN(new_n382));
  NAND2_X1  g181(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(G113gat), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT1), .B1(new_n384), .B2(new_n370), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT73), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n380), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n374), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT74), .B1(new_n340), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n340), .A2(new_n390), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n340), .A2(KEYINPUT74), .A3(new_n390), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n393), .A2(KEYINPUT34), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT74), .ZN(new_n397));
  INV_X1    g196(.A(new_n374), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n380), .A2(new_n385), .A3(new_n388), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n388), .B1(new_n380), .B2(new_n385), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n326), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n326), .A2(new_n401), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n402), .A2(new_n395), .A3(new_n394), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT34), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n396), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT32), .ZN(new_n408));
  XNOR2_X1  g207(.A(G15gat), .B(G43gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(G71gat), .B(G99gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(KEYINPUT75), .B(KEYINPUT33), .Z(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n408), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n402), .A2(new_n395), .A3(new_n403), .ZN(new_n417));
  INV_X1    g216(.A(new_n394), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n417), .A2(new_n418), .B1(new_n408), .B2(new_n414), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n407), .B(new_n420), .C1(new_n421), .C2(new_n411), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n404), .B(KEYINPUT34), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(new_n418), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n414), .A2(new_n408), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n411), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n426), .B2(new_n419), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n427), .A3(KEYINPUT77), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT77), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n423), .B(new_n429), .C1(new_n426), .C2(new_n419), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n398), .B(new_n227), .C1(new_n399), .C2(new_n400), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT4), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n387), .A2(new_n389), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n398), .A4(new_n227), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n227), .B(KEYINPUT3), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n401), .ZN(new_n439));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n432), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT5), .ZN(new_n444));
  INV_X1    g243(.A(new_n227), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n401), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n432), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n444), .B1(new_n447), .B2(new_n441), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n433), .A2(new_n436), .B1(new_n438), .B2(new_n401), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n441), .A2(KEYINPUT5), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n443), .A2(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XOR2_X1   g250(.A(G57gat), .B(G85gat), .Z(new_n452));
  XNOR2_X1  g251(.A(G1gat), .B(G29gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n451), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n448), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n449), .A2(new_n450), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n456), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n457), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n451), .B2(new_n456), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n362), .A2(new_n431), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT76), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n424), .A2(new_n425), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n419), .B1(new_n470), .B2(new_n412), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n471), .B2(new_n407), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n423), .B(KEYINPUT76), .C1(new_n426), .C2(new_n419), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n422), .A2(new_n266), .A3(new_n274), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT87), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n422), .A2(new_n274), .A3(new_n266), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n472), .A4(new_n473), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n461), .A2(KEYINPUT83), .A3(new_n462), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT83), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n451), .B2(new_n456), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n482), .A3(new_n465), .ZN(new_n483));
  INV_X1    g282(.A(new_n458), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n361), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n476), .A2(new_n479), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n468), .B1(new_n486), .B2(KEYINPUT35), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n348), .A2(KEYINPUT78), .A3(new_n349), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT78), .B1(new_n348), .B2(new_n349), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT37), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT38), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n348), .A2(new_n349), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n491), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n354), .B1(KEYINPUT37), .B2(new_n491), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n492), .B(new_n491), .C1(KEYINPUT37), .C2(new_n354), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n490), .A2(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n275), .B1(new_n466), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n488), .A2(new_n489), .A3(new_n354), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n359), .A2(new_n360), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n463), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(KEYINPUT40), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n440), .B1(new_n437), .B2(new_n439), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n446), .A2(new_n440), .A3(new_n432), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT39), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n456), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n449), .A2(KEYINPUT39), .A3(new_n440), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n506), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT39), .B(new_n508), .C1(new_n449), .C2(new_n440), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT39), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n507), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n506), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n513), .A2(new_n515), .A3(new_n456), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n501), .B1(new_n504), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n512), .A2(new_n517), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n520), .A2(KEYINPUT86), .A3(new_n463), .A4(new_n361), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n500), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n483), .A2(new_n484), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n275), .B1(new_n523), .B2(new_n361), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n472), .A2(KEYINPUT36), .A3(new_n422), .A4(new_n473), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n431), .B2(KEYINPUT36), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n487), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G113gat), .B(G141gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT11), .ZN(new_n530));
  INV_X1    g329(.A(G169gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G197gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT12), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536));
  INV_X1    g335(.A(G1gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT16), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(G1gat), .B2(new_n536), .ZN(new_n540));
  INV_X1    g339(.A(G8gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(new_n536), .B2(G1gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT91), .ZN(new_n545));
  OAI221_X1 g344(.A(new_n539), .B1(new_n542), .B2(G8gat), .C1(G1gat), .C2(new_n536), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n550));
  INV_X1    g349(.A(G29gat), .ZN(new_n551));
  INV_X1    g350(.A(G36gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT88), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT88), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n555), .A2(new_n550), .A3(new_n551), .A4(new_n552), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G29gat), .A2(G36gat), .ZN(new_n559));
  INV_X1    g358(.A(G43gat), .ZN(new_n560));
  INV_X1    g359(.A(G50gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G43gat), .A2(G50gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT15), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n566), .A3(new_n563), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n558), .A2(new_n559), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n553), .A2(new_n557), .B1(G29gat), .B2(G36gat), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT89), .B(KEYINPUT17), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n568), .A2(new_n570), .A3(KEYINPUT17), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT92), .B1(new_n549), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n544), .A2(new_n546), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT91), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n544), .A2(new_n546), .A3(new_n545), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n572), .B1(new_n568), .B2(new_n570), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n568), .A2(new_n570), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(KEYINPUT17), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT92), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT93), .Z(new_n588));
  INV_X1    g387(.A(new_n578), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n571), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n577), .A2(new_n586), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT18), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n588), .A2(KEYINPUT18), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n577), .A2(new_n586), .A3(new_n590), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n583), .A2(new_n578), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n588), .B(KEYINPUT94), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT13), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n535), .B1(new_n593), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT95), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n591), .A2(new_n592), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n604), .A2(new_n600), .A3(new_n534), .A4(new_n595), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(KEYINPUT95), .B(new_n535), .C1(new_n593), .C2(new_n601), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n528), .A2(KEYINPUT96), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n487), .A2(new_n527), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(new_n608), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT101), .B(G183gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G211gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n620));
  XOR2_X1   g419(.A(G57gat), .B(G64gat), .Z(new_n621));
  NAND2_X1  g420(.A1(G71gat), .A2(G78gat), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT9), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT98), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n622), .A2(new_n626), .A3(new_n623), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n621), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n622), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(KEYINPUT97), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n630), .B1(new_n628), .B2(new_n631), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n620), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n636), .A2(KEYINPUT99), .A3(new_n632), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT21), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G127gat), .B(G155gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT20), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n635), .A2(new_n637), .A3(new_n638), .A4(new_n640), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n645), .B1(new_n642), .B2(new_n646), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n619), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n649), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n647), .A3(new_n618), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n589), .B1(new_n653), .B2(KEYINPUT21), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n650), .B2(new_n652), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n616), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n650), .A2(new_n652), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n654), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n615), .A3(new_n656), .ZN(new_n662));
  XNOR2_X1  g461(.A(G134gat), .B(G162gat), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n664));
  INV_X1    g463(.A(G232gat), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n665), .B2(new_n258), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n663), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G190gat), .B(G218gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT102), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT103), .Z(new_n670));
  NAND2_X1  g469(.A1(G85gat), .A2(G92gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT7), .ZN(new_n672));
  NAND2_X1  g471(.A1(G99gat), .A2(G106gat), .ZN(new_n673));
  INV_X1    g472(.A(G85gat), .ZN(new_n674));
  AOI22_X1  g473(.A1(KEYINPUT8), .A2(new_n673), .B1(new_n674), .B2(new_n353), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(G99gat), .B(G106gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n574), .A3(new_n575), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n664), .A2(new_n665), .A3(new_n258), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n678), .B2(new_n571), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n670), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n667), .B1(new_n683), .B2(KEYINPUT104), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n684), .A2(KEYINPUT105), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n680), .A2(new_n670), .A3(new_n682), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(KEYINPUT105), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n685), .B2(new_n688), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n637), .A2(new_n635), .A3(new_n679), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT10), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(new_n677), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n677), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n696), .B(new_n697), .C1(new_n634), .C2(new_n633), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n692), .A2(new_n693), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n653), .A2(KEYINPUT10), .A3(new_n678), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(G230gat), .A2(G233gat), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n692), .A2(new_n698), .ZN(new_n704));
  INV_X1    g503(.A(new_n702), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(G120gat), .B(G148gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G176gat), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(G204gat), .Z(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n703), .A2(new_n706), .A3(new_n710), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(KEYINPUT107), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n707), .A2(new_n715), .A3(new_n711), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n659), .A2(new_n662), .A3(new_n691), .A4(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT108), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n614), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n483), .A2(new_n484), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(new_n537), .ZN(G1324gat));
  INV_X1    g526(.A(new_n724), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT16), .B(G8gat), .Z(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(new_n361), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n728), .A2(KEYINPUT42), .A3(new_n361), .A4(new_n729), .ZN(new_n733));
  INV_X1    g532(.A(new_n361), .ZN(new_n734));
  OAI21_X1  g533(.A(G8gat), .B1(new_n724), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(G1325gat));
  INV_X1    g535(.A(new_n431), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n724), .A2(G15gat), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n526), .B(KEYINPUT109), .ZN(new_n739));
  OAI21_X1  g538(.A(G15gat), .B1(new_n724), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(G1326gat));
  INV_X1    g540(.A(new_n275), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n724), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT43), .B(G22gat), .Z(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1327gat));
  NAND2_X1  g544(.A1(new_n659), .A2(new_n662), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n714), .A2(new_n716), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n747), .A2(new_n691), .A3(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n614), .A2(new_n551), .A3(new_n523), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT45), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n608), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n606), .A2(KEYINPUT110), .A3(new_n607), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n717), .B(KEYINPUT111), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n758), .A3(new_n746), .ZN(new_n759));
  INV_X1    g558(.A(new_n691), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n487), .B2(new_n527), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT44), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT112), .B(KEYINPUT44), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n760), .B(new_n763), .C1(new_n487), .C2(new_n527), .ZN(new_n764));
  AOI211_X1 g563(.A(new_n725), .B(new_n759), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G29gat), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n751), .B1(new_n767), .B2(new_n768), .ZN(G1328gat));
  NAND3_X1  g568(.A1(new_n749), .A2(new_n552), .A3(new_n361), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n610), .B2(new_n613), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT46), .ZN(new_n772));
  AOI211_X1 g571(.A(new_n734), .B(new_n759), .C1(new_n762), .C2(new_n764), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G36gat), .B1(new_n773), .B2(new_n774), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(G1329gat));
  AND2_X1   g576(.A1(new_n614), .A2(new_n749), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n737), .A2(G43gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI211_X1 g579(.A(new_n526), .B(new_n759), .C1(new_n762), .C2(new_n764), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n780), .B(KEYINPUT47), .C1(new_n560), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n762), .A2(new_n764), .ZN(new_n783));
  INV_X1    g582(.A(new_n739), .ZN(new_n784));
  INV_X1    g583(.A(new_n759), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n778), .A2(new_n779), .B1(new_n786), .B2(G43gat), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n788));
  OAI21_X1  g587(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(G1330gat));
  NAND4_X1  g588(.A1(new_n614), .A2(new_n561), .A3(new_n275), .A4(new_n749), .ZN(new_n790));
  AOI211_X1 g589(.A(new_n742), .B(new_n759), .C1(new_n762), .C2(new_n764), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n561), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT116), .B1(new_n791), .B2(new_n561), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(KEYINPUT48), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT48), .ZN(new_n795));
  OAI221_X1 g594(.A(new_n790), .B1(KEYINPUT116), .B2(new_n795), .C1(new_n561), .C2(new_n791), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n794), .A2(new_n796), .ZN(G1331gat));
  NAND3_X1  g596(.A1(new_n755), .A2(new_n747), .A3(new_n691), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n612), .A2(new_n758), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n523), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT117), .B(G57gat), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1332gat));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n361), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n804));
  XOR2_X1   g603(.A(KEYINPUT49), .B(G64gat), .Z(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n803), .B2(new_n805), .ZN(G1333gat));
  NAND2_X1  g605(.A1(new_n799), .A2(new_n784), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n737), .A2(G71gat), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n807), .A2(G71gat), .B1(new_n799), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g609(.A1(new_n799), .A2(new_n275), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g611(.A1(new_n756), .A2(new_n747), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n760), .C1(new_n487), .C2(new_n527), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n814), .A2(new_n815), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(new_n717), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n674), .A3(new_n523), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n813), .A2(new_n748), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n762), .B2(new_n764), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G85gat), .B1(new_n824), .B2(new_n725), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(G1336gat));
  NAND3_X1  g625(.A1(new_n757), .A2(new_n353), .A3(new_n361), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT118), .Z(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n817), .B2(new_n818), .ZN(new_n829));
  AOI211_X1 g628(.A(new_n734), .B(new_n822), .C1(new_n762), .C2(new_n764), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n353), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n831), .A2(KEYINPUT119), .A3(KEYINPUT52), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT119), .B1(new_n831), .B2(KEYINPUT52), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n830), .A2(new_n353), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n819), .B2(new_n827), .ZN(new_n836));
  OAI22_X1  g635(.A1(new_n832), .A2(new_n833), .B1(new_n834), .B2(new_n836), .ZN(G1337gat));
  INV_X1    g636(.A(G99gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n820), .A2(new_n838), .A3(new_n431), .ZN(new_n839));
  OAI21_X1  g638(.A(G99gat), .B1(new_n824), .B2(new_n739), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1338gat));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843));
  INV_X1    g642(.A(new_n822), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n783), .A2(new_n275), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G106gat), .ZN(new_n846));
  INV_X1    g645(.A(G106gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n757), .A2(new_n847), .A3(new_n275), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n528), .A2(KEYINPUT51), .A3(new_n760), .A4(new_n813), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n816), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n843), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n847), .B1(new_n823), .B2(new_n275), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(KEYINPUT120), .A3(new_n850), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n842), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n846), .A2(new_n843), .A3(new_n851), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT120), .B1(new_n853), .B2(new_n850), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n855), .A2(new_n858), .ZN(G1339gat));
  NAND3_X1  g658(.A1(new_n699), .A2(new_n705), .A3(new_n700), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n703), .A2(new_n860), .A3(KEYINPUT54), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n705), .B1(new_n699), .B2(new_n700), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n710), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT55), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n713), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n861), .A2(KEYINPUT55), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n753), .A2(new_n754), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n577), .A2(new_n590), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n588), .B1(new_n872), .B2(new_n586), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n597), .A2(new_n599), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n533), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n714), .A2(new_n716), .A3(new_n605), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n760), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n605), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n869), .A2(new_n691), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n746), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n719), .A2(new_n755), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n275), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n725), .A2(new_n361), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n431), .A3(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n369), .A3(new_n608), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n476), .A2(new_n479), .A3(new_n734), .ZN(new_n886));
  AOI211_X1 g685(.A(new_n725), .B(new_n886), .C1(new_n880), .C2(new_n881), .ZN(new_n887));
  AOI21_X1  g686(.A(G113gat), .B1(new_n887), .B2(new_n756), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n885), .A2(new_n888), .ZN(G1340gat));
  OAI21_X1  g688(.A(G120gat), .B1(new_n884), .B2(new_n758), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n887), .A2(new_n382), .A3(new_n383), .A4(new_n748), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1341gat));
  OAI21_X1  g691(.A(G127gat), .B1(new_n884), .B2(new_n746), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n887), .A2(new_n363), .A3(new_n747), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT121), .ZN(G1342gat));
  NAND3_X1  g695(.A1(new_n887), .A2(new_n365), .A3(new_n760), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT56), .ZN(new_n898));
  OAI21_X1  g697(.A(G134gat), .B1(new_n884), .B2(new_n691), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(KEYINPUT56), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G1343gat));
  NAND4_X1  g700(.A1(new_n606), .A2(new_n867), .A3(new_n607), .A4(new_n868), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n760), .B1(new_n902), .B2(new_n876), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n746), .B1(new_n903), .B2(new_n879), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n742), .B1(new_n904), .B2(new_n881), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT57), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n526), .B(new_n883), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n742), .B1(new_n880), .B2(new_n881), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n210), .B1(new_n909), .B2(new_n756), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n725), .B1(new_n880), .B2(new_n881), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n739), .A2(new_n275), .A3(new_n734), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n608), .A2(G141gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  INV_X1    g717(.A(new_n916), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n210), .B1(new_n909), .B2(new_n609), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n917), .A2(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1344gat));
  NAND3_X1  g721(.A1(new_n915), .A2(new_n208), .A3(new_n748), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G148gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n925), .B1(new_n909), .B2(new_n748), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n609), .B1(new_n720), .B2(new_n722), .ZN(new_n927));
  INV_X1    g726(.A(new_n904), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n906), .B(new_n275), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n526), .A2(new_n748), .A3(new_n883), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n929), .B(new_n930), .C1(new_n908), .C2(new_n906), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n924), .B1(new_n931), .B2(G148gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n923), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g734(.A(KEYINPUT122), .B(new_n923), .C1(new_n926), .C2(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1345gat));
  INV_X1    g736(.A(new_n909), .ZN(new_n938));
  OAI21_X1  g737(.A(G155gat), .B1(new_n938), .B2(new_n746), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n915), .A2(new_n219), .A3(new_n747), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1346gat));
  OAI21_X1  g740(.A(G162gat), .B1(new_n938), .B2(new_n691), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n915), .A2(new_n220), .A3(new_n760), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1347gat));
  NAND2_X1  g743(.A1(new_n725), .A2(new_n361), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(KEYINPUT123), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(KEYINPUT123), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n431), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n882), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n952), .A2(new_n531), .A3(new_n608), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n523), .B1(new_n880), .B2(new_n881), .ZN(new_n954));
  AND4_X1   g753(.A1(new_n361), .A2(new_n954), .A3(new_n476), .A4(new_n479), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n756), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n953), .B1(new_n956), .B2(new_n531), .ZN(G1348gat));
  INV_X1    g756(.A(G176gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n958), .A3(new_n748), .ZN(new_n959));
  OAI21_X1  g758(.A(G176gat), .B1(new_n952), .B2(new_n758), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1349gat));
  NAND3_X1  g760(.A1(new_n955), .A2(new_n284), .A3(new_n747), .ZN(new_n962));
  OAI21_X1  g761(.A(G183gat), .B1(new_n952), .B2(new_n746), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT60), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT60), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n962), .A2(new_n966), .A3(new_n963), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1350gat));
  INV_X1    g767(.A(G190gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n955), .A2(new_n969), .A3(new_n760), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n951), .A2(new_n882), .A3(new_n760), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G190gat), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT125), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n971), .A2(new_n975), .A3(G190gat), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n974), .B1(new_n973), .B2(new_n976), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n970), .B1(new_n977), .B2(new_n978), .ZN(G1351gat));
  AND2_X1   g778(.A1(new_n739), .A2(new_n948), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n929), .B(new_n980), .C1(new_n908), .C2(new_n906), .ZN(new_n981));
  INV_X1    g780(.A(G197gat), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n981), .A2(new_n982), .A3(new_n608), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n954), .A2(new_n275), .A3(new_n361), .A4(new_n739), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n986), .A2(new_n756), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n983), .B1(new_n988), .B2(new_n982), .ZN(G1352gat));
  NOR3_X1   g788(.A1(new_n984), .A2(G204gat), .A3(new_n717), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(G204gat), .B1(new_n981), .B2(new_n758), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(G1353gat));
  OAI21_X1  g794(.A(G211gat), .B1(new_n981), .B2(new_n746), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT63), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND4_X1  g797(.A1(new_n986), .A2(new_n230), .A3(new_n747), .A4(new_n987), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1354gat));
  NOR3_X1   g799(.A1(new_n981), .A2(new_n231), .A3(new_n691), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n760), .A3(new_n987), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n1001), .B1(new_n1002), .B2(new_n231), .ZN(G1355gat));
endmodule


