//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n579, new_n580, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1228, new_n1229, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n461), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n461), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  OAI22_X1  g053(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(G136), .B2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT67), .Z(G162));
  OAI211_X1 g057(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT68), .B1(new_n461), .B2(G114), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT69), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n486), .A2(new_n489), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n492), .B(new_n483), .C1(new_n493), .C2(new_n485), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n461), .A2(G138), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n472), .B2(new_n473), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT71), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT4), .B1(new_n497), .B2(KEYINPUT70), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n461), .A2(G138), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(KEYINPUT70), .C1(new_n463), .C2(new_n462), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n499), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n501), .B1(new_n463), .B2(new_n462), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n507), .A2(KEYINPUT71), .A3(KEYINPUT4), .A4(new_n502), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n495), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT73), .B1(new_n514), .B2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(KEYINPUT72), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n519), .B2(G651), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  AOI211_X1 g096(.A(KEYINPUT73), .B(new_n521), .C1(new_n516), .C2(new_n518), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n513), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n515), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT72), .B(KEYINPUT6), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n527), .B2(new_n521), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n519), .A2(new_n529), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(KEYINPUT74), .A3(new_n513), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n525), .A2(G88), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  INV_X1    g109(.A(G62), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n511), .B2(new_n512), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(KEYINPUT75), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(KEYINPUT75), .ZN(new_n538));
  NAND2_X1  g113(.A1(G75), .A2(G543), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n528), .B2(new_n530), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n540), .A2(G651), .B1(new_n542), .B2(G50), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n533), .A2(new_n534), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n534), .B1(new_n533), .B2(new_n543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(G303));
  INV_X1    g121(.A(G303), .ZN(G166));
  AOI21_X1  g122(.A(KEYINPUT74), .B1(new_n531), .B2(new_n513), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n511), .A2(new_n512), .ZN(new_n549));
  AOI211_X1 g124(.A(new_n524), .B(new_n549), .C1(new_n528), .C2(new_n530), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G89), .ZN(new_n552));
  NAND3_X1  g127(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT7), .Z(new_n554));
  AND3_X1   g129(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n555));
  AOI211_X1 g130(.A(new_n554), .B(new_n555), .C1(new_n542), .C2(G51), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G286));
  INV_X1    g132(.A(G286), .ZN(G168));
  NAND2_X1  g133(.A1(G77), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G64), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n549), .B2(new_n560), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(KEYINPUT77), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n521), .B1(new_n561), .B2(KEYINPUT77), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n562), .A2(new_n563), .B1(G52), .B2(new_n542), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n525), .A2(new_n532), .ZN(new_n565));
  INV_X1    g140(.A(G90), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(G301));
  INV_X1    g142(.A(G301), .ZN(G171));
  NAND2_X1  g143(.A1(new_n551), .A2(G81), .ZN(new_n569));
  NAND2_X1  g144(.A1(G68), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G56), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n549), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n542), .A2(G43), .B1(G651), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  NAND4_X1  g151(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT78), .ZN(G176));
  NAND2_X1  g153(.A1(G1), .A2(G3), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT8), .ZN(new_n580));
  NAND4_X1  g155(.A1(G319), .A2(G483), .A3(G661), .A4(new_n580), .ZN(G188));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  AND2_X1   g157(.A1(KEYINPUT79), .A2(G53), .ZN(new_n583));
  AND3_X1   g158(.A1(new_n542), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n582), .B1(new_n542), .B2(new_n583), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n584), .A2(new_n585), .B1(new_n521), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n525), .A2(G91), .A3(new_n532), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G299));
  OAI21_X1  g165(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n592));
  AND2_X1   g167(.A1(G49), .A2(G543), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n531), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n592), .B1(new_n531), .B2(new_n593), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n551), .B2(G87), .ZN(new_n600));
  INV_X1    g175(.A(G87), .ZN(new_n601));
  NOR4_X1   g176(.A1(new_n548), .A2(new_n550), .A3(KEYINPUT80), .A4(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n598), .B1(new_n600), .B2(new_n602), .ZN(G288));
  AOI22_X1  g178(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n604), .A2(new_n605), .A3(new_n521), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n604), .B2(new_n521), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n606), .A2(new_n607), .B1(new_n542), .B2(G48), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n525), .A2(G86), .A3(new_n532), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(G305));
  NAND2_X1  g185(.A1(new_n551), .A2(G85), .ZN(new_n611));
  NAND2_X1  g186(.A1(G72), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G60), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n549), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n542), .A2(G47), .B1(G651), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(G301), .A2(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n542), .A2(G54), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n521), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n621));
  INV_X1    g196(.A(G92), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n565), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n551), .A2(KEYINPUT10), .A3(G92), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n617), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n617), .B1(new_n625), .B2(G868), .ZN(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n589), .B2(G868), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(new_n589), .B2(G868), .ZN(G280));
  NAND2_X1  g205(.A1(new_n623), .A2(new_n624), .ZN(new_n631));
  INV_X1    g206(.A(new_n620), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G860), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(G559), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT83), .ZN(G148));
  INV_X1    g211(.A(G868), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n574), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n633), .A2(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n638), .B1(new_n639), .B2(new_n637), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n480), .A2(G135), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n461), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  INV_X1    g219(.A(G123), .ZN(new_n645));
  OAI221_X1 g220(.A(new_n642), .B1(new_n643), .B2(new_n644), .C1(new_n645), .C2(new_n475), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT85), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2096), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n474), .A2(new_n468), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT13), .B(G2100), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n648), .A2(new_n653), .ZN(G156));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n668), .A3(G14), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT86), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2084), .B(G2090), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT87), .ZN(new_n674));
  XOR2_X1   g249(.A(G2067), .B(G2678), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(KEYINPUT17), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n672), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n672), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n679), .B2(new_n680), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT88), .B(G2096), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT89), .ZN(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(new_n693), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n696), .A2(new_n689), .A3(new_n697), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n695), .B(new_n698), .C1(new_n689), .C2(new_n696), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT90), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1991), .B(G1996), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n702), .A2(new_n703), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n708), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n707), .A2(new_n710), .ZN(G229));
  NAND2_X1  g286(.A1(G168), .A2(G16), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(KEYINPUT96), .C1(G16), .C2(G21), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(KEYINPUT96), .B2(new_n712), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(G1966), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G32), .ZN(new_n717));
  INV_X1    g292(.A(new_n475), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G129), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n468), .A2(G105), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n480), .A2(G141), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND4_X1  g298(.A1(new_n719), .A2(new_n720), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n717), .B1(new_n725), .B2(new_n716), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT27), .ZN(new_n727));
  INV_X1    g302(.A(G1996), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n716), .A2(G26), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n480), .A2(G140), .ZN(new_n732));
  OR2_X1    g307(.A1(G104), .A2(G2105), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n733), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n734));
  INV_X1    g309(.A(G128), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n734), .C1(new_n475), .C2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n731), .B1(new_n738), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G2067), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n716), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n716), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2078), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n715), .A2(new_n729), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n714), .A2(G1966), .ZN(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G35), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G162), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT29), .ZN(new_n749));
  INV_X1    g324(.A(G2090), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AND3_X1   g326(.A1(new_n745), .A2(new_n746), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n480), .A2(G139), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n754), .B(new_n755), .C1(new_n461), .C2(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT95), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G29), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G33), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT94), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2072), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n647), .A2(G29), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT97), .Z(new_n765));
  XOR2_X1   g340(.A(KEYINPUT31), .B(G11), .Z(new_n766));
  INV_X1    g341(.A(G28), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(KEYINPUT30), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT98), .ZN(new_n769));
  AOI21_X1  g344(.A(G29), .B1(new_n767), .B2(KEYINPUT30), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n772), .B2(KEYINPUT24), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(KEYINPUT24), .B2(new_n772), .ZN(new_n774));
  INV_X1    g349(.A(G160), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n716), .ZN(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n771), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n777), .B2(new_n776), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n763), .A2(new_n765), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G1961), .ZN(new_n781));
  INV_X1    g356(.A(G16), .ZN(new_n782));
  NOR2_X1   g357(.A1(G171), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G5), .B2(new_n782), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n780), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(G20), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT23), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n589), .B2(new_n782), .ZN(new_n788));
  INV_X1    g363(.A(G1956), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G16), .A2(G19), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n575), .B2(G16), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1341), .Z(new_n793));
  AND3_X1   g368(.A1(new_n785), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n784), .A2(new_n781), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT99), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n782), .A2(G4), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n625), .B2(new_n782), .ZN(new_n798));
  INV_X1    g373(.A(G1348), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n752), .A2(new_n794), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT36), .ZN(new_n802));
  INV_X1    g377(.A(G290), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(new_n782), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n782), .B2(G24), .ZN(new_n805));
  INV_X1    g380(.A(G1986), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n716), .A2(G25), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n718), .A2(G119), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n480), .A2(G131), .ZN(new_n811));
  OR2_X1    g386(.A1(G95), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n809), .B1(new_n815), .B2(new_n716), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n807), .A2(new_n808), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n782), .A2(G23), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT80), .B1(new_n565), .B2(new_n601), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n551), .A2(new_n599), .A3(G87), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n597), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n820), .B1(new_n823), .B2(new_n782), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT33), .B(G1976), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n824), .B(new_n825), .Z(new_n826));
  AND2_X1   g401(.A1(new_n608), .A2(new_n609), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G16), .ZN(new_n828));
  OR2_X1    g403(.A1(G6), .A2(G16), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT32), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT32), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n828), .A2(new_n832), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G1981), .ZN(new_n835));
  INV_X1    g410(.A(G1981), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n831), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n826), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(G303), .A2(G16), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n782), .A2(G22), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT91), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G1971), .ZN(new_n843));
  INV_X1    g418(.A(G1971), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n839), .A2(new_n844), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n843), .A2(KEYINPUT92), .A3(new_n845), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n838), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n819), .B1(new_n850), .B2(KEYINPUT34), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT34), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n838), .A2(new_n852), .A3(new_n848), .A4(new_n849), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n802), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n851), .A2(new_n802), .A3(new_n853), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n801), .B1(new_n855), .B2(new_n856), .ZN(G311));
  INV_X1    g432(.A(new_n801), .ZN(new_n858));
  INV_X1    g433(.A(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n859), .B2(new_n854), .ZN(G150));
  NAND2_X1  g435(.A1(new_n625), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n551), .A2(G93), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT100), .B(G55), .Z(new_n864));
  NAND2_X1  g439(.A1(G80), .A2(G543), .ZN(new_n865));
  INV_X1    g440(.A(G67), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n549), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n542), .A2(new_n864), .B1(G651), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n569), .A2(new_n863), .A3(new_n573), .A4(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n569), .A2(new_n573), .B1(new_n863), .B2(new_n868), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n862), .B(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n634), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G93), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n868), .B1(new_n565), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G860), .ZN(new_n879));
  XOR2_X1   g454(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n881), .ZN(G145));
  XNOR2_X1  g457(.A(new_n647), .B(G160), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G162), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n484), .A2(new_n490), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n738), .A2(new_n504), .A3(new_n508), .A4(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n736), .B(KEYINPUT93), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n504), .A2(new_n508), .A3(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n886), .A2(new_n725), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n725), .B1(new_n886), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n758), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g469(.A(KEYINPUT102), .B(new_n758), .C1(new_n890), .C2(new_n891), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n890), .A2(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n757), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n651), .ZN(new_n899));
  INV_X1    g474(.A(G130), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n461), .A2(G118), .ZN(new_n901));
  OAI21_X1  g476(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n475), .A2(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(G142), .B2(new_n480), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n815), .B(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT103), .ZN(new_n906));
  INV_X1    g481(.A(new_n651), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n894), .A2(new_n897), .A3(new_n907), .A4(new_n895), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n899), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n899), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n884), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n899), .A2(new_n908), .ZN(new_n912));
  INV_X1    g487(.A(new_n906), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n884), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n899), .A2(new_n906), .A3(new_n908), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n911), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g495(.A1(new_n878), .A2(new_n637), .ZN(new_n921));
  NAND2_X1  g496(.A1(G288), .A2(KEYINPUT105), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n823), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n803), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n924), .A3(G290), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(G305), .B1(new_n544), .B2(new_n545), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n533), .A2(new_n543), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT76), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n533), .A2(new_n534), .A3(new_n543), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n827), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n929), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n929), .B2(new_n933), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n928), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n926), .A2(new_n935), .A3(new_n927), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT42), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n872), .B(new_n639), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n625), .A2(new_n589), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n625), .A2(new_n589), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n942), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n945), .B2(new_n943), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n633), .A2(G299), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n944), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n946), .B1(new_n953), .B2(new_n942), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n941), .B(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n921), .B1(new_n955), .B2(new_n637), .ZN(G295));
  OAI21_X1  g531(.A(new_n921), .B1(new_n955), .B2(new_n637), .ZN(G331));
  AOI21_X1  g532(.A(G286), .B1(G171), .B2(KEYINPUT107), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n574), .A2(new_n878), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n961));
  NAND2_X1  g536(.A1(G301), .A2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n960), .A2(new_n869), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n960), .B2(new_n869), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n962), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n870), .B2(new_n871), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(new_n869), .A3(new_n962), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n958), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n953), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n945), .A2(new_n943), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n965), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n971), .A2(new_n938), .A3(new_n939), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n918), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n971), .A2(new_n973), .B1(new_n938), .B2(new_n939), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT43), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n978));
  INV_X1    g553(.A(new_n970), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n950), .A2(new_n944), .A3(new_n948), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n972), .B2(KEYINPUT41), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n973), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n940), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n918), .A4(new_n974), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n977), .A2(new_n978), .A3(new_n985), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n969), .A2(new_n965), .B1(new_n949), .B2(new_n952), .ZN(new_n987));
  INV_X1    g562(.A(new_n973), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n940), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n989), .A2(new_n984), .A3(new_n918), .A4(new_n974), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n988), .A2(new_n987), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n938), .A2(new_n939), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n995), .A2(KEYINPUT108), .A3(new_n984), .A4(new_n989), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n982), .A2(new_n940), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n997), .B2(new_n975), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n992), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n986), .B1(KEYINPUT44), .B2(new_n999), .ZN(G397));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n1001));
  NAND4_X1  g576(.A1(G303), .A2(new_n1001), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT113), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n931), .A2(G8), .A3(new_n932), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1002), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n888), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n467), .A2(new_n469), .ZN(new_n1013));
  INV_X1    g588(.A(G125), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n472), .B2(new_n473), .ZN(new_n1015));
  INV_X1    g590(.A(new_n465), .ZN(new_n1016));
  OAI21_X1  g591(.A(G2105), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1017), .A3(G40), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1011), .A2(new_n1012), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n888), .B2(new_n1009), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT115), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n509), .A2(new_n1024), .A3(new_n1009), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1023), .A2(new_n1027), .A3(new_n750), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n509), .A2(new_n1009), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n888), .A2(KEYINPUT45), .A3(new_n1009), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1022), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n844), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1029), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1008), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n888), .A2(new_n1024), .A3(new_n1009), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1022), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1024), .B1(new_n509), .B2(new_n1009), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1010), .A2(new_n1031), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n1009), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n1022), .ZN(new_n1045));
  INV_X1    g620(.A(G1966), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n777), .A2(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1047), .A2(new_n1048), .A3(G286), .ZN(new_n1049));
  INV_X1    g624(.A(G1976), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G288), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1010), .A2(new_n1026), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n1048), .ZN(new_n1054));
  OAI211_X1 g629(.A(G1976), .B(new_n598), .C1(new_n600), .C2(new_n602), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1054), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT52), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n836), .B1(new_n608), .B2(new_n609), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n608), .A2(new_n609), .A3(new_n836), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(KEYINPUT49), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT49), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1061), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(new_n1059), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1065), .A3(new_n1054), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1056), .A2(new_n1058), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1002), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1040), .A2(G2090), .A3(new_n1041), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1048), .B1(new_n1070), .B2(new_n1035), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1038), .A2(new_n1049), .A3(new_n1067), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT116), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1077), .A3(new_n1074), .ZN(new_n1078));
  NOR4_X1   g653(.A1(new_n1047), .A2(new_n1074), .A3(new_n1048), .A4(G286), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT45), .B1(new_n509), .B2(new_n1009), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(new_n1026), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1971), .B1(new_n1081), .B2(new_n1033), .ZN(new_n1082));
  OAI21_X1  g657(.A(G8), .B1(new_n1082), .B2(new_n1069), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(new_n1004), .A3(new_n1007), .A4(new_n1002), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1067), .A2(new_n1072), .A3(new_n1079), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT117), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1041), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1087), .A2(new_n777), .A3(new_n1022), .A4(new_n1039), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1043), .A2(new_n1044), .A3(new_n1022), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(G1966), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1090), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1008), .B2(new_n1083), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1072), .A4(new_n1067), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1076), .A2(new_n1078), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1026), .B1(new_n1010), .B2(new_n1031), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1966), .B1(new_n1097), .B2(new_n1044), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1040), .A2(G2084), .A3(new_n1041), .ZN(new_n1099));
  OAI211_X1 g674(.A(G8), .B(G286), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT120), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1090), .A2(new_n1102), .A3(G8), .A4(G286), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1088), .B(G168), .C1(new_n1089), .C2(G1966), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(KEYINPUT51), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1105), .A2(G8), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1048), .B1(new_n1047), .B2(G168), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT121), .B(KEYINPUT51), .Z(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1104), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1038), .A2(new_n1072), .A3(new_n1067), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1023), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1033), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1116), .A2(new_n1080), .A3(new_n1026), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT56), .B(G2072), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1115), .A2(new_n789), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n589), .B(KEYINPUT57), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n799), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1053), .A2(new_n740), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(new_n633), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1121), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT58), .B(G1341), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1034), .A2(G1996), .B1(new_n1053), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n575), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT59), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1132), .A3(new_n575), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1123), .A2(KEYINPUT60), .A3(new_n1124), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1123), .A2(KEYINPUT119), .A3(KEYINPUT60), .A4(new_n1124), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1137), .A2(new_n625), .A3(new_n1138), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1137), .A2(new_n625), .B1(KEYINPUT60), .B2(new_n1125), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1134), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1115), .A2(new_n789), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(KEYINPUT118), .ZN(new_n1145));
  AND4_X1   g720(.A1(new_n1120), .A2(new_n1142), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1127), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(G2078), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1150), .A2(KEYINPUT53), .ZN(new_n1151));
  AND3_X1   g726(.A1(G160), .A2(G40), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1043), .A2(new_n1033), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT123), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n781), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1043), .A2(new_n1156), .A3(new_n1033), .A4(new_n1152), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1160), .B1(new_n1117), .B2(new_n1150), .ZN(new_n1161));
  OAI21_X1  g736(.A(G171), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1162), .A2(KEYINPUT125), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(KEYINPUT125), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1097), .A2(new_n1044), .A3(new_n1151), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1155), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1159), .B1(new_n1034), .B2(G2078), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(G301), .A3(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1163), .A2(KEYINPUT54), .A3(new_n1164), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1158), .A2(new_n1161), .A3(G171), .ZN(new_n1171));
  AOI21_X1  g746(.A(G301), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(KEYINPUT124), .B(new_n1170), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1114), .A2(new_n1149), .A3(new_n1169), .A4(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1038), .A2(new_n1072), .A3(new_n1067), .A4(new_n1172), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1179), .B1(new_n1112), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(KEYINPUT62), .B1(new_n1104), .B2(new_n1111), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g759(.A(KEYINPUT126), .B(KEYINPUT62), .C1(new_n1104), .C2(new_n1111), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1181), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1066), .A2(new_n1050), .A3(new_n823), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1054), .B1(new_n1187), .B2(new_n1064), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1067), .A2(new_n1071), .A3(new_n1068), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1188), .A2(new_n1189), .A3(KEYINPUT114), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT114), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1096), .A2(new_n1178), .A3(new_n1186), .A4(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1022), .A2(new_n1010), .A3(new_n1031), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT110), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n887), .A2(new_n740), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n738), .A2(G2067), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1199), .A2(KEYINPUT111), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(KEYINPUT111), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n724), .B(G1996), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1195), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n814), .B(new_n817), .ZN(new_n1205));
  XOR2_X1   g780(.A(new_n1205), .B(KEYINPUT112), .Z(new_n1206));
  AND2_X1   g781(.A1(new_n1195), .A2(new_n1206), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(G290), .B(G1986), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1208), .B1(new_n1195), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1193), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1195), .A2(new_n806), .A3(new_n803), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT48), .Z(new_n1213));
  NAND2_X1  g788(.A1(new_n1195), .A2(new_n728), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT46), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1196), .A2(new_n1197), .A3(new_n725), .ZN(new_n1216));
  AOI22_X1  g791(.A1(new_n1214), .A2(new_n1215), .B1(new_n1195), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1217), .B1(new_n1215), .B2(new_n1214), .ZN(new_n1218));
  AND2_X1   g793(.A1(new_n1218), .A2(KEYINPUT47), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1218), .A2(KEYINPUT47), .ZN(new_n1220));
  OAI22_X1  g795(.A1(new_n1208), .A2(new_n1213), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n815), .A2(new_n817), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1196), .B1(new_n1204), .B2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1223), .B(KEYINPUT127), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1221), .B1(new_n1224), .B2(new_n1195), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1211), .A2(new_n1225), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g801(.A1(new_n686), .A2(G319), .A3(new_n670), .ZN(new_n1228));
  AOI21_X1  g802(.A(new_n1228), .B1(new_n707), .B2(new_n710), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n977), .A2(new_n985), .ZN(new_n1230));
  NAND3_X1  g804(.A1(new_n1229), .A2(new_n919), .A3(new_n1230), .ZN(G225));
  INV_X1    g805(.A(G225), .ZN(G308));
endmodule


