//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1184, new_n1185, new_n1186, new_n1187, new_n1189,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1240, new_n1241, new_n1242, new_n1243;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n209), .B(new_n215), .C1(G58), .C2(G232), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G1), .B2(G20), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT1), .Z(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G1), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n224), .A2(new_n221), .A3(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NOR3_X1   g0027(.A1(new_n218), .A2(new_n223), .A3(new_n227), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  INV_X1    g0031(.A(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n208), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G107), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n207), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G58), .ZN(new_n244));
  INV_X1    g0044(.A(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n242), .B(new_n246), .Z(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n222), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n252), .A2(new_n254), .B1(G150), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n203), .A2(G20), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n250), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n224), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n258), .A2(KEYINPUT68), .B1(new_n202), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n224), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n250), .A2(new_n262), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n261), .B1(KEYINPUT68), .B2(new_n258), .C1(new_n202), .C2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1698), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n268), .A2(G222), .B1(G77), .B2(new_n267), .ZN(new_n269));
  INV_X1    g0069(.A(G223), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n269), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n222), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT66), .B1(new_n276), .B2(new_n222), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT66), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n275), .A2(new_n280), .A3(G1), .A4(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n224), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G226), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n279), .B2(new_n281), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n285), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n278), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT67), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n264), .B1(new_n293), .B2(G169), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n291), .A2(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n292), .ZN(new_n296));
  AOI21_X1  g0096(.A(G179), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(G190), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n264), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n295), .A2(G200), .A3(new_n296), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n264), .A2(new_n300), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n299), .A2(new_n301), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n302), .A2(new_n303), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(new_n301), .A4(new_n299), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n298), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT72), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  OAI211_X1 g0111(.A(G226), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n312));
  OAI211_X1 g0112(.A(G223), .B(new_n271), .C1(new_n265), .C2(new_n266), .ZN(new_n313));
  INV_X1    g0113(.A(G87), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n312), .B(new_n313), .C1(new_n253), .C2(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n277), .B1(new_n289), .B2(new_n285), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n282), .A2(G232), .A3(new_n284), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n311), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n277), .ZN(new_n319));
  AND4_X1   g0119(.A1(G179), .A2(new_n319), .A3(new_n290), .A4(new_n317), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n310), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(G179), .A3(new_n317), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n319), .A2(new_n290), .A3(new_n317), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n322), .B(KEYINPUT72), .C1(new_n323), .C2(new_n311), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT7), .B1(new_n267), .B2(new_n221), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  NOR4_X1   g0127(.A1(new_n265), .A2(new_n266), .A3(new_n327), .A4(G20), .ZN(new_n328));
  OAI21_X1  g0128(.A(G68), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n255), .A2(G159), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G58), .A2(G68), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(G20), .B1(new_n332), .B2(new_n201), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n329), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n330), .A4(new_n333), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n249), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n252), .A2(new_n262), .A3(new_n250), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n251), .A2(new_n260), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT18), .B1(new_n325), .B2(new_n341), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n325), .A2(KEYINPUT18), .A3(new_n341), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT73), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n325), .A2(KEYINPUT18), .A3(new_n341), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT73), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n323), .A2(G190), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n338), .A2(new_n348), .A3(new_n339), .A4(new_n340), .ZN(new_n349));
  INV_X1    g0149(.A(G200), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n323), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT17), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OR3_X1    g0152(.A1(new_n349), .A2(KEYINPUT17), .A3(new_n351), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n345), .A2(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OR2_X1    g0154(.A1(KEYINPUT3), .A2(G33), .ZN(new_n355));
  NAND2_X1  g0155(.A1(KEYINPUT3), .A2(G33), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(G232), .A3(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n271), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n358), .B(new_n359), .C1(new_n360), .C2(new_n232), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n277), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT69), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n286), .A2(G238), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(KEYINPUT69), .A3(new_n277), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .A4(new_n290), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n367), .A2(KEYINPUT13), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(KEYINPUT13), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n260), .A2(KEYINPUT12), .A3(new_n211), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT12), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n259), .B2(G68), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n373), .B(new_n375), .C1(new_n263), .C2(new_n211), .ZN(new_n376));
  XOR2_X1   g0176(.A(new_n376), .B(KEYINPUT71), .Z(new_n377));
  AOI22_X1  g0177(.A1(new_n254), .A2(G77), .B1(new_n255), .B2(G50), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n211), .A2(G20), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n250), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g0180(.A(KEYINPUT70), .B(KEYINPUT11), .Z(new_n381));
  XNOR2_X1  g0181(.A(new_n380), .B(new_n381), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n350), .B1(new_n368), .B2(new_n369), .ZN(new_n384));
  OR3_X1    g0184(.A1(new_n372), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n309), .A2(new_n354), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n370), .A2(G169), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT14), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n368), .A2(G179), .A3(new_n369), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT14), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n370), .A2(new_n390), .A3(G169), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n383), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n357), .A2(G232), .A3(new_n271), .ZN(new_n394));
  INV_X1    g0194(.A(G107), .ZN(new_n395));
  OAI221_X1 g0195(.A(new_n394), .B1(new_n395), .B2(new_n357), .C1(new_n273), .C2(new_n212), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n277), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n286), .A2(G244), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n290), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n311), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n252), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n401));
  INV_X1    g0201(.A(new_n254), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT15), .B(G87), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(new_n249), .B1(new_n245), .B2(new_n260), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n245), .B2(new_n263), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n400), .B(new_n406), .C1(G179), .C2(new_n399), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n406), .B1(new_n399), .B2(G200), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n371), .B2(new_n399), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n393), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n386), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT78), .B(G116), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n413), .A2(G20), .A3(new_n253), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT23), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n221), .B2(G107), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n395), .A2(KEYINPUT23), .A3(G20), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n221), .B(G87), .C1(new_n265), .C2(new_n266), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT22), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT82), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT82), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(new_n422), .A3(KEYINPUT22), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT85), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT84), .ZN(new_n426));
  XOR2_X1   g0226(.A(KEYINPUT83), .B(KEYINPUT22), .Z(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(new_n419), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(G20), .B1(new_n355), .B2(new_n356), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(KEYINPUT84), .A3(G87), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n424), .A2(new_n425), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n425), .B1(new_n424), .B2(new_n432), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n418), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT86), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(KEYINPUT86), .B(new_n418), .C1(new_n433), .C2(new_n434), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(KEYINPUT24), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT24), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n249), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n260), .A2(new_n395), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT25), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n250), .B(new_n259), .C1(G1), .C2(new_n253), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT75), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n445), .B(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n447), .B2(G107), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT87), .B1(new_n273), .B2(new_n214), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT87), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n272), .A2(new_n451), .A3(G257), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G294), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n268), .A2(G250), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n450), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT5), .B(G41), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n283), .A2(new_n459), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n455), .A2(new_n277), .B1(G264), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n289), .A2(new_n459), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n311), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(G179), .B2(new_n463), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n449), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT19), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n221), .B1(new_n359), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G97), .A2(G107), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n314), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n472), .A2(KEYINPUT79), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n429), .A2(G68), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(KEYINPUT79), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n468), .B1(new_n402), .B2(new_n213), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n473), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n477), .A2(new_n249), .B1(new_n260), .B2(new_n403), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n445), .B(KEYINPUT75), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n403), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n357), .A2(G244), .A3(G1698), .ZN(new_n481));
  OAI221_X1 g0281(.A(new_n481), .B1(new_n253), .B2(new_n413), .C1(new_n360), .C2(new_n212), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n277), .ZN(new_n483));
  INV_X1    g0283(.A(G250), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT77), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n458), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n282), .B(new_n486), .C1(new_n485), .C2(new_n458), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n458), .A2(KEYINPUT66), .A3(G274), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n483), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n311), .ZN(new_n490));
  INV_X1    g0290(.A(G179), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n483), .A2(new_n491), .A3(new_n487), .A4(new_n488), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n480), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT6), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n213), .A2(new_n395), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(new_n470), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n395), .A2(KEYINPUT6), .A3(G97), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(new_n221), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n327), .B1(new_n357), .B2(G20), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n395), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n245), .A2(G20), .A3(G33), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n499), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n250), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT74), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n259), .A2(G97), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n479), .A2(new_n213), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n268), .B(G244), .C1(KEYINPUT76), .C2(KEYINPUT4), .ZN(new_n510));
  NOR2_X1   g0310(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n511));
  INV_X1    g0311(.A(G244), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n360), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n272), .A2(G250), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n510), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n277), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n460), .A2(G257), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n462), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G200), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n507), .A2(new_n506), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n517), .A2(G190), .A3(new_n518), .A4(new_n462), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n509), .A2(new_n520), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n489), .A2(G200), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n447), .A2(G87), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n483), .A2(G190), .A3(new_n487), .A4(new_n488), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n524), .A2(new_n478), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n507), .A2(new_n506), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n447), .B2(G97), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n529), .B(new_n521), .C1(new_n504), .C2(new_n250), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n519), .A2(new_n311), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n517), .A2(new_n491), .A3(new_n518), .A4(new_n462), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND4_X1   g0333(.A1(new_n493), .A2(new_n523), .A3(new_n527), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n463), .A2(new_n350), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G190), .B2(new_n463), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n442), .A2(new_n448), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n445), .A2(new_n207), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n515), .B(new_n221), .C1(G33), .C2(new_n213), .ZN(new_n539));
  INV_X1    g0339(.A(new_n413), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n249), .B(new_n539), .C1(new_n540), .C2(new_n221), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT20), .ZN(new_n542));
  OR2_X1    g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n538), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n540), .A2(new_n259), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n272), .A2(G264), .ZN(new_n549));
  XNOR2_X1  g0349(.A(KEYINPUT80), .B(G303), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n267), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n549), .B(new_n551), .C1(new_n214), .C2(new_n360), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n277), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n460), .A2(G270), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n462), .A3(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n548), .A2(new_n555), .A3(KEYINPUT21), .A4(G169), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT81), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(new_n491), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n556), .A2(new_n557), .B1(new_n558), .B2(new_n548), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n311), .B1(new_n545), .B2(new_n547), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n555), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n555), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G190), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n555), .A2(G200), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n565), .A2(new_n547), .A3(new_n545), .A4(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n560), .A2(KEYINPUT81), .A3(KEYINPUT21), .A4(new_n555), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n559), .A2(new_n563), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n467), .A2(new_n534), .A3(new_n537), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n412), .A2(new_n571), .ZN(G372));
  NAND2_X1  g0372(.A1(new_n393), .A2(new_n407), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n372), .A2(new_n383), .A3(new_n384), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n352), .B2(new_n353), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n342), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n346), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n298), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n559), .A2(new_n563), .A3(new_n568), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n467), .A2(KEYINPUT88), .A3(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n537), .A2(new_n534), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT88), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n465), .B1(new_n442), .B2(new_n448), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n588), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n493), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n527), .A2(new_n493), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n533), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT26), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT26), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n597), .B2(new_n533), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n596), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n411), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n587), .A2(new_n605), .ZN(G369));
  INV_X1    g0406(.A(G13), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(G20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n224), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n609), .A2(KEYINPUT27), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(KEYINPUT27), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(G213), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(G343), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n442), .B2(new_n448), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT89), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n467), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n537), .B1(new_n616), .B2(new_n617), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n588), .A2(new_n615), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n467), .A2(new_n614), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT90), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n620), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n593), .B1(new_n617), .B2(new_n616), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(new_n588), .A3(new_n615), .A4(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT90), .ZN(new_n628));
  INV_X1    g0428(.A(new_n623), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n548), .A2(new_n614), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n570), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n589), .B2(new_n632), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G330), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n625), .A2(new_n626), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n593), .A2(new_n614), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n631), .A2(new_n639), .ZN(G399));
  NOR2_X1   g0440(.A1(new_n471), .A2(G116), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT91), .ZN(new_n642));
  INV_X1    g0442(.A(new_n225), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(G41), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n644), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n645), .A2(new_n224), .B1(new_n220), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT92), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT28), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n604), .A2(new_n615), .ZN(new_n650));
  XOR2_X1   g0450(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n651));
  AOI21_X1  g0451(.A(new_n588), .B1(new_n449), .B2(new_n466), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n537), .A2(new_n534), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n603), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(KEYINPUT29), .A3(new_n615), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT95), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n534), .B(new_n537), .C1(new_n593), .C2(new_n588), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n614), .B1(new_n657), .B2(new_n603), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT95), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT29), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n650), .A2(new_n651), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n517), .A2(new_n518), .A3(new_n462), .ZN(new_n663));
  INV_X1    g0463(.A(new_n489), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n558), .A2(new_n663), .A3(new_n664), .A4(new_n461), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT30), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n519), .A2(new_n489), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(KEYINPUT30), .A3(new_n461), .A4(new_n558), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n564), .A2(G179), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n463), .A3(new_n489), .A4(new_n519), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(KEYINPUT31), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n615), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n571), .B2(KEYINPUT31), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n614), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT93), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n676), .B(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(G330), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n662), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n649), .B1(new_n681), .B2(G1), .ZN(G364));
  INV_X1    g0482(.A(new_n635), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n224), .B1(new_n608), .B2(G45), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n644), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(G330), .B2(new_n634), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n643), .A2(new_n357), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n219), .A2(new_n457), .A3(G50), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n689), .B(new_n690), .C1(new_n246), .C2(new_n457), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n643), .A2(new_n267), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G355), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n691), .B(new_n693), .C1(G116), .C2(new_n225), .ZN(new_n694));
  NOR2_X1   g0494(.A1(G13), .A2(G33), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G20), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n222), .B1(G20), .B2(new_n311), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n686), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n491), .A2(G200), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT98), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n221), .A2(new_n371), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n706), .A2(G303), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n221), .A2(G190), .ZN(new_n708));
  NOR2_X1   g0508(.A1(G179), .A2(G200), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT101), .Z(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(G329), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n491), .A2(G200), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n704), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT96), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n715), .A2(KEYINPUT96), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n707), .B(new_n713), .C1(G322), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n708), .A2(new_n714), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G311), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n703), .A2(new_n708), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT99), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G283), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n221), .A2(new_n491), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G200), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G190), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G317), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(KEYINPUT33), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(KEYINPUT33), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n729), .A2(new_n371), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n357), .B1(new_n735), .B2(G326), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n221), .B1(new_n709), .B2(G190), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT100), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT100), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n737), .B1(G294), .B2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n721), .A2(new_n724), .A3(new_n727), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(G97), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n211), .B2(new_n731), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n267), .B(new_n746), .C1(G50), .C2(new_n735), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n726), .A2(G107), .ZN(new_n748));
  INV_X1    g0548(.A(G58), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n719), .A2(new_n749), .B1(new_n314), .B2(new_n705), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n723), .A2(KEYINPUT97), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n723), .A2(KEYINPUT97), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(G77), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n747), .A2(new_n748), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n710), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G159), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT32), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n744), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n701), .B1(new_n760), .B2(new_n698), .ZN(new_n761));
  INV_X1    g0561(.A(new_n697), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n700), .B(new_n761), .C1(new_n634), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n688), .A2(new_n763), .ZN(G396));
  NOR2_X1   g0564(.A1(new_n407), .A2(new_n614), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n406), .A2(new_n614), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n409), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(new_n767), .B2(new_n407), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n650), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n614), .B1(new_n595), .B2(new_n603), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n768), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n679), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n676), .B(KEYINPUT93), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT31), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n569), .B1(new_n449), .B2(new_n466), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(new_n591), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n775), .B1(new_n778), .B2(new_n674), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n770), .A2(G330), .A3(new_n779), .A4(new_n772), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n774), .A2(new_n701), .A3(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n754), .A2(G159), .B1(G137), .B2(new_n735), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n720), .A2(G143), .ZN(new_n783));
  INV_X1    g0583(.A(G150), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n731), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT34), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n357), .B1(new_n705), .B2(new_n202), .C1(new_n741), .C2(new_n749), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G68), .B2(new_n726), .ZN(new_n788));
  INV_X1    g0588(.A(G132), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n786), .B(new_n788), .C1(new_n789), .C2(new_n711), .ZN(new_n790));
  INV_X1    g0590(.A(G294), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n745), .B1(new_n791), .B2(new_n719), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT103), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n711), .A2(new_n794), .B1(new_n395), .B2(new_n705), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n267), .B1(new_n753), .B2(new_n413), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n730), .A2(KEYINPUT102), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n730), .A2(KEYINPUT102), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n795), .B(new_n796), .C1(G283), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n735), .A2(G303), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n726), .A2(G87), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n793), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n790), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n701), .B1(new_n805), .B2(new_n698), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n698), .A2(new_n695), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n245), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n806), .B(new_n808), .C1(new_n696), .C2(new_n768), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n781), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n810), .A2(KEYINPUT104), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(KEYINPUT104), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G384));
  AOI21_X1  g0614(.A(new_n586), .B1(new_n661), .B2(new_n411), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT106), .Z(new_n816));
  NAND2_X1  g0616(.A1(new_n383), .A2(new_n614), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n390), .B1(new_n370), .B2(G169), .ZN(new_n818));
  AOI211_X1 g0618(.A(KEYINPUT14), .B(new_n311), .C1(new_n368), .C2(new_n369), .ZN(new_n819));
  INV_X1    g0619(.A(new_n389), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n383), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n385), .B(new_n817), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n383), .B(new_n614), .C1(new_n392), .C2(new_n574), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n676), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n768), .B(new_n825), .C1(new_n675), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n612), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n341), .B1(new_n325), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n338), .A2(new_n339), .ZN(new_n830));
  INV_X1    g0630(.A(new_n351), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n830), .A2(new_n831), .A3(new_n348), .A4(new_n340), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT37), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n829), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n341), .A2(new_n828), .ZN(new_n838));
  OAI211_X1 g0638(.A(KEYINPUT38), .B(new_n837), .C1(new_n354), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n834), .A2(new_n836), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n353), .A2(new_n352), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n838), .B1(new_n578), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT40), .B1(new_n827), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n325), .A2(new_n344), .A3(new_n341), .A4(KEYINPUT18), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n347), .A2(new_n577), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n838), .B1(new_n849), .B2(new_n842), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n850), .B2(new_n841), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT40), .B1(new_n851), .B2(new_n839), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n676), .B1(new_n778), .B2(new_n674), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n852), .A2(new_n768), .A3(new_n853), .A4(new_n825), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n411), .A2(new_n853), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(G330), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n816), .B(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n825), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n765), .B(KEYINPUT105), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(new_n772), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n851), .A2(new_n839), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(KEYINPUT39), .B2(new_n845), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n393), .A2(new_n614), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n577), .A2(new_n346), .A3(new_n612), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n864), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n859), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n224), .B2(new_n608), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT35), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n221), .B(new_n222), .C1(new_n498), .C2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n874), .B(G116), .C1(new_n873), .C2(new_n498), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT36), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n331), .A2(G77), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n220), .A2(new_n877), .B1(G50), .B2(new_n211), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(G1), .A3(new_n607), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n872), .A2(new_n876), .A3(new_n879), .ZN(G367));
  NAND2_X1  g0680(.A1(new_n599), .A2(new_n614), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n530), .A2(new_n614), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n523), .A2(new_n533), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n622), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n885), .A2(KEYINPUT42), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n533), .B1(new_n467), .B2(new_n883), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n615), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(KEYINPUT42), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n478), .A2(new_n525), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n614), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n598), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n493), .B2(new_n892), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT43), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n638), .A3(new_n884), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n638), .A2(new_n884), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n890), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n894), .A2(KEYINPUT43), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n900), .B(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n644), .B(KEYINPUT41), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n884), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n624), .B2(new_n630), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT45), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n624), .A2(new_n630), .A3(new_n905), .ZN(new_n909));
  XNOR2_X1  g0709(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT108), .Z(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n909), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n638), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n906), .B(KEYINPUT45), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n909), .B(new_n911), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n916), .A3(new_n639), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n636), .A2(new_n637), .A3(new_n621), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n627), .ZN(new_n919));
  OR3_X1    g0719(.A1(new_n919), .A2(KEYINPUT109), .A3(new_n635), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n635), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT109), .B1(new_n919), .B2(new_n635), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n923), .A2(new_n680), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n914), .A2(new_n917), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n904), .B1(new_n925), .B2(new_n681), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n902), .B1(new_n926), .B2(new_n685), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT110), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(KEYINPUT110), .B(new_n902), .C1(new_n926), .C2(new_n685), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT46), .B1(new_n706), .B2(new_n540), .ZN(new_n932));
  INV_X1    g0732(.A(new_n725), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n720), .A2(new_n550), .B1(new_n933), .B2(G97), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n706), .A2(KEYINPUT46), .A3(G116), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n357), .B1(new_n735), .B2(G311), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n932), .B(new_n937), .C1(G294), .C2(new_n800), .ZN(new_n938));
  INV_X1    g0738(.A(G283), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n753), .A2(new_n939), .B1(new_n741), .B2(new_n395), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT111), .Z(new_n941));
  OAI211_X1 g0741(.A(new_n938), .B(new_n941), .C1(new_n732), .C2(new_n710), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n742), .A2(G68), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n267), .B1(new_n735), .B2(G143), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(new_n202), .C2(new_n753), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(G159), .B2(new_n800), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n719), .A2(new_n784), .B1(new_n749), .B2(new_n705), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G77), .B2(new_n933), .ZN(new_n948));
  INV_X1    g0748(.A(G137), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n946), .B(new_n948), .C1(new_n949), .C2(new_n710), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n942), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT112), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT47), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n698), .ZN(new_n954));
  INV_X1    g0754(.A(new_n689), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n699), .B1(new_n225), .B2(new_n403), .C1(new_n237), .C2(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n894), .A2(new_n762), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n954), .A2(new_n686), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT113), .Z(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n931), .A2(new_n960), .ZN(G387));
  XOR2_X1   g0761(.A(KEYINPUT115), .B(G322), .Z(new_n962));
  AOI22_X1  g0762(.A1(new_n800), .A2(G311), .B1(new_n735), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT116), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n754), .A2(new_n550), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(new_n732), .C2(new_n719), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT48), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n939), .B2(new_n741), .C1(new_n791), .C2(new_n705), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT49), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n757), .A2(G326), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n969), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n357), .B1(new_n933), .B2(new_n540), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n710), .A2(new_n784), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n719), .A2(new_n202), .B1(new_n245), .B2(new_n705), .ZN(new_n976));
  INV_X1    g0776(.A(G159), .ZN(new_n977));
  INV_X1    g0777(.A(new_n735), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n977), .A2(new_n978), .B1(new_n731), .B2(new_n251), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n357), .B1(new_n722), .B2(new_n211), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n976), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n726), .A2(G97), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n741), .A2(new_n403), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n974), .B1(new_n975), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n701), .B1(new_n986), .B2(new_n698), .ZN(new_n987));
  INV_X1    g0787(.A(new_n233), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n955), .B1(new_n988), .B2(G45), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n642), .B1(new_n989), .B2(new_n692), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n252), .A2(new_n202), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT114), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT50), .ZN(new_n993));
  AOI21_X1  g0793(.A(G45), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n993), .B2(new_n992), .C1(new_n211), .C2(new_n245), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n989), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n990), .B(new_n996), .C1(G107), .C2(new_n225), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n699), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n636), .A2(new_n637), .A3(new_n697), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n987), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n923), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n644), .B1(new_n1001), .B2(new_n681), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1000), .B1(new_n684), .B2(new_n923), .C1(new_n1002), .C2(new_n924), .ZN(G393));
  OAI22_X1  g0803(.A1(new_n719), .A2(new_n794), .B1(new_n732), .B2(new_n978), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT52), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n723), .A2(G294), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n357), .B1(new_n757), .B2(new_n962), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n705), .B2(new_n939), .C1(new_n741), .C2(new_n413), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n550), .B2(new_n800), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1005), .A2(new_n748), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n741), .A2(new_n245), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n800), .B2(G50), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n357), .B1(new_n705), .B2(new_n211), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n754), .B2(new_n252), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n757), .A2(G143), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n1014), .A3(new_n803), .A4(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n719), .A2(new_n977), .B1(new_n784), .B2(new_n978), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT51), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n1010), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n701), .B1(new_n1019), .B2(new_n698), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n699), .B1(new_n213), .B2(new_n225), .C1(new_n241), .C2(new_n955), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n762), .C2(new_n884), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n914), .A2(new_n917), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n1023), .B2(new_n684), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n924), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n646), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1024), .B1(new_n1026), .B2(new_n925), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(G390));
  NAND4_X1  g0828(.A1(new_n853), .A2(G330), .A3(new_n768), .A4(new_n825), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n654), .A2(new_n615), .A3(new_n768), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n861), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n867), .B1(new_n1031), .B2(new_n825), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT117), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n1033), .A3(new_n845), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n867), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n861), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n658), .B2(new_n768), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1035), .B(new_n845), .C1(new_n1037), .C2(new_n860), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT117), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n614), .B(new_n769), .C1(new_n595), .C2(new_n603), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n825), .B1(new_n1041), .B2(new_n1036), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n866), .B1(new_n1042), .B2(new_n1035), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1029), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n862), .B2(new_n867), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n779), .A2(G330), .A3(new_n768), .A4(new_n825), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1047), .A2(new_n1039), .A3(new_n1034), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n411), .A2(G330), .A3(new_n853), .ZN(new_n1052));
  OAI211_X1 g0852(.A(G330), .B(new_n768), .C1(new_n675), .C2(new_n826), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n860), .ZN(new_n1054));
  AND3_X1   g0854(.A1(new_n1054), .A2(new_n1037), .A3(new_n1048), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1036), .B1(new_n771), .B2(new_n768), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n860), .B1(new_n679), .B2(new_n769), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n1029), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n815), .B(new_n1052), .C1(new_n1055), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1051), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1044), .A2(new_n1050), .A3(new_n1059), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n644), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(G125), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n357), .B1(new_n202), .B2(new_n725), .C1(new_n711), .C2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT118), .ZN(new_n1066));
  XOR2_X1   g0866(.A(KEYINPUT54), .B(G143), .Z(new_n1067));
  AOI22_X1  g0867(.A1(new_n754), .A2(new_n1067), .B1(new_n720), .B2(G132), .ZN(new_n1068));
  INV_X1    g0868(.A(G128), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n978), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n799), .A2(new_n949), .B1(new_n977), .B2(new_n741), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n706), .A2(G150), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT53), .ZN(new_n1073));
  OR4_X1    g0873(.A1(new_n1066), .A2(new_n1070), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n267), .B1(new_n939), .B2(new_n978), .C1(new_n799), .C2(new_n395), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1011), .B(new_n1075), .C1(G87), .C2(new_n706), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n726), .A2(G68), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n754), .A2(G97), .B1(new_n712), .B2(G294), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n719), .A2(new_n207), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1074), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n701), .B1(new_n1081), .B2(new_n698), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n866), .B2(new_n696), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n251), .B2(new_n807), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1051), .B2(new_n685), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1063), .A2(new_n1085), .ZN(G378));
  NAND2_X1  g0886(.A1(new_n264), .A2(new_n828), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT119), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n309), .A2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(KEYINPUT119), .B(new_n298), .C1(new_n305), .C2(new_n308), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n585), .B1(new_n580), .B2(new_n581), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(KEYINPUT119), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n309), .A2(new_n1091), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n1089), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n855), .B2(G330), .ZN(new_n1101));
  INV_X1    g0901(.A(G330), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1102), .B(new_n1099), .C1(new_n847), .C2(new_n854), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT120), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n870), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n827), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n853), .A2(new_n768), .A3(new_n845), .A4(new_n825), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1107), .A2(new_n852), .B1(new_n1108), .B2(KEYINPUT40), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1099), .B1(new_n1109), .B2(new_n1102), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n855), .A2(G330), .A3(new_n1100), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1110), .A2(new_n870), .A3(new_n1105), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1059), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n815), .A2(new_n1052), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1106), .A2(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT57), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1115), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1061), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1110), .A2(new_n870), .A3(new_n1111), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT122), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n870), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT122), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1110), .A2(new_n870), .A3(new_n1125), .A4(new_n1111), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1120), .A2(new_n1127), .A3(KEYINPUT57), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1118), .A2(new_n644), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n685), .B1(new_n1106), .B2(new_n1113), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1100), .A2(new_n695), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n807), .A2(new_n202), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1064), .A2(new_n978), .B1(new_n731), .B2(new_n789), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n719), .A2(new_n1069), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(new_n706), .C2(new_n1067), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n949), .B2(new_n722), .C1(new_n784), .C2(new_n741), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT59), .Z(new_n1137));
  AOI21_X1  g0937(.A(G41), .B1(new_n933), .B2(G159), .ZN(new_n1138));
  AOI21_X1  g0938(.A(G33), .B1(new_n757), .B2(G124), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n202), .B1(new_n265), .B2(G41), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n933), .A2(G58), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n245), .B2(new_n705), .C1(new_n719), .C2(new_n395), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G283), .B2(new_n712), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n267), .B1(new_n722), .B2(new_n403), .C1(new_n978), .C2(new_n207), .ZN(new_n1145));
  AOI211_X1 g0945(.A(G41), .B(new_n1145), .C1(G97), .C2(new_n730), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n943), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT58), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1140), .A2(new_n1141), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n701), .B1(new_n1149), .B2(new_n698), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1131), .A2(new_n1132), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1130), .A2(KEYINPUT121), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT121), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1110), .A2(new_n1105), .A3(new_n1111), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n1123), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n684), .B1(new_n1155), .B2(new_n1112), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1151), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1153), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1152), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1129), .A2(new_n1159), .ZN(G375));
  NOR2_X1   g0960(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1115), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n903), .A3(new_n1059), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n800), .A2(new_n1067), .B1(G137), .B2(new_n720), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n789), .B2(new_n978), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT123), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n722), .A2(new_n784), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n711), .A2(new_n1069), .B1(new_n977), .B2(new_n705), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(G50), .C2(new_n742), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1166), .A2(new_n357), .A3(new_n1142), .A4(new_n1169), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n267), .B1(new_n791), .B2(new_n978), .C1(new_n799), .C2(new_n413), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n983), .B(new_n1171), .C1(G107), .C2(new_n754), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n712), .A2(G303), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n726), .A2(G77), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n720), .A2(G283), .B1(new_n706), .B2(G97), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1170), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n701), .B1(new_n1177), .B2(new_n698), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n825), .B2(new_n696), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n211), .B2(new_n807), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1161), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n685), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1163), .A2(new_n1182), .ZN(G381));
  NOR4_X1   g0983(.A1(G387), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n1184));
  XOR2_X1   g0984(.A(G375), .B(KEYINPUT124), .Z(new_n1185));
  INV_X1    g0985(.A(G378), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(G384), .A2(G381), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(G407));
  NAND3_X1  g0988(.A1(new_n1185), .A2(new_n613), .A3(new_n1186), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(G407), .A2(G213), .A3(new_n1189), .ZN(G409));
  NAND2_X1  g0990(.A1(G387), .A2(new_n1027), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n931), .A2(new_n960), .A3(G390), .ZN(new_n1192));
  XOR2_X1   g0992(.A(G393), .B(G396), .Z(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(KEYINPUT126), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G390), .B1(new_n931), .B2(new_n960), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n959), .B(new_n1027), .C1(new_n929), .C2(new_n930), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1193), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(KEYINPUT126), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1195), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT60), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n646), .B1(new_n1162), .B2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1202), .B(new_n1059), .C1(new_n1201), .C2(new_n1162), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n813), .B1(new_n1203), .B2(new_n1182), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n813), .A3(new_n1182), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n613), .A2(G213), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1129), .A2(new_n1159), .A3(G378), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1127), .A2(new_n685), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1116), .B2(new_n904), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1186), .B1(new_n1211), .B2(new_n1157), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1209), .A2(KEYINPUT125), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT125), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1207), .B(new_n1208), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT62), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT62), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT61), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1208), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1206), .ZN(new_n1222));
  INV_X1    g1022(.A(G2897), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n1222), .A2(new_n1204), .B1(new_n1223), .B2(new_n1208), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1208), .A2(new_n1223), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1205), .A2(new_n1206), .A3(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1221), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1219), .A2(new_n1220), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1200), .B1(new_n1216), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT63), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1208), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1232), .B2(new_n1227), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1215), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1195), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1218), .A2(new_n1231), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1220), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1230), .B1(new_n1235), .B2(new_n1238), .ZN(G405));
  XNOR2_X1  g1039(.A(new_n1207), .B(KEYINPUT127), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G375), .A2(new_n1186), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1209), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1240), .B(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(new_n1236), .ZN(G402));
endmodule


