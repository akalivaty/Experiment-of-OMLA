//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1330, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1391, new_n1392;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(KEYINPUT64), .A2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(KEYINPUT64), .A2(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G58), .A2(G232), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n213), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT66), .Z(new_n230));
  NOR2_X1   g0030(.A1(new_n213), .A2(G13), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT0), .Z(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n211), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n202), .A2(new_n203), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n233), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  AND3_X1   g0039(.A1(new_n228), .A2(new_n230), .A3(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  INV_X1    g0041(.A(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT2), .B(G226), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G264), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G358));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n250), .B(new_n251), .Z(new_n252));
  XOR2_X1   g0052(.A(G87), .B(G97), .Z(new_n253));
  XNOR2_X1  g0053(.A(G107), .B(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n260), .A2(G222), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n264), .B1(new_n269), .B2(G77), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n263), .B1(new_n262), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G223), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT69), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n269), .B2(new_n261), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n260), .A2(KEYINPUT69), .A3(G1698), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n259), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G179), .ZN(new_n278));
  AND2_X1   g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  OAI21_X1  g0079(.A(G274), .B1(new_n279), .B2(new_n234), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n210), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(G1), .A2(G13), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n210), .A2(new_n288), .B1(new_n289), .B2(new_n257), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n285), .B1(G226), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n277), .A2(new_n278), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(G169), .B1(new_n277), .B2(new_n291), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n234), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT8), .B(G58), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OR3_X1    g0099(.A1(new_n298), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT71), .B1(new_n267), .B2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT71), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(new_n211), .A3(G33), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n299), .A2(new_n300), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G20), .A2(G33), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n296), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n294), .B(new_n234), .C1(G1), .C2(new_n211), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G50), .ZN(new_n310));
  INV_X1    g0110(.A(G13), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n311), .A2(new_n211), .A3(G1), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n201), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n292), .A2(new_n293), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(KEYINPUT9), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT9), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n307), .B2(new_n314), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n277), .A2(G190), .A3(new_n291), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT74), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G200), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n277), .B2(new_n291), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT10), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT73), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT10), .B1(new_n326), .B2(KEYINPUT74), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n326), .A2(KEYINPUT10), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(new_n321), .A3(new_n320), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n316), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT17), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n299), .A2(new_n300), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(new_n309), .ZN(new_n334));
  INV_X1    g0134(.A(new_n312), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AND2_X1   g0137(.A1(KEYINPUT64), .A2(G68), .ZN(new_n338));
  OAI21_X1  g0138(.A(G58), .B1(new_n338), .B2(new_n214), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT77), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT77), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(G58), .C1(new_n338), .C2(new_n214), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n236), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G20), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n260), .A2(new_n345), .A3(G20), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT7), .B1(new_n269), .B2(new_n211), .ZN(new_n347));
  OAI21_X1  g0147(.A(G68), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n305), .A2(G159), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n344), .A2(KEYINPUT16), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n295), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n343), .A2(G20), .B1(G159), .B2(new_n305), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT78), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n267), .B2(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n265), .A2(KEYINPUT78), .A3(G33), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n268), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n345), .A2(G20), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n345), .B1(new_n260), .B2(G20), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n217), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT16), .B1(new_n352), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n337), .B1(new_n351), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT79), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n272), .A2(new_n261), .ZN(new_n365));
  INV_X1    g0165(.A(G226), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G1698), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n266), .A2(new_n365), .A3(new_n268), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G87), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n258), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n258), .A2(G232), .A3(new_n281), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n283), .A2(new_n284), .ZN(new_n373));
  INV_X1    g0173(.A(G274), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n289), .B2(new_n257), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(G200), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  NOR4_X1   g0177(.A1(new_n370), .A2(new_n285), .A3(G190), .A4(new_n371), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n364), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G190), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n372), .A2(new_n380), .A3(new_n376), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n370), .A2(new_n285), .A3(new_n371), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n381), .B(KEYINPUT79), .C1(G200), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n332), .B1(new_n363), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n361), .A2(new_n344), .A3(new_n349), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n359), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n387), .B1(new_n390), .B2(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n296), .B1(new_n352), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n336), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n393), .A2(KEYINPUT17), .A3(new_n379), .A4(new_n383), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n385), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n382), .A2(G179), .ZN(new_n396));
  INV_X1    g0196(.A(G169), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(new_n382), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT18), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n363), .A2(new_n401), .A3(new_n398), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT76), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n215), .A2(G20), .A3(new_n216), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n311), .A2(G1), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT12), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n406), .A2(new_n408), .B1(new_n312), .B2(KEYINPUT12), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n203), .B1(new_n308), .B2(KEYINPUT12), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n301), .A2(new_n303), .A3(G77), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n305), .A2(G50), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n406), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT11), .B1(new_n414), .B2(new_n295), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n405), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n417), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n419), .A2(KEYINPUT76), .A3(new_n415), .A4(new_n411), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT75), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT14), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n373), .A2(new_n375), .B1(new_n290), .B2(G238), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n366), .A2(new_n261), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n242), .A2(G1698), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n266), .A2(new_n425), .A3(new_n268), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n259), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT13), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n424), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n424), .B2(new_n430), .ZN(new_n433));
  OAI211_X1 g0233(.A(G169), .B(new_n423), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n290), .A2(G238), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n376), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n258), .B1(new_n427), .B2(new_n428), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT13), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n424), .A2(new_n430), .A3(new_n431), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(G179), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n439), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n423), .B1(new_n442), .B2(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n421), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n219), .B1(new_n274), .B2(new_n275), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n260), .A2(G232), .A3(new_n261), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n207), .B2(new_n260), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n259), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT72), .ZN(new_n449));
  INV_X1    g0249(.A(new_n290), .ZN(new_n450));
  INV_X1    g0250(.A(G244), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n452), .B2(new_n285), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n376), .B(KEYINPUT72), .C1(new_n451), .C2(new_n450), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n448), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n455), .A2(G200), .ZN(new_n456));
  INV_X1    g0256(.A(G77), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n312), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n457), .B2(new_n308), .ZN(new_n459));
  INV_X1    g0259(.A(new_n297), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n460), .A2(new_n305), .B1(G20), .B2(G77), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n211), .A2(G33), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT15), .B(G87), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n459), .B1(new_n464), .B2(new_n295), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n455), .B2(new_n380), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n456), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n438), .A2(G190), .A3(new_n439), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n416), .A2(new_n417), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n432), .A2(new_n433), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n468), .B(new_n469), .C1(new_n470), .C2(new_n323), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n465), .B1(new_n455), .B2(new_n397), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n448), .A2(new_n453), .A3(new_n278), .A4(new_n454), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND4_X1   g0274(.A1(new_n444), .A2(new_n467), .A3(new_n471), .A4(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n331), .A2(new_n404), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT80), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT80), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n331), .A2(new_n478), .A3(new_n404), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n266), .A2(new_n268), .A3(G244), .A4(new_n261), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n488), .A2(new_n259), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n287), .A2(G1), .ZN(new_n490));
  AND2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NOR2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(G257), .A3(new_n258), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT5), .B(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n375), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n397), .B1(new_n489), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n488), .A2(new_n259), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT84), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT84), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n499), .A2(new_n501), .A3(new_n278), .A4(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n360), .A2(G107), .B1(G77), .B2(new_n305), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G97), .A2(G107), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT81), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  AND2_X1   g0308(.A1(KEYINPUT6), .A2(G107), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n208), .B(new_n506), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT82), .ZN(new_n511));
  INV_X1    g0311(.A(new_n506), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n512), .A2(new_n513), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n510), .B2(new_n514), .ZN(new_n516));
  OAI21_X1  g0316(.A(G20), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n296), .B1(new_n505), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT86), .ZN(new_n519));
  OR3_X1    g0319(.A1(new_n335), .A2(KEYINPUT83), .A3(G97), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT83), .B1(new_n335), .B2(G97), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n267), .A2(G1), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n312), .A2(new_n295), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n520), .A2(new_n521), .B1(G97), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n510), .A2(new_n514), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n211), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n305), .A2(G77), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n265), .A2(G33), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n211), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n345), .A2(new_n534), .B1(new_n356), .B2(new_n357), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n531), .B1(new_n535), .B2(new_n207), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n295), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT86), .B1(new_n537), .B2(new_n524), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n504), .B1(new_n526), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT85), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n518), .A2(new_n525), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n497), .B1(new_n488), .B2(new_n259), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT85), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n540), .A2(new_n546), .A3(G200), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n542), .A2(new_n543), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n539), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n428), .ZN(new_n550));
  AND2_X1   g0350(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n551));
  NOR2_X1   g0351(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G87), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n553), .A2(new_n211), .B1(new_n554), .B2(new_n513), .ZN(new_n555));
  OR2_X1    g0355(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n556));
  NAND2_X1  g0356(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n556), .B(new_n557), .C1(new_n462), .C2(new_n206), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n266), .A2(new_n268), .A3(new_n211), .A4(G68), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n295), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n463), .A2(new_n312), .ZN(new_n562));
  INV_X1    g0362(.A(new_n463), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n523), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT88), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT88), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n561), .A2(new_n567), .A3(new_n562), .A4(new_n564), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n375), .A2(new_n490), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n210), .A2(G45), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n258), .A2(G250), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n266), .A2(new_n268), .A3(G244), .A4(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n266), .A2(new_n268), .A3(G238), .A4(new_n261), .ZN(new_n574));
  INV_X1    g0374(.A(G116), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n267), .C2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n572), .B1(new_n576), .B2(new_n259), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n278), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n259), .ZN(new_n579));
  INV_X1    g0379(.A(new_n572), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n397), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n566), .A2(new_n568), .A3(new_n578), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(G190), .A3(new_n580), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT89), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n577), .A2(KEYINPUT89), .A3(G190), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n523), .A2(G87), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n561), .A2(new_n562), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n581), .A2(G200), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n586), .A2(new_n587), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n549), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n493), .A2(G264), .A3(new_n258), .ZN(new_n594));
  INV_X1    g0394(.A(G294), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n267), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(G250), .A2(G1698), .ZN(new_n597));
  INV_X1    g0397(.A(G257), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(new_n599), .B2(new_n260), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n259), .B1(new_n600), .B2(KEYINPUT92), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(G1698), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G250), .B2(G1698), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n603), .A2(new_n269), .B1(new_n267), .B2(new_n595), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT92), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n496), .B(new_n594), .C1(new_n601), .C2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT93), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n605), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n600), .A2(KEYINPUT92), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(new_n259), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n612), .A2(KEYINPUT93), .A3(new_n496), .A4(new_n594), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(G169), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n607), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G179), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n260), .A2(new_n211), .A3(G87), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT22), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT22), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n260), .A2(new_n620), .A3(new_n211), .A4(G87), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n267), .A2(new_n575), .A3(G20), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT23), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n211), .B2(G107), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT24), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT24), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n622), .A2(new_n630), .A3(new_n627), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n295), .ZN(new_n633));
  INV_X1    g0433(.A(new_n523), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n312), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT25), .B1(new_n312), .B2(new_n207), .ZN(new_n636));
  OAI22_X1  g0436(.A1(new_n634), .A2(new_n207), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n617), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n632), .B2(new_n295), .ZN(new_n641));
  AOI21_X1  g0441(.A(G190), .B1(new_n609), .B2(new_n613), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n615), .A2(G200), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n266), .A2(new_n268), .A3(G257), .A4(new_n261), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT91), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT91), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n260), .A2(new_n647), .A3(G257), .A4(new_n261), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n266), .A2(new_n268), .A3(G1698), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n650), .A2(G264), .B1(G303), .B2(new_n269), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n259), .ZN(new_n653));
  INV_X1    g0453(.A(new_n496), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n493), .A2(G270), .A3(new_n258), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT90), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n493), .A2(KEYINPUT90), .A3(G270), .A4(new_n258), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n335), .A2(G116), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n523), .B2(G116), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n487), .B(new_n211), .C1(G33), .C2(new_n206), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n575), .A2(G20), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n295), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT20), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n663), .A2(KEYINPUT20), .A3(new_n295), .A4(new_n664), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n660), .A2(new_n670), .A3(new_n278), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n397), .B1(new_n662), .B2(new_n669), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n660), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT21), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT21), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n660), .A2(new_n675), .A3(new_n672), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n671), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n660), .A2(G200), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n678), .B(new_n670), .C1(new_n380), .C2(new_n660), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n640), .A2(new_n644), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n481), .A2(new_n593), .A3(new_n680), .ZN(G372));
  NAND2_X1  g0481(.A1(new_n640), .A2(new_n677), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n549), .A2(new_n591), .A3(new_n682), .A4(new_n644), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT94), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n577), .B2(G169), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n581), .A2(KEYINPUT94), .A3(new_n397), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(new_n565), .A4(new_n578), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT26), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n591), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n498), .B(new_n503), .C1(new_n518), .C2(new_n525), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(KEYINPUT95), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n498), .A2(new_n503), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n519), .B1(new_n518), .B2(new_n525), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n537), .A2(KEYINPUT86), .A3(new_n524), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n592), .A3(KEYINPUT26), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT95), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n698), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n692), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n683), .A2(new_n687), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n480), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n400), .A2(new_n402), .ZN(new_n703));
  INV_X1    g0503(.A(new_n471), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n444), .B1(new_n704), .B2(new_n474), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n706), .B2(new_n395), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n325), .A2(new_n330), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n316), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n702), .A2(new_n710), .ZN(G369));
  NAND2_X1  g0511(.A1(new_n674), .A2(new_n676), .ZN(new_n712));
  INV_X1    g0512(.A(new_n671), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT27), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n407), .A2(new_n715), .A3(new_n211), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT96), .Z(new_n717));
  INV_X1    g0517(.A(G213), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n407), .A2(new_n211), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(KEYINPUT27), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G343), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n670), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT97), .B1(new_n714), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n677), .A2(new_n679), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(new_n725), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n714), .A2(KEYINPUT97), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(KEYINPUT98), .A3(G330), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT98), .ZN(new_n733));
  INV_X1    g0533(.A(G330), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n640), .B(new_n644), .C1(new_n641), .C2(new_n724), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n617), .A2(new_n639), .A3(new_n723), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT99), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n737), .A2(KEYINPUT99), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n677), .A2(new_n723), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n741), .B2(new_n742), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n640), .A2(new_n723), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n744), .A2(new_n749), .ZN(G399));
  INV_X1    g0550(.A(KEYINPUT100), .ZN(new_n751));
  INV_X1    g0551(.A(new_n231), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n752), .B2(G41), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n231), .A2(KEYINPUT100), .A3(new_n286), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(G1), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(new_n237), .B2(new_n755), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT28), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n640), .A2(new_n677), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n539), .A2(new_n644), .A3(new_n548), .A4(new_n591), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n687), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n689), .A2(new_n690), .A3(new_n688), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n696), .A2(new_n592), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n763), .B1(new_n688), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n724), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(KEYINPUT29), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n594), .B1(new_n601), .B2(new_n606), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n579), .A2(G179), .A3(new_n580), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n657), .A2(new_n658), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n496), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n258), .B1(new_n649), .B2(new_n651), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n770), .A2(new_n774), .A3(KEYINPUT30), .A4(new_n544), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT30), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n544), .A2(new_n653), .A3(new_n659), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n612), .A2(new_n577), .A3(G179), .A4(new_n594), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n577), .A2(G179), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n660), .A2(new_n540), .A3(new_n780), .A4(new_n607), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n775), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n723), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT31), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(KEYINPUT31), .A3(new_n723), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n539), .A2(new_n548), .A3(new_n592), .A4(new_n724), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n785), .B(new_n786), .C1(new_n680), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G330), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT29), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n701), .A2(new_n790), .A3(new_n724), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n767), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n759), .B1(new_n793), .B2(G1), .ZN(G364));
  INV_X1    g0594(.A(new_n755), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n311), .A2(G20), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n210), .B1(new_n796), .B2(G45), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n231), .A2(new_n260), .ZN(new_n800));
  INV_X1    g0600(.A(G355), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n801), .B1(G116), .B2(new_n231), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n752), .A2(new_n260), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n287), .B2(new_n238), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n252), .A2(new_n287), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G13), .A2(G33), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n234), .B1(G20), .B2(new_n397), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n799), .B1(new_n807), .B2(new_n813), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n380), .A2(G179), .A3(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n211), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n211), .A2(new_n278), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G190), .A2(G200), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n817), .A2(G294), .B1(new_n821), .B2(G311), .ZN(new_n822));
  INV_X1    g0622(.A(G326), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n818), .A2(G200), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n380), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n822), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT101), .Z(new_n828));
  NAND3_X1  g0628(.A1(new_n818), .A2(G190), .A3(new_n323), .ZN(new_n829));
  INV_X1    g0629(.A(G322), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n269), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n211), .A2(G179), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n819), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(G329), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n824), .A2(G190), .ZN(new_n836));
  INV_X1    g0636(.A(G317), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT33), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(KEYINPUT33), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n832), .A2(G190), .A3(G200), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n832), .A2(new_n380), .A3(G200), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n842), .A2(G303), .B1(new_n844), .B2(G283), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n828), .A2(new_n835), .A3(new_n840), .A4(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT102), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n841), .A2(new_n554), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n834), .A2(G159), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(KEYINPUT32), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(G68), .C2(new_n836), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n260), .B1(new_n820), .B2(new_n457), .ZN(new_n853));
  INV_X1    g0653(.A(new_n829), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(G58), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n843), .A2(new_n207), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n850), .B2(KEYINPUT32), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G97), .A2(new_n817), .B1(new_n825), .B2(G50), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n852), .A2(new_n855), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n846), .A2(new_n847), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n848), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n814), .B1(new_n861), .B2(new_n811), .ZN(new_n862));
  INV_X1    g0662(.A(new_n810), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n731), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n799), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n731), .B2(G330), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n864), .B1(new_n736), .B2(new_n866), .ZN(G396));
  NAND3_X1  g0667(.A1(new_n467), .A2(new_n474), .A3(new_n724), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n701), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n687), .ZN(new_n871));
  INV_X1    g0671(.A(new_n761), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n682), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n723), .B1(new_n873), .B2(new_n700), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n472), .A2(new_n473), .A3(new_n724), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n456), .A2(new_n466), .B1(new_n465), .B2(new_n724), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n876), .B2(new_n474), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n870), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n799), .B1(new_n878), .B2(new_n789), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n789), .B2(new_n878), .ZN(new_n880));
  INV_X1    g0680(.A(new_n811), .ZN(new_n881));
  INV_X1    g0681(.A(G132), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n260), .B1(new_n833), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(G50), .B2(new_n842), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n817), .A2(G58), .B1(new_n844), .B2(G68), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n854), .A2(G143), .B1(new_n821), .B2(G159), .ZN(new_n886));
  INV_X1    g0686(.A(G137), .ZN(new_n887));
  INV_X1    g0687(.A(G150), .ZN(new_n888));
  INV_X1    g0688(.A(new_n836), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n886), .B1(new_n826), .B2(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT34), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n884), .B(new_n885), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n889), .A2(KEYINPUT103), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n889), .A2(KEYINPUT103), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(G283), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n817), .A2(G97), .B1(new_n844), .B2(G87), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n825), .A2(G303), .B1(new_n842), .B2(G107), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n260), .B1(new_n854), .B2(G294), .ZN(new_n901));
  AOI22_X1  g0701(.A1(G116), .A2(new_n821), .B1(new_n834), .B2(G311), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n899), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n892), .A2(new_n893), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n881), .B1(new_n904), .B2(KEYINPUT104), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(KEYINPUT104), .B2(new_n904), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n881), .A2(new_n809), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n906), .B(new_n799), .C1(G77), .C2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT105), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n809), .B2(new_n877), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n880), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(G384));
  NOR2_X1   g0712(.A1(new_n515), .A2(new_n516), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n914), .A2(KEYINPUT35), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(KEYINPUT35), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n915), .A2(new_n916), .A3(G116), .A4(new_n235), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT36), .Z(new_n918));
  NAND4_X1  g0718(.A1(new_n340), .A2(G77), .A3(new_n238), .A4(new_n342), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n201), .A2(G68), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n210), .B(G13), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n344), .A2(new_n349), .A3(new_n348), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n387), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n336), .B1(new_n924), .B2(new_n392), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n363), .A2(new_n384), .B1(new_n925), .B2(new_n721), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n399), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT37), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n393), .A2(new_n379), .A3(new_n383), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n363), .A2(new_n398), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n721), .B(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n363), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT37), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n929), .A2(new_n930), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n925), .A2(new_n721), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n395), .B2(new_n403), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n935), .A2(new_n937), .A3(KEYINPUT38), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n935), .B2(new_n937), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT108), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n937), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT38), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT108), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n935), .A2(new_n937), .A3(KEYINPUT38), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n444), .A2(KEYINPUT106), .A3(new_n471), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n418), .A2(new_n723), .A3(new_n420), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n471), .ZN(new_n950));
  INV_X1    g0750(.A(new_n423), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n470), .B2(new_n397), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(new_n440), .A3(new_n434), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT106), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n444), .A2(new_n955), .A3(new_n471), .ZN(new_n956));
  INV_X1    g0756(.A(new_n949), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n948), .A2(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND4_X1   g0758(.A1(KEYINPUT110), .A2(new_n788), .A3(new_n877), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n948), .A2(new_n954), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n956), .A2(new_n957), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n960), .A2(new_n961), .A3(new_n877), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT110), .B1(new_n962), .B2(new_n788), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT40), .B1(new_n947), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n932), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT109), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n385), .A2(new_n967), .A3(new_n394), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n703), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n967), .B1(new_n385), .B2(new_n394), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT37), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n934), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n942), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n945), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n680), .A2(new_n787), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n785), .A2(new_n786), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT40), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n960), .A2(new_n961), .A3(new_n877), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n965), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n481), .A2(new_n980), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n734), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n984), .B2(new_n985), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n953), .A2(new_n421), .A3(new_n724), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n943), .A2(KEYINPUT39), .A3(new_n945), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n938), .B1(new_n975), .B2(new_n942), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n989), .B(new_n990), .C1(new_n991), .C2(KEYINPUT39), .ZN(new_n992));
  INV_X1    g0792(.A(new_n958), .ZN(new_n993));
  INV_X1    g0793(.A(new_n875), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n870), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n947), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n703), .A2(new_n931), .ZN(new_n997));
  AND3_X1   g0797(.A1(new_n992), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n710), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n767), .A2(new_n791), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n480), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n998), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n987), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n210), .B2(new_n796), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n987), .A2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n922), .B1(new_n1004), .B2(new_n1005), .ZN(G367));
  OAI21_X1  g0806(.A(new_n723), .B1(new_n518), .B2(new_n525), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n693), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n549), .A2(new_n1007), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT111), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n549), .A2(KEYINPUT111), .A3(new_n1007), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n747), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n539), .B1(new_n1013), .B2(new_n640), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1015), .A2(KEYINPUT42), .B1(new_n1016), .B2(new_n724), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1015), .A2(KEYINPUT42), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n724), .A2(new_n589), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n871), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n689), .B2(new_n1019), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1017), .A2(new_n1018), .B1(KEYINPUT43), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(KEYINPUT43), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n744), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n1014), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1024), .B(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n755), .B(KEYINPUT41), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT113), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n743), .A2(new_n745), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n748), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n1014), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT112), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT112), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n749), .A2(new_n1034), .A3(new_n1014), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(KEYINPUT45), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT44), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n749), .B2(new_n1014), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1013), .B(KEYINPUT44), .C1(new_n747), .C2(new_n748), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT45), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1029), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n744), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1029), .B(new_n1025), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n736), .B(KEYINPUT115), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n747), .A2(KEYINPUT114), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n743), .B2(new_n745), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n743), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(KEYINPUT114), .A3(new_n746), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(KEYINPUT115), .B1(new_n732), .B2(new_n735), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1048), .A2(new_n1053), .A3(new_n1050), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n792), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1044), .A2(new_n1045), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1028), .B1(new_n1056), .B2(new_n793), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1027), .B1(new_n1057), .B2(new_n798), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1021), .A2(new_n863), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n896), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(G159), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n820), .A2(new_n201), .B1(new_n833), .B2(new_n887), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n269), .B(new_n1062), .C1(G150), .C2(new_n854), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n825), .A2(G143), .B1(new_n844), .B2(G77), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n817), .A2(G68), .B1(new_n842), .B2(G58), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n841), .A2(new_n575), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT46), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(KEYINPUT46), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n896), .C2(new_n595), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(KEYINPUT116), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n817), .A2(G107), .B1(new_n844), .B2(G97), .ZN(new_n1072));
  INV_X1    g0872(.A(G311), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1072), .B1(new_n1073), .B2(new_n826), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n269), .B1(new_n833), .B2(new_n837), .ZN(new_n1075));
  INV_X1    g0875(.A(G303), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n829), .A2(new_n1076), .B1(new_n820), .B2(new_n897), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1071), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1070), .A2(KEYINPUT116), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1066), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT47), .Z(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n881), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n803), .A2(new_n248), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n813), .B1(new_n752), .B2(new_n563), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n865), .B(new_n1083), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT117), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1059), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1058), .A2(new_n1089), .ZN(G387));
  OAI22_X1  g0890(.A1(new_n800), .A2(new_n756), .B1(G107), .B2(new_n231), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n245), .A2(new_n287), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n756), .ZN(new_n1093));
  AOI211_X1 g0893(.A(G45), .B(new_n1093), .C1(G68), .C2(G77), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n297), .A2(G50), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT50), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n804), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1091), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n269), .B1(new_n833), .B2(new_n823), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n854), .A2(G317), .B1(new_n821), .B2(G303), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n830), .B2(new_n826), .C1(new_n896), .C2(new_n1073), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT48), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n817), .A2(G283), .B1(new_n842), .B2(G294), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT49), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1099), .B(new_n1108), .C1(G116), .C2(new_n844), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n269), .B1(new_n834), .B2(G150), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n457), .B2(new_n841), .C1(new_n206), .C2(new_n843), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT118), .Z(new_n1113));
  AOI22_X1  g0913(.A1(new_n854), .A2(G50), .B1(new_n821), .B2(G68), .ZN(new_n1114));
  INV_X1    g0914(.A(G159), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1114), .B1(new_n463), .B2(new_n816), .C1(new_n1115), .C2(new_n826), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n333), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n836), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1109), .A2(new_n1110), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n799), .B1(new_n813), .B2(new_n1098), .C1(new_n1119), .C2(new_n881), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1049), .B2(new_n810), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n798), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1055), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n795), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1122), .A2(new_n793), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(G393));
  AND2_X1   g0927(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT45), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1032), .A2(KEYINPUT112), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1034), .B1(new_n749), .B2(new_n1014), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1128), .A2(KEYINPUT119), .A3(new_n744), .A4(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1132), .A2(new_n744), .A3(new_n1040), .A4(new_n1036), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT119), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1025), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1133), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n795), .B(new_n1056), .C1(new_n1138), .C2(new_n1055), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1013), .A2(new_n810), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n812), .B1(new_n206), .B2(new_n231), .C1(new_n804), .C2(new_n255), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n799), .A2(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n826), .A2(new_n837), .B1(new_n1073), .B2(new_n829), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT52), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n856), .B1(G116), .B2(new_n817), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n897), .B2(new_n841), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n269), .B1(new_n833), .B2(new_n830), .C1(new_n595), .C2(new_n820), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1144), .B(new_n1148), .C1(new_n1076), .C2(new_n896), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n826), .A2(new_n888), .B1(new_n1115), .B2(new_n829), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT51), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n817), .A2(G77), .B1(new_n821), .B2(new_n460), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(new_n201), .C2(new_n896), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n269), .B1(new_n834), .B2(G143), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n554), .B2(new_n843), .C1(new_n218), .C2(new_n841), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT120), .Z(new_n1156));
  OAI21_X1  g0956(.A(new_n1149), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1142), .B1(new_n1157), .B2(new_n811), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1138), .A2(new_n798), .B1(new_n1140), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1139), .A2(new_n1159), .ZN(G390));
  NAND3_X1  g0960(.A1(new_n480), .A2(G330), .A3(new_n788), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n876), .A2(new_n474), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n724), .B(new_n1162), .C1(new_n762), .C2(new_n765), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n994), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n788), .A2(G330), .A3(new_n877), .A4(new_n958), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n877), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n993), .B1(new_n789), .B2(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n875), .B1(new_n701), .B2(new_n869), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1168), .B2(new_n1166), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1001), .B(new_n1161), .C1(new_n1169), .C2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT39), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT38), .B1(new_n971), .B2(new_n974), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n938), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n868), .B1(new_n873), .B2(new_n700), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n958), .B1(new_n1176), .B2(new_n875), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1175), .A2(new_n990), .B1(new_n1177), .B2(new_n988), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n993), .B1(new_n1163), .B2(new_n994), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1179), .A2(new_n991), .A3(new_n989), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1166), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1175), .A2(new_n990), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1177), .A2(new_n988), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n977), .B(new_n988), .C1(new_n1165), .C2(new_n993), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1166), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1172), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1168), .A2(new_n1166), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1171), .B1(new_n1165), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1000), .A2(new_n480), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n710), .A3(new_n1161), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1181), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1185), .A2(new_n1186), .A3(new_n1166), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1188), .A2(new_n795), .A3(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n798), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1183), .A2(new_n808), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n799), .B1(new_n1117), .B2(new_n907), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1060), .A2(G107), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n269), .B1(new_n829), .B2(new_n575), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G97), .B2(new_n821), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n825), .A2(G283), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n849), .B1(G77), .B2(new_n817), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n843), .A2(new_n203), .B1(new_n833), .B2(new_n595), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT122), .Z(new_n1208));
  NOR2_X1   g1008(.A1(new_n829), .A2(new_n882), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n269), .B(new_n1209), .C1(G125), .C2(new_n834), .ZN(new_n1210));
  OAI21_X1  g1010(.A(KEYINPUT53), .B1(new_n841), .B2(new_n888), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT54), .B(G143), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT121), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n821), .ZN(new_n1214));
  OR3_X1    g1014(.A1(new_n841), .A2(KEYINPUT53), .A3(new_n888), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1210), .A2(new_n1211), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n825), .A2(G128), .B1(new_n844), .B2(G50), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n1115), .B2(new_n816), .C1(new_n896), .C2(new_n887), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1206), .A2(new_n1208), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1200), .B1(new_n1219), .B2(new_n811), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1199), .A2(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1198), .A2(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1197), .A2(KEYINPUT123), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT123), .B1(new_n1197), .B2(new_n1222), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(G378));
  AOI21_X1  g1025(.A(new_n734), .B1(new_n977), .B2(new_n983), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n315), .A2(new_n721), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n331), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n331), .A2(new_n1229), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1227), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1232), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1227), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1234), .A2(new_n1230), .A3(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT110), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n980), .B2(new_n982), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n962), .A2(KEYINPUT110), .A3(new_n788), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n940), .B2(new_n946), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1226), .B(new_n1237), .C1(new_n1242), .C2(KEYINPUT40), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n983), .ZN(new_n1245));
  OAI21_X1  g1045(.A(G330), .B1(new_n1245), .B2(new_n991), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n965), .B2(new_n1246), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1243), .A2(new_n1247), .A3(new_n998), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n998), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n798), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1244), .A2(new_n808), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n799), .B1(G50), .B2(new_n907), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n854), .A2(G128), .B1(new_n821), .B2(G137), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n882), .B2(new_n889), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G150), .A2(new_n817), .B1(new_n825), .B2(G125), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT124), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(new_n842), .C2(new_n1213), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT59), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n844), .A2(G159), .ZN(new_n1261));
  AOI211_X1 g1061(.A(G33), .B(G41), .C1(new_n834), .C2(G124), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n889), .A2(new_n206), .B1(new_n202), .B2(new_n843), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G116), .B2(new_n825), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n269), .A2(new_n286), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G283), .B2(new_n834), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n854), .A2(G107), .B1(new_n821), .B2(new_n563), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n817), .A2(G68), .B1(new_n842), .B2(G77), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1265), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT58), .ZN(new_n1271));
  OR2_X1    g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1266), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1263), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1252), .B1(new_n1275), .B2(new_n811), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1251), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1250), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT57), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1192), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1196), .A2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n795), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n992), .A2(new_n996), .A3(new_n997), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n947), .A2(new_n964), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n981), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1237), .B1(new_n1286), .B2(new_n1226), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n965), .A2(new_n1246), .A3(new_n1244), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1284), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1243), .A2(new_n1247), .A3(new_n998), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1196), .A2(new_n1281), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT57), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1279), .B1(new_n1283), .B2(new_n1293), .ZN(G375));
  NAND2_X1  g1094(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1028), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1172), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1297), .B(KEYINPUT125), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1060), .A2(new_n1213), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n269), .B1(new_n854), .B2(G137), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(G150), .A2(new_n821), .B1(new_n834), .B2(G128), .ZN(new_n1301));
  OAI22_X1  g1101(.A1(new_n826), .A2(new_n882), .B1(new_n202), .B2(new_n843), .ZN(new_n1302));
  OAI22_X1  g1102(.A1(new_n816), .A2(new_n201), .B1(new_n841), .B2(new_n1115), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1060), .A2(G116), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n829), .A2(new_n897), .B1(new_n820), .B2(new_n207), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n260), .B(new_n1307), .C1(G303), .C2(new_n834), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n817), .A2(new_n563), .B1(new_n844), .B2(G77), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n825), .A2(G294), .B1(new_n842), .B2(G97), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1306), .A2(new_n1308), .A3(new_n1309), .A4(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1305), .A2(new_n1311), .ZN(new_n1312));
  OAI221_X1 g1112(.A(new_n799), .B1(G68), .B2(new_n907), .C1(new_n1312), .C2(new_n881), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1313), .B1(new_n993), .B2(new_n808), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1190), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1315), .B2(new_n798), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1298), .A2(new_n1316), .ZN(G381));
  NOR4_X1   g1117(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1318));
  INV_X1    g1118(.A(G390), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1197), .A2(new_n1222), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT57), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n755), .B1(new_n1325), .B2(new_n1292), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1278), .B1(new_n1324), .B2(new_n1326), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1318), .A2(new_n1319), .A3(new_n1321), .A4(new_n1327), .ZN(new_n1328));
  OR2_X1    g1128(.A1(new_n1328), .A2(G387), .ZN(G407));
  NAND3_X1  g1129(.A1(new_n1327), .A2(new_n722), .A3(new_n1321), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(G407), .A2(G213), .A3(new_n1330), .ZN(G409));
  XNOR2_X1  g1131(.A(G393), .B(G396), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1058), .A2(G390), .A3(new_n1089), .ZN(new_n1333));
  AOI21_X1  g1133(.A(G390), .B1(new_n1058), .B2(new_n1089), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1332), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(G387), .A2(new_n1319), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1332), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1058), .A2(G390), .A3(new_n1089), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1336), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1335), .A2(new_n1339), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n718), .A2(G343), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT123), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1320), .A2(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1197), .A2(KEYINPUT123), .A3(new_n1222), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(G375), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT126), .ZN(new_n1348));
  AOI22_X1  g1148(.A1(new_n1289), .A2(new_n1290), .B1(new_n1196), .B2(new_n1281), .ZN(new_n1349));
  AOI22_X1  g1149(.A1(new_n1278), .A2(new_n1348), .B1(new_n1296), .B2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1250), .A2(KEYINPUT126), .A3(new_n1277), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1320), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1342), .B1(new_n1347), .B2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT60), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1295), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n795), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1354), .B1(new_n1172), .B2(new_n1295), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1316), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1358));
  OR2_X1    g1158(.A1(new_n1358), .A2(new_n911), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n911), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1341), .A2(G2897), .ZN(new_n1362));
  XNOR2_X1  g1162(.A(new_n1361), .B(new_n1362), .ZN(new_n1363));
  AOI21_X1  g1163(.A(KEYINPUT61), .B1(new_n1353), .B2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1327), .A2(G378), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n797), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1277), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1348), .B1(new_n1366), .B2(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1349), .A2(new_n1296), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1368), .A2(new_n1351), .A3(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1370), .A2(new_n1321), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1341), .B1(new_n1365), .B2(new_n1371), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1361), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1372), .A2(KEYINPUT63), .A3(new_n1373), .ZN(new_n1374));
  OAI211_X1 g1174(.A(new_n1342), .B(new_n1373), .C1(new_n1347), .C2(new_n1352), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT63), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1375), .A2(new_n1376), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1340), .A2(new_n1364), .A3(new_n1374), .A4(new_n1377), .ZN(new_n1378));
  AOI21_X1  g1178(.A(KEYINPUT62), .B1(new_n1372), .B2(new_n1373), .ZN(new_n1379));
  AOI22_X1  g1179(.A1(new_n1327), .A2(G378), .B1(new_n1370), .B2(new_n1321), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT62), .ZN(new_n1381));
  NOR4_X1   g1181(.A1(new_n1380), .A2(new_n1381), .A3(new_n1341), .A4(new_n1361), .ZN(new_n1382));
  OAI211_X1 g1182(.A(new_n1364), .B(KEYINPUT127), .C1(new_n1379), .C2(new_n1382), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1335), .A2(new_n1339), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1383), .A2(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1375), .A2(new_n1381), .ZN(new_n1386));
  NAND3_X1  g1186(.A1(new_n1372), .A2(KEYINPUT62), .A3(new_n1373), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1386), .A2(new_n1387), .ZN(new_n1388));
  AOI21_X1  g1188(.A(KEYINPUT127), .B1(new_n1388), .B2(new_n1364), .ZN(new_n1389));
  OAI21_X1  g1189(.A(new_n1378), .B1(new_n1385), .B2(new_n1389), .ZN(G405));
  OAI21_X1  g1190(.A(new_n1365), .B1(new_n1320), .B2(new_n1327), .ZN(new_n1391));
  XNOR2_X1  g1191(.A(new_n1391), .B(new_n1373), .ZN(new_n1392));
  XNOR2_X1  g1192(.A(new_n1392), .B(new_n1384), .ZN(G402));
endmodule


