//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT72), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  AOI21_X1  g008(.A(G128), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(KEYINPUT1), .A3(G146), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n190), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n192), .A2(new_n194), .A3(new_n199), .A4(G128), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n196), .B(KEYINPUT67), .C1(new_n201), .C2(G128), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n198), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT3), .A3(G104), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT73), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n207), .B2(G104), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(KEYINPUT73), .A3(G107), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n209), .A2(new_n210), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n205), .A2(G107), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n207), .A2(G104), .ZN(new_n216));
  OAI21_X1  g030(.A(G101), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n203), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n214), .A2(new_n217), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n200), .B(new_n196), .C1(G128), .C2(new_n201), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT11), .B1(new_n224), .B2(G134), .ZN(new_n225));
  INV_X1    g039(.A(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G137), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G137), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT11), .A4(G134), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n227), .A2(new_n228), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n228), .B1(new_n227), .B2(new_n232), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT12), .B1(new_n223), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT12), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n233), .A2(new_n234), .ZN(new_n238));
  AOI211_X1 g052(.A(new_n237), .B(new_n238), .C1(new_n219), .C2(new_n222), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT10), .B1(new_n203), .B2(new_n218), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT10), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n220), .A2(new_n242), .A3(new_n221), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT74), .A2(G101), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(KEYINPUT4), .A3(new_n247), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT0), .A4(G128), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n201), .A2(KEYINPUT64), .A3(KEYINPUT0), .A4(G128), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT0), .B(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n201), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT68), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n258), .B1(new_n254), .B2(new_n255), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n251), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n244), .A2(new_n238), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n244), .A2(new_n265), .A3(KEYINPUT75), .A4(new_n238), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n240), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G140), .ZN(new_n272));
  INV_X1    g086(.A(G953), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n273), .A2(G227), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n272), .B(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n270), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n244), .A2(new_n265), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n235), .ZN(new_n279));
  AOI211_X1 g093(.A(KEYINPUT68), .B(new_n258), .C1(new_n254), .C2(new_n255), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n263), .B1(new_n256), .B2(new_n259), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n282), .A2(new_n251), .B1(new_n241), .B2(new_n243), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT75), .B1(new_n283), .B2(new_n238), .ZN(new_n284));
  INV_X1    g098(.A(new_n269), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n279), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT76), .B1(new_n286), .B2(new_n275), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n268), .A2(new_n269), .ZN(new_n288));
  INV_X1    g102(.A(new_n240), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n288), .A2(new_n276), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n277), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n288), .A2(new_n276), .A3(new_n279), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n295), .B(G469), .C1(new_n276), .C2(new_n270), .ZN(new_n296));
  NAND2_X1  g110(.A1(G469), .A2(G902), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n189), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n300), .B(KEYINPUT77), .Z(new_n301));
  NOR2_X1   g115(.A1(G237), .A2(G953), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n302), .A2(G143), .A3(G214), .ZN(new_n303));
  AOI21_X1  g117(.A(G143), .B1(new_n302), .B2(G214), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT18), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n306), .A2(new_n228), .A3(KEYINPUT82), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n305), .B(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n309), .B1(new_n314), .B2(G146), .ZN(new_n315));
  XNOR2_X1  g129(.A(G125), .B(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(KEYINPUT70), .A3(new_n191), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n318), .B1(new_n191), .B2(new_n316), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n308), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n305), .A2(new_n228), .ZN(new_n321));
  OAI21_X1  g135(.A(G131), .B1(new_n303), .B2(new_n304), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(KEYINPUT83), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n316), .A2(KEYINPUT16), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(G146), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n316), .B(KEYINPUT19), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n191), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT83), .B1(new_n321), .B2(new_n322), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n320), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G113), .B(G122), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(new_n205), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n333), .B(KEYINPUT84), .Z(new_n336));
  AND3_X1   g150(.A1(new_n324), .A2(G146), .A3(new_n325), .ZN(new_n337));
  AOI21_X1  g151(.A(G146), .B1(new_n324), .B2(new_n325), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT17), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n321), .A2(new_n340), .A3(new_n322), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n339), .B(new_n341), .C1(new_n340), .C2(new_n322), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n342), .A3(new_n320), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(G475), .A2(G902), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT20), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n348), .A3(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G234), .ZN(new_n351));
  INV_X1    g165(.A(G237), .ZN(new_n352));
  AND2_X1   g166(.A1(KEYINPUT87), .A2(G952), .ZN(new_n353));
  NOR2_X1   g167(.A1(KEYINPUT87), .A2(G952), .ZN(new_n354));
  OAI221_X1 g168(.A(new_n273), .B1(new_n351), .B2(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT21), .B(G898), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT88), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI211_X1 g173(.A(new_n293), .B(new_n273), .C1(G234), .C2(G237), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n356), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G217), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n187), .A2(new_n363), .A3(G953), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(G116), .B(G122), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT85), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n366), .A2(new_n367), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n207), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(G128), .B(G143), .Z(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(G134), .ZN(new_n373));
  INV_X1    g187(.A(G116), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT14), .A3(G122), .ZN(new_n375));
  XOR2_X1   g189(.A(G116), .B(G122), .Z(new_n376));
  OAI211_X1 g190(.A(G107), .B(new_n375), .C1(new_n376), .C2(KEYINPUT14), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n371), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(KEYINPUT85), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n368), .A3(G107), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n193), .A2(G128), .B1(KEYINPUT86), .B2(KEYINPUT13), .ZN(new_n381));
  AND2_X1   g195(.A1(KEYINPUT86), .A2(KEYINPUT13), .ZN(new_n382));
  OAI21_X1  g196(.A(G134), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n383), .A2(new_n372), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n372), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n371), .A2(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n365), .B1(new_n378), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n371), .A2(new_n380), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n385), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n371), .A2(new_n373), .A3(new_n377), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(new_n364), .ZN(new_n392));
  AOI21_X1  g206(.A(G902), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G478), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT15), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n393), .B(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n343), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n333), .B1(new_n342), .B2(new_n320), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n293), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G475), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n350), .A2(new_n362), .A3(new_n396), .A4(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G210), .B1(G237), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G119), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G116), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n374), .A2(G119), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT2), .B(G113), .Z(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n406), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT2), .B(G113), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n251), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT5), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G113), .B1(new_n405), .B2(KEYINPUT5), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n419), .A2(new_n409), .A3(new_n214), .A4(new_n217), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G122), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n414), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n200), .A2(new_n312), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n198), .A3(new_n202), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT78), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n423), .A2(new_n198), .A3(KEYINPUT78), .A4(new_n202), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT79), .B(G224), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n273), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT7), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n260), .B2(G125), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n409), .B1(new_n415), .B2(new_n417), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n218), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n420), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n421), .B(KEYINPUT8), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n426), .A2(new_n427), .B1(G125), .B2(new_n260), .ZN(new_n439));
  INV_X1    g253(.A(new_n431), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n433), .B(new_n438), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n422), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n260), .A2(G125), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n428), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n431), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n428), .A2(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT80), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(KEYINPUT81), .B(new_n293), .C1(new_n443), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n414), .A2(new_n420), .ZN(new_n450));
  INV_X1    g264(.A(new_n421), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT6), .A3(new_n422), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n439), .B(new_n430), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(new_n455), .A3(new_n451), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n449), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n441), .A2(new_n442), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n446), .A2(KEYINPUT80), .A3(new_n447), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n422), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT81), .B1(new_n461), .B2(new_n293), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n403), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n293), .B1(new_n443), .B2(new_n448), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT81), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n466), .A2(new_n402), .A3(new_n457), .A4(new_n449), .ZN(new_n467));
  AOI211_X1 g281(.A(new_n301), .B(new_n401), .C1(new_n463), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n233), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n198), .A2(new_n200), .A3(new_n202), .ZN(new_n470));
  AOI21_X1  g284(.A(G134), .B1(new_n229), .B2(new_n231), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n226), .A2(G137), .ZN(new_n472));
  OAI21_X1  g286(.A(G131), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n475));
  OAI22_X1  g289(.A1(new_n262), .A2(new_n475), .B1(new_n233), .B2(new_n234), .ZN(new_n476));
  AOI211_X1 g290(.A(KEYINPUT65), .B(new_n258), .C1(new_n254), .C2(new_n255), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT30), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n261), .A2(new_n235), .A3(new_n264), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(KEYINPUT30), .A3(new_n474), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n482), .A3(new_n413), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n413), .B(KEYINPUT69), .Z(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n484), .A3(new_n474), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n302), .A2(G210), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT27), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT26), .B(G101), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n483), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT31), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n483), .A2(KEYINPUT31), .A3(new_n485), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT28), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n485), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n478), .A2(new_n413), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n497), .A2(new_n485), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n496), .B1(new_n498), .B2(new_n495), .ZN(new_n499));
  INV_X1    g313(.A(new_n489), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(G472), .A2(G902), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(KEYINPUT32), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n492), .A2(new_n493), .B1(new_n499), .B2(new_n500), .ZN(new_n506));
  INV_X1    g320(.A(new_n503), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n495), .B1(new_n497), .B2(new_n485), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n282), .B2(new_n235), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT28), .B1(new_n511), .B2(new_n484), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n509), .A2(new_n512), .A3(new_n500), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n489), .B1(new_n483), .B2(new_n485), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n513), .A2(KEYINPUT29), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n481), .A2(new_n474), .ZN(new_n516));
  INV_X1    g330(.A(new_n484), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n485), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT28), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT29), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n500), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n496), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n293), .ZN(new_n524));
  OAI21_X1  g338(.A(G472), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n504), .A2(new_n508), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n363), .B1(G234), .B2(new_n293), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n404), .B2(G128), .ZN(new_n531));
  INV_X1    g345(.A(G128), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT23), .A3(G119), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n531), .B(new_n533), .C1(G119), .C2(new_n532), .ZN(new_n534));
  XNOR2_X1  g348(.A(G119), .B(G128), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT24), .B(G110), .Z(new_n536));
  AOI22_X1  g350(.A1(new_n534), .A2(G110), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n337), .B2(new_n338), .ZN(new_n538));
  OAI22_X1  g352(.A1(new_n534), .A2(G110), .B1(new_n535), .B2(new_n536), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n318), .A3(new_n326), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT22), .B(G137), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n538), .A2(new_n540), .A3(new_n544), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n293), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n546), .A2(KEYINPUT25), .A3(new_n293), .A4(new_n547), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n529), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n528), .A2(G902), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(new_n547), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n526), .A2(new_n527), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n527), .B1(new_n526), .B2(new_n557), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n299), .B(new_n468), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT89), .B(G101), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(G3));
  INV_X1    g376(.A(KEYINPUT91), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n463), .A2(new_n563), .A3(new_n467), .ZN(new_n564));
  INV_X1    g378(.A(new_n301), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n458), .A2(new_n462), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(KEYINPUT91), .A3(new_n402), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n350), .A2(new_n400), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n378), .A2(new_n386), .A3(new_n365), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n364), .B1(new_n390), .B2(new_n391), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n293), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(new_n394), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT93), .B1(new_n393), .B2(G478), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n394), .A2(G902), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT33), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n579), .B(new_n580), .C1(new_n387), .C2(new_n392), .ZN(new_n581));
  AND4_X1   g395(.A1(KEYINPUT92), .A2(new_n387), .A3(new_n392), .A4(new_n578), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n577), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n576), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n576), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n569), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n362), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(KEYINPUT90), .A2(G472), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n502), .A2(new_n293), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n591), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n506), .B2(G902), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n556), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n568), .A2(new_n299), .A3(new_n590), .A4(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT34), .B(G104), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G6));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n600));
  INV_X1    g414(.A(new_n569), .ZN(new_n601));
  INV_X1    g415(.A(new_n396), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n361), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n568), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n606));
  INV_X1    g420(.A(new_n603), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n362), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT95), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n299), .A3(new_n596), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G107), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n545), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n541), .B(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n616), .A2(new_n554), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n552), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n614), .B1(new_n595), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n618), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n592), .A2(new_n594), .A3(KEYINPUT96), .A4(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n619), .A2(new_n468), .A3(new_n299), .A4(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT37), .B(G110), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT97), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n622), .B(new_n624), .ZN(G12));
  NAND2_X1  g439(.A1(new_n526), .A2(new_n620), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n606), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n360), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n355), .B1(new_n628), .B2(G900), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT98), .Z(new_n630));
  NOR2_X1   g444(.A1(new_n603), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n299), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G128), .ZN(G30));
  NOR2_X1   g448(.A1(new_n601), .A2(new_n396), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n565), .A3(new_n618), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(KEYINPUT100), .Z(new_n637));
  NAND2_X1  g451(.A1(new_n463), .A2(new_n467), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT38), .Z(new_n639));
  NOR2_X1   g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n630), .B(KEYINPUT39), .Z(new_n641));
  NAND2_X1  g455(.A1(new_n299), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT40), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n293), .B1(new_n519), .B2(new_n489), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n500), .B1(new_n483), .B2(new_n485), .ZN(new_n645));
  OAI21_X1  g459(.A(G472), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n504), .A2(new_n508), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT99), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n642), .A2(KEYINPUT40), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n640), .A2(new_n643), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G143), .ZN(G45));
  INV_X1    g465(.A(G472), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n496), .B(new_n489), .C1(new_n498), .C2(new_n495), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n483), .A2(new_n485), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n500), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n655), .A3(new_n521), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n512), .B1(new_n519), .B2(KEYINPUT28), .ZN(new_n657));
  AOI21_X1  g471(.A(G902), .B1(new_n657), .B2(new_n522), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n652), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n502), .A2(new_n503), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n659), .B1(new_n660), .B2(new_n505), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n618), .B1(new_n661), .B2(new_n504), .ZN(new_n662));
  INV_X1    g476(.A(new_n630), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n569), .B(new_n663), .C1(new_n585), .C2(new_n586), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n568), .A2(new_n662), .A3(new_n299), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G146), .ZN(G48));
  AND3_X1   g481(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n668), .A2(new_n669), .A3(new_n189), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n556), .B1(new_n661), .B2(new_n504), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n568), .A2(new_n670), .A3(new_n671), .A4(new_n590), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NAND2_X1  g488(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n605), .B2(new_n609), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT101), .B(G116), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G18));
  INV_X1    g492(.A(new_n401), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n568), .A2(new_n670), .A3(new_n679), .A4(new_n662), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  NAND4_X1  g495(.A1(new_n564), .A2(new_n567), .A3(new_n565), .A4(new_n635), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n189), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n271), .A2(new_n288), .A3(new_n276), .A4(new_n289), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n270), .A2(new_n276), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n268), .A2(new_n269), .B1(new_n235), .B2(new_n278), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n271), .B1(new_n687), .B2(new_n276), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n685), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(G469), .B1(new_n689), .B2(G902), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n684), .A2(new_n690), .A3(new_n294), .A4(new_n362), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n494), .B1(new_n489), .B2(new_n657), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n503), .B(KEYINPUT102), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n506), .B2(G902), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n556), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n683), .A2(new_n691), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  NOR3_X1   g513(.A1(new_n696), .A2(new_n618), .A3(new_n664), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n568), .A2(new_n670), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  NAND3_X1  g516(.A1(new_n463), .A2(new_n565), .A3(new_n467), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT103), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n463), .A2(new_n467), .A3(new_n705), .A4(new_n565), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n299), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n671), .A3(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n299), .A2(new_n704), .A3(new_n665), .A4(new_n706), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n506), .A2(new_n505), .A3(new_n507), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n508), .B(new_n525), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n504), .A2(KEYINPUT104), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n557), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT42), .B1(new_n710), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n709), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n228), .ZN(G33));
  NAND4_X1  g532(.A1(new_n671), .A2(new_n299), .A3(new_n706), .A4(new_n704), .ZN(new_n719));
  INV_X1    g533(.A(new_n631), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT105), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n707), .A2(new_n722), .A3(new_n671), .A4(new_n631), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  AND2_X1   g539(.A1(new_n704), .A2(new_n706), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n585), .A2(new_n586), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n601), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(KEYINPUT43), .Z(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n595), .A3(new_n620), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n732), .B2(new_n731), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n734), .A2(KEYINPUT106), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(KEYINPUT106), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n295), .B1(new_n276), .B2(new_n270), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(G469), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n297), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n668), .B1(new_n742), .B2(new_n743), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n189), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(new_n641), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n735), .A2(new_n736), .A3(new_n748), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT107), .B(G137), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G39));
  OR2_X1    g565(.A1(new_n747), .A2(KEYINPUT47), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n747), .A2(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n727), .A2(new_n526), .A3(new_n557), .A4(new_n664), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(KEYINPUT108), .B(G140), .Z(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G42));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n730), .A2(new_n356), .A3(new_n697), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(new_n301), .A3(new_n639), .A4(new_n670), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n690), .A2(new_n684), .A3(new_n294), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n727), .A2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n767), .A2(new_n356), .A3(new_n730), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n620), .A3(new_n695), .A4(new_n694), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n761), .A2(new_n762), .A3(KEYINPUT50), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n648), .A2(new_n556), .A3(new_n355), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(new_n767), .ZN(new_n772));
  INV_X1    g586(.A(new_n728), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n601), .A3(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n765), .A2(new_n769), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n760), .A2(new_n726), .ZN(new_n776));
  INV_X1    g590(.A(new_n754), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n668), .A2(new_n669), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n189), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT113), .Z(new_n780));
  AOI21_X1  g594(.A(new_n776), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n759), .B1(new_n775), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT115), .ZN(new_n783));
  INV_X1    g597(.A(new_n715), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n768), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(KEYINPUT48), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n772), .A2(new_n588), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n273), .B1(new_n353), .B2(new_n354), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n606), .A2(new_n766), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n789), .B1(new_n760), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n786), .A2(KEYINPUT48), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n787), .A2(new_n788), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n775), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n777), .A2(new_n779), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n776), .B1(new_n796), .B2(KEYINPUT117), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n759), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n793), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n783), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n569), .A2(new_n602), .A3(new_n630), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n526), .A2(new_n620), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n665), .A2(new_n695), .A3(new_n620), .A4(new_n694), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n707), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n301), .B1(new_n463), .B2(new_n467), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n361), .B1(new_n603), .B2(new_n587), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n596), .A2(new_n299), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n622), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n294), .A2(new_n298), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n807), .A3(new_n684), .A4(new_n679), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n526), .A2(new_n557), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT71), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n526), .A2(new_n527), .A3(new_n557), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n724), .A2(new_n806), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n299), .A2(new_n704), .A3(new_n706), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n804), .B2(new_n803), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n810), .A3(new_n816), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(KEYINPUT112), .A3(new_n724), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n698), .A2(new_n672), .A3(new_n680), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n717), .A2(new_n826), .A3(new_n676), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT109), .B1(new_n618), .B2(new_n663), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT109), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n552), .A2(new_n617), .A3(new_n829), .A4(new_n630), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n189), .B(new_n831), .C1(new_n294), .C2(new_n298), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n683), .A2(KEYINPUT110), .A3(new_n647), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  INV_X1    g648(.A(new_n831), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n811), .A2(new_n684), .A3(new_n647), .A4(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n834), .B1(new_n836), .B2(new_n682), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n633), .A2(new_n666), .A3(new_n701), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT52), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n833), .A2(new_n837), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n627), .A2(new_n632), .B1(new_n790), .B2(new_n700), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n666), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n633), .A2(new_n701), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(new_n846), .B2(KEYINPUT52), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n827), .A2(new_n840), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n825), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n840), .A2(new_n844), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n826), .A2(new_n676), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n709), .A2(new_n716), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n823), .A3(new_n852), .A4(new_n724), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n845), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT111), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT111), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n856), .B(new_n845), .C1(new_n850), .C2(new_n853), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n849), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n806), .A2(new_n560), .A3(new_n622), .A4(new_n809), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n723), .B2(new_n721), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n827), .A3(new_n844), .A4(new_n840), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n846), .A2(KEYINPUT52), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n845), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n845), .B2(new_n863), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n860), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n801), .A2(new_n867), .B1(G952), .B2(G953), .ZN(new_n868));
  OR4_X1    g682(.A1(new_n556), .A2(new_n729), .A3(new_n189), .A4(new_n301), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n778), .B(KEYINPUT49), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n639), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n868), .B1(new_n648), .B2(new_n872), .ZN(G75));
  OAI21_X1  g687(.A(KEYINPUT119), .B1(new_n858), .B2(new_n293), .ZN(new_n874));
  INV_X1    g688(.A(new_n850), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n827), .A2(new_n847), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n820), .A4(new_n824), .ZN(new_n877));
  INV_X1    g691(.A(new_n857), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n856), .B1(new_n863), .B2(new_n845), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n881), .A3(G902), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n874), .A2(new_n882), .A3(new_n403), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n874), .A2(new_n882), .A3(KEYINPUT120), .A4(new_n403), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n453), .A2(new_n456), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(new_n454), .Z(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(KEYINPUT56), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n885), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n273), .A2(G952), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n880), .A2(G210), .A3(G902), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT118), .B1(new_n896), .B2(new_n889), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n898));
  INV_X1    g712(.A(new_n889), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n898), .B(new_n899), .C1(new_n894), .C2(new_n895), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n893), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n891), .A2(new_n901), .ZN(G51));
  NAND2_X1  g716(.A1(new_n880), .A2(KEYINPUT54), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n860), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n297), .B(KEYINPUT57), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n291), .B(KEYINPUT121), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n741), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n874), .A2(new_n882), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n892), .B1(new_n908), .B2(new_n910), .ZN(G54));
  NAND4_X1  g725(.A1(new_n874), .A2(new_n882), .A3(KEYINPUT58), .A4(G475), .ZN(new_n912));
  INV_X1    g726(.A(new_n344), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n892), .ZN(G60));
  OR2_X1    g730(.A1(new_n581), .A2(new_n582), .ZN(new_n917));
  XNOR2_X1  g731(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n904), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n917), .B1(new_n867), .B2(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n892), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT60), .Z(new_n925));
  NAND2_X1  g739(.A1(new_n880), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n616), .B(KEYINPUT123), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n893), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT61), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n546), .A2(new_n547), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n932), .B(new_n893), .C1(new_n926), .C2(new_n927), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n930), .B(new_n933), .ZN(G66));
  INV_X1    g748(.A(new_n429), .ZN(new_n935));
  OAI21_X1  g749(.A(G953), .B1(new_n359), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n851), .A2(new_n817), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n938), .B2(G953), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT125), .Z(new_n940));
  OAI21_X1  g754(.A(new_n887), .B1(G898), .B2(new_n273), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G69));
  NAND2_X1  g756(.A1(new_n480), .A2(new_n482), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT126), .Z(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n327), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n558), .A2(new_n559), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n607), .A2(new_n588), .ZN(new_n947));
  NOR4_X1   g761(.A1(new_n727), .A2(new_n946), .A3(new_n642), .A4(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n754), .B2(new_n755), .ZN(new_n949));
  INV_X1    g763(.A(new_n839), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n650), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n749), .A2(new_n949), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n945), .B1(new_n954), .B2(new_n273), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n749), .A2(new_n852), .A3(new_n724), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n748), .A2(new_n683), .A3(new_n784), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n756), .A2(new_n950), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n273), .ZN(new_n960));
  INV_X1    g774(.A(new_n945), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(G900), .B2(G953), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n955), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n273), .B1(G227), .B2(G900), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n963), .B(new_n964), .Z(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n954), .B2(new_n937), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n645), .ZN(new_n969));
  INV_X1    g783(.A(new_n967), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n655), .A2(new_n490), .ZN(new_n971));
  OR3_X1    g785(.A1(new_n866), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n969), .A2(new_n972), .A3(new_n893), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n959), .B2(new_n938), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT127), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n654), .A2(new_n489), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G57));
endmodule


