

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747;

  OR2_X1 U373 ( .A1(n538), .A2(n515), .ZN(n524) );
  XNOR2_X1 U374 ( .A(n386), .B(n560), .ZN(n385) );
  NAND2_X1 U375 ( .A1(n385), .A2(n566), .ZN(n384) );
  NAND2_X1 U376 ( .A1(n596), .A2(n582), .ZN(n583) );
  XNOR2_X2 U377 ( .A(n576), .B(n577), .ZN(n596) );
  NOR2_X2 U378 ( .A1(n745), .A2(n365), .ZN(n591) );
  XNOR2_X1 U379 ( .A(n553), .B(KEYINPUT42), .ZN(n747) );
  NAND2_X2 U380 ( .A1(n678), .A2(n676), .ZN(n551) );
  NAND2_X2 U381 ( .A1(n694), .A2(n615), .ZN(n363) );
  XOR2_X2 U382 ( .A(n707), .B(KEYINPUT59), .Z(n708) );
  XNOR2_X2 U383 ( .A(n446), .B(n445), .ZN(n449) );
  XNOR2_X2 U384 ( .A(n447), .B(G101), .ZN(n448) );
  XNOR2_X2 U385 ( .A(n459), .B(n458), .ZN(n720) );
  XNOR2_X2 U386 ( .A(n449), .B(n448), .ZN(n459) );
  OR2_X1 U387 ( .A1(n570), .A2(n552), .ZN(n537) );
  NAND2_X2 U388 ( .A1(n587), .A2(n586), .ZN(n366) );
  XNOR2_X2 U389 ( .A(n524), .B(n523), .ZN(n570) );
  NOR2_X1 U390 ( .A1(n520), .A2(n656), .ZN(n544) );
  NAND2_X1 U391 ( .A1(n656), .A2(KEYINPUT70), .ZN(n377) );
  INV_X1 U392 ( .A(n592), .ZN(n513) );
  AND2_X1 U393 ( .A1(n573), .A2(n687), .ZN(n574) );
  XNOR2_X1 U394 ( .A(n367), .B(KEYINPUT35), .ZN(n745) );
  BUF_X1 U395 ( .A(n578), .Z(n660) );
  XNOR2_X1 U396 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n439) );
  XNOR2_X1 U397 ( .A(KEYINPUT66), .B(G131), .ZN(n482) );
  XNOR2_X1 U398 ( .A(n388), .B(KEYINPUT81), .ZN(n351) );
  XNOR2_X1 U399 ( .A(n388), .B(KEYINPUT81), .ZN(n611) );
  NAND2_X1 U400 ( .A1(n385), .A2(n566), .ZN(n352) );
  NOR2_X1 U401 ( .A1(n383), .A2(n351), .ZN(n353) );
  BUF_X1 U402 ( .A(n678), .Z(n354) );
  NOR2_X1 U403 ( .A1(n383), .A2(n611), .ZN(n382) );
  BUF_X1 U404 ( .A(n747), .Z(n355) );
  BUF_X1 U405 ( .A(n459), .Z(n356) );
  XNOR2_X1 U406 ( .A(n352), .B(n390), .ZN(n357) );
  XNOR2_X1 U407 ( .A(n384), .B(n390), .ZN(n389) );
  XNOR2_X2 U408 ( .A(G119), .B(G116), .ZN(n446) );
  XNOR2_X2 U409 ( .A(n538), .B(KEYINPUT38), .ZN(n546) );
  INV_X1 U410 ( .A(KEYINPUT33), .ZN(n378) );
  NAND2_X1 U411 ( .A1(n371), .A2(n370), .ZN(n379) );
  NOR2_X1 U412 ( .A1(n373), .A2(n372), .ZN(n371) );
  NAND2_X1 U413 ( .A1(n375), .A2(n374), .ZN(n370) );
  NOR2_X1 U414 ( .A1(n655), .A2(KEYINPUT70), .ZN(n374) );
  XNOR2_X1 U415 ( .A(n387), .B(KEYINPUT80), .ZN(n383) );
  XNOR2_X1 U416 ( .A(G134), .B(KEYINPUT7), .ZN(n495) );
  XNOR2_X1 U417 ( .A(n483), .B(KEYINPUT12), .ZN(n484) );
  XNOR2_X1 U418 ( .A(G113), .B(G143), .ZN(n481) );
  XNOR2_X1 U419 ( .A(n514), .B(KEYINPUT101), .ZN(n562) );
  NAND2_X1 U420 ( .A1(n513), .A2(n395), .ZN(n514) );
  XNOR2_X1 U421 ( .A(n492), .B(n391), .ZN(n549) );
  OR2_X1 U422 ( .A1(n707), .A2(G902), .ZN(n492) );
  OR2_X1 U423 ( .A1(n702), .A2(G902), .ZN(n405) );
  INV_X1 U424 ( .A(KEYINPUT67), .ZN(n445) );
  NAND2_X1 U425 ( .A1(n376), .A2(n513), .ZN(n372) );
  XNOR2_X1 U426 ( .A(G137), .B(KEYINPUT95), .ZN(n440) );
  XOR2_X1 U427 ( .A(KEYINPUT96), .B(G122), .Z(n494) );
  XOR2_X1 U428 ( .A(KEYINPUT97), .B(KEYINPUT9), .Z(n496) );
  XNOR2_X1 U429 ( .A(n461), .B(KEYINPUT10), .ZN(n476) );
  XOR2_X1 U430 ( .A(KEYINPUT17), .B(KEYINPUT74), .Z(n462) );
  INV_X1 U431 ( .A(KEYINPUT82), .ZN(n390) );
  AND2_X1 U432 ( .A1(n588), .A2(n674), .ZN(n455) );
  INV_X1 U433 ( .A(G237), .ZN(n454) );
  XNOR2_X1 U434 ( .A(n425), .B(n424), .ZN(n578) );
  NOR2_X1 U435 ( .A1(n716), .A2(G902), .ZN(n425) );
  XNOR2_X1 U436 ( .A(n486), .B(KEYINPUT16), .ZN(n458) );
  XNOR2_X1 U437 ( .A(KEYINPUT77), .B(KEYINPUT24), .ZN(n408) );
  XNOR2_X1 U438 ( .A(G119), .B(G128), .ZN(n406) );
  XNOR2_X1 U439 ( .A(G140), .B(G137), .ZN(n417) );
  INV_X1 U440 ( .A(G953), .ZN(n726) );
  NAND2_X1 U441 ( .A1(n361), .A2(n370), .ZN(n597) );
  AND2_X1 U442 ( .A1(n676), .A2(n661), .ZN(n582) );
  INV_X1 U443 ( .A(KEYINPUT64), .ZN(n399) );
  XNOR2_X1 U444 ( .A(n383), .B(n741), .ZN(n742) );
  XNOR2_X1 U445 ( .A(n380), .B(G107), .ZN(n397) );
  INV_X1 U446 ( .A(G110), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n505), .B(n504), .ZN(n712) );
  XNOR2_X1 U448 ( .A(n503), .B(KEYINPUT98), .ZN(n504) );
  XNOR2_X1 U449 ( .A(n491), .B(n490), .ZN(n707) );
  XNOR2_X1 U450 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U451 ( .A(n485), .B(n484), .ZN(n491) );
  OR2_X1 U452 ( .A1(n411), .A2(G952), .ZN(n699) );
  XNOR2_X1 U453 ( .A(n556), .B(n555), .ZN(n623) );
  XNOR2_X1 U454 ( .A(n519), .B(n393), .ZN(n520) );
  NAND2_X1 U455 ( .A1(n369), .A2(n368), .ZN(n367) );
  INV_X1 U456 ( .A(n581), .ZN(n368) );
  XNOR2_X1 U457 ( .A(n379), .B(n378), .ZN(n652) );
  INV_X1 U458 ( .A(n656), .ZN(n375) );
  XNOR2_X1 U459 ( .A(KEYINPUT75), .B(n569), .ZN(n358) );
  XOR2_X1 U460 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n359) );
  OR2_X1 U461 ( .A1(G953), .A2(G237), .ZN(n360) );
  XNOR2_X1 U462 ( .A(n588), .B(n510), .ZN(n592) );
  AND2_X1 U463 ( .A1(n377), .A2(n376), .ZN(n361) );
  AND2_X2 U464 ( .A1(n608), .A2(n607), .ZN(n381) );
  NOR2_X1 U465 ( .A1(n624), .A2(n610), .ZN(n473) );
  INV_X1 U466 ( .A(n595), .ZN(n587) );
  NAND2_X1 U467 ( .A1(n382), .A2(n362), .ZN(n364) );
  AND2_X2 U468 ( .A1(n725), .A2(n610), .ZN(n362) );
  NAND2_X2 U469 ( .A1(n364), .A2(n363), .ZN(n706) );
  NAND2_X1 U470 ( .A1(n351), .A2(n725), .ZN(n694) );
  XNOR2_X2 U471 ( .A(n381), .B(n609), .ZN(n725) );
  NAND2_X1 U472 ( .A1(n746), .A2(n640), .ZN(n365) );
  XNOR2_X2 U473 ( .A(n366), .B(KEYINPUT32), .ZN(n746) );
  XNOR2_X1 U474 ( .A(n580), .B(KEYINPUT34), .ZN(n369) );
  INV_X1 U475 ( .A(n377), .ZN(n373) );
  NAND2_X1 U476 ( .A1(n655), .A2(KEYINPUT70), .ZN(n376) );
  NAND2_X1 U477 ( .A1(n353), .A2(n725), .ZN(n693) );
  NAND2_X1 U478 ( .A1(n558), .A2(n559), .ZN(n386) );
  NAND2_X1 U479 ( .A1(n357), .A2(n568), .ZN(n387) );
  NAND2_X1 U480 ( .A1(n389), .A2(n358), .ZN(n388) );
  NOR2_X2 U481 ( .A1(n747), .A2(n623), .ZN(n557) );
  XNOR2_X2 U482 ( .A(n547), .B(KEYINPUT103), .ZN(n678) );
  NOR2_X2 U483 ( .A1(n673), .A2(n552), .ZN(n553) );
  XNOR2_X2 U484 ( .A(n551), .B(n550), .ZN(n673) );
  XOR2_X1 U485 ( .A(KEYINPUT13), .B(G475), .Z(n391) );
  XOR2_X1 U486 ( .A(KEYINPUT69), .B(KEYINPUT39), .Z(n392) );
  XOR2_X1 U487 ( .A(n518), .B(KEYINPUT36), .Z(n393) );
  AND2_X1 U488 ( .A1(n578), .A2(n435), .ZN(n394) );
  AND2_X1 U489 ( .A1(n646), .A2(n525), .ZN(n395) );
  INV_X1 U490 ( .A(KEYINPUT48), .ZN(n560) );
  XNOR2_X1 U491 ( .A(n734), .B(G146), .ZN(n451) );
  XNOR2_X2 U492 ( .A(G143), .B(G128), .ZN(n502) );
  XNOR2_X1 U493 ( .A(n502), .B(KEYINPUT4), .ZN(n463) );
  INV_X1 U494 ( .A(G134), .ZN(n509) );
  XNOR2_X1 U495 ( .A(n482), .B(n509), .ZN(n396) );
  XNOR2_X1 U496 ( .A(n463), .B(n396), .ZN(n734) );
  XNOR2_X1 U497 ( .A(n397), .B(KEYINPUT85), .ZN(n721) );
  XNOR2_X1 U498 ( .A(n721), .B(KEYINPUT68), .ZN(n460) );
  XNOR2_X1 U499 ( .A(G104), .B(G101), .ZN(n398) );
  XNOR2_X1 U500 ( .A(n417), .B(n398), .ZN(n401) );
  XNOR2_X2 U501 ( .A(n399), .B(G953), .ZN(n411) );
  NAND2_X1 U502 ( .A1(n411), .A2(G227), .ZN(n400) );
  XNOR2_X1 U503 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U504 ( .A(n460), .B(n402), .ZN(n403) );
  XNOR2_X1 U505 ( .A(n451), .B(n403), .ZN(n702) );
  INV_X1 U506 ( .A(G469), .ZN(n404) );
  XNOR2_X2 U507 ( .A(n405), .B(n404), .ZN(n599) );
  INV_X1 U508 ( .A(n599), .ZN(n436) );
  XOR2_X1 U509 ( .A(KEYINPUT86), .B(G110), .Z(n407) );
  XNOR2_X1 U510 ( .A(n407), .B(n406), .ZN(n410) );
  XNOR2_X1 U511 ( .A(n359), .B(n408), .ZN(n409) );
  XOR2_X1 U512 ( .A(n410), .B(n409), .Z(n416) );
  NAND2_X1 U513 ( .A1(G234), .A2(n411), .ZN(n414) );
  XNOR2_X1 U514 ( .A(KEYINPUT8), .B(KEYINPUT65), .ZN(n412) );
  XNOR2_X1 U515 ( .A(n412), .B(KEYINPUT78), .ZN(n413) );
  XNOR2_X1 U516 ( .A(n414), .B(n413), .ZN(n499) );
  NAND2_X1 U517 ( .A1(G221), .A2(n499), .ZN(n415) );
  XNOR2_X1 U518 ( .A(n416), .B(n415), .ZN(n419) );
  XNOR2_X2 U519 ( .A(G146), .B(G125), .ZN(n461) );
  INV_X1 U520 ( .A(n417), .ZN(n418) );
  XNOR2_X1 U521 ( .A(n476), .B(n418), .ZN(n736) );
  XNOR2_X1 U522 ( .A(n419), .B(n736), .ZN(n716) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(KEYINPUT89), .Z(n423) );
  XNOR2_X1 U524 ( .A(G902), .B(KEYINPUT15), .ZN(n612) );
  NAND2_X1 U525 ( .A1(n612), .A2(G234), .ZN(n421) );
  XNOR2_X1 U526 ( .A(KEYINPUT88), .B(KEYINPUT20), .ZN(n420) );
  XNOR2_X1 U527 ( .A(n421), .B(n420), .ZN(n426) );
  NAND2_X1 U528 ( .A1(G217), .A2(n426), .ZN(n422) );
  XNOR2_X1 U529 ( .A(n423), .B(n422), .ZN(n424) );
  NAND2_X1 U530 ( .A1(G221), .A2(n426), .ZN(n428) );
  XOR2_X1 U531 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n427) );
  XNOR2_X1 U532 ( .A(n428), .B(n427), .ZN(n661) );
  NAND2_X1 U533 ( .A1(G237), .A2(G234), .ZN(n429) );
  XNOR2_X1 U534 ( .A(n429), .B(KEYINPUT14), .ZN(n687) );
  AND2_X1 U535 ( .A1(n661), .A2(n687), .ZN(n434) );
  INV_X1 U536 ( .A(G900), .ZN(n430) );
  NAND2_X1 U537 ( .A1(n430), .A2(G902), .ZN(n431) );
  OR2_X1 U538 ( .A1(n411), .A2(n431), .ZN(n432) );
  NAND2_X1 U539 ( .A1(n726), .A2(G952), .ZN(n571) );
  NAND2_X1 U540 ( .A1(n432), .A2(n571), .ZN(n433) );
  NAND2_X1 U541 ( .A1(n434), .A2(n433), .ZN(n512) );
  INV_X1 U542 ( .A(n512), .ZN(n435) );
  NAND2_X1 U543 ( .A1(n436), .A2(n394), .ZN(n438) );
  INV_X1 U544 ( .A(KEYINPUT72), .ZN(n437) );
  XNOR2_X1 U545 ( .A(n438), .B(n437), .ZN(n457) );
  XNOR2_X1 U546 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U547 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n441) );
  XNOR2_X1 U548 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U549 ( .A(n360), .B(KEYINPUT71), .ZN(n487) );
  NAND2_X1 U550 ( .A1(n487), .A2(G210), .ZN(n443) );
  XNOR2_X1 U551 ( .A(n444), .B(n443), .ZN(n450) );
  XNOR2_X2 U552 ( .A(G113), .B(KEYINPUT3), .ZN(n447) );
  XNOR2_X1 U553 ( .A(n450), .B(n356), .ZN(n452) );
  XNOR2_X1 U554 ( .A(n452), .B(n451), .ZN(n617) );
  OR2_X2 U555 ( .A1(n617), .A2(G902), .ZN(n453) );
  XNOR2_X2 U556 ( .A(n453), .B(G472), .ZN(n588) );
  INV_X1 U557 ( .A(G902), .ZN(n506) );
  NAND2_X1 U558 ( .A1(n506), .A2(n454), .ZN(n471) );
  NAND2_X1 U559 ( .A1(n471), .A2(G214), .ZN(n674) );
  XNOR2_X1 U560 ( .A(n455), .B(KEYINPUT30), .ZN(n456) );
  NAND2_X1 U561 ( .A1(n457), .A2(n456), .ZN(n539) );
  INV_X1 U562 ( .A(n539), .ZN(n474) );
  XOR2_X1 U563 ( .A(G104), .B(G122), .Z(n486) );
  XNOR2_X1 U564 ( .A(n720), .B(n460), .ZN(n470) );
  XNOR2_X1 U565 ( .A(n462), .B(n461), .ZN(n464) );
  XOR2_X1 U566 ( .A(n464), .B(n463), .Z(n468) );
  XOR2_X1 U567 ( .A(KEYINPUT18), .B(KEYINPUT73), .Z(n466) );
  NAND2_X1 U568 ( .A1(G224), .A2(n411), .ZN(n465) );
  XNOR2_X1 U569 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U570 ( .A(n468), .B(n467), .Z(n469) );
  XNOR2_X1 U571 ( .A(n470), .B(n469), .ZN(n624) );
  INV_X1 U572 ( .A(n612), .ZN(n610) );
  AND2_X1 U573 ( .A1(n471), .A2(G210), .ZN(n472) );
  XNOR2_X2 U574 ( .A(n473), .B(n472), .ZN(n538) );
  NAND2_X1 U575 ( .A1(n474), .A2(n546), .ZN(n475) );
  XNOR2_X2 U576 ( .A(n475), .B(n392), .ZN(n554) );
  NAND2_X1 U577 ( .A1(n476), .A2(G140), .ZN(n480) );
  INV_X1 U578 ( .A(n476), .ZN(n478) );
  INV_X1 U579 ( .A(G140), .ZN(n477) );
  NAND2_X1 U580 ( .A1(n478), .A2(n477), .ZN(n479) );
  NAND2_X1 U581 ( .A1(n480), .A2(n479), .ZN(n485) );
  XNOR2_X1 U582 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U583 ( .A(n486), .B(KEYINPUT11), .ZN(n489) );
  NAND2_X1 U584 ( .A1(G214), .A2(n487), .ZN(n488) );
  XNOR2_X1 U585 ( .A(G116), .B(G107), .ZN(n493) );
  XNOR2_X1 U586 ( .A(n494), .B(n493), .ZN(n498) );
  XNOR2_X1 U587 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U588 ( .A(n498), .B(n497), .Z(n501) );
  NAND2_X1 U589 ( .A1(n499), .A2(G217), .ZN(n500) );
  XNOR2_X1 U590 ( .A(n501), .B(n500), .ZN(n505) );
  INV_X1 U591 ( .A(n502), .ZN(n503) );
  NAND2_X1 U592 ( .A1(n712), .A2(n506), .ZN(n507) );
  XNOR2_X1 U593 ( .A(n507), .B(G478), .ZN(n548) );
  INV_X1 U594 ( .A(n548), .ZN(n511) );
  OR2_X1 U595 ( .A1(n549), .A2(n511), .ZN(n508) );
  XNOR2_X1 U596 ( .A(n508), .B(KEYINPUT99), .ZN(n648) );
  AND2_X1 U597 ( .A1(n554), .A2(n648), .ZN(n567) );
  XNOR2_X1 U598 ( .A(n567), .B(n509), .ZN(G36) );
  XNOR2_X1 U599 ( .A(KEYINPUT100), .B(KEYINPUT6), .ZN(n510) );
  AND2_X2 U600 ( .A1(n549), .A2(n511), .ZN(n646) );
  NOR2_X1 U601 ( .A1(n578), .A2(n512), .ZN(n525) );
  XNOR2_X1 U602 ( .A(n562), .B(KEYINPUT104), .ZN(n517) );
  INV_X1 U603 ( .A(n674), .ZN(n515) );
  INV_X1 U604 ( .A(n524), .ZN(n516) );
  NAND2_X1 U605 ( .A1(n517), .A2(n516), .ZN(n519) );
  INV_X1 U606 ( .A(KEYINPUT84), .ZN(n518) );
  XNOR2_X2 U607 ( .A(n599), .B(KEYINPUT1), .ZN(n656) );
  XOR2_X1 U608 ( .A(KEYINPUT110), .B(KEYINPUT37), .Z(n521) );
  XOR2_X1 U609 ( .A(n521), .B(G125), .Z(n522) );
  XNOR2_X1 U610 ( .A(n544), .B(n522), .ZN(G27) );
  INV_X1 U611 ( .A(KEYINPUT19), .ZN(n523) );
  NAND2_X1 U612 ( .A1(n588), .A2(n525), .ZN(n526) );
  XNOR2_X1 U613 ( .A(n526), .B(KEYINPUT28), .ZN(n527) );
  OR2_X1 U614 ( .A1(n527), .A2(n599), .ZN(n552) );
  INV_X1 U615 ( .A(n537), .ZN(n528) );
  NAND2_X1 U616 ( .A1(n646), .A2(n528), .ZN(n645) );
  NAND2_X1 U617 ( .A1(KEYINPUT76), .A2(n645), .ZN(n529) );
  NOR2_X1 U618 ( .A1(n529), .A2(KEYINPUT47), .ZN(n532) );
  INV_X1 U619 ( .A(n648), .ZN(n530) );
  NOR2_X1 U620 ( .A1(n537), .A2(n530), .ZN(n641) );
  INV_X1 U621 ( .A(n641), .ZN(n531) );
  NAND2_X1 U622 ( .A1(n532), .A2(n531), .ZN(n536) );
  NAND2_X1 U623 ( .A1(n537), .A2(KEYINPUT76), .ZN(n533) );
  NOR2_X1 U624 ( .A1(n646), .A2(n648), .ZN(n605) );
  INV_X1 U625 ( .A(n605), .ZN(n677) );
  AND2_X1 U626 ( .A1(n533), .A2(n677), .ZN(n534) );
  NAND2_X1 U627 ( .A1(n534), .A2(KEYINPUT47), .ZN(n535) );
  NAND2_X1 U628 ( .A1(n536), .A2(n535), .ZN(n543) );
  NOR2_X1 U629 ( .A1(n537), .A2(KEYINPUT76), .ZN(n541) );
  NAND2_X1 U630 ( .A1(n549), .A2(n548), .ZN(n581) );
  OR2_X1 U631 ( .A1(n538), .A2(n581), .ZN(n540) );
  NOR2_X1 U632 ( .A1(n540), .A2(n539), .ZN(n643) );
  NOR2_X1 U633 ( .A1(n541), .A2(n643), .ZN(n542) );
  NAND2_X1 U634 ( .A1(n543), .A2(n542), .ZN(n545) );
  NOR2_X1 U635 ( .A1(n545), .A2(n544), .ZN(n559) );
  NAND2_X1 U636 ( .A1(n546), .A2(n674), .ZN(n547) );
  NOR2_X1 U637 ( .A1(n549), .A2(n548), .ZN(n676) );
  INV_X1 U638 ( .A(KEYINPUT41), .ZN(n550) );
  NAND2_X1 U639 ( .A1(n554), .A2(n646), .ZN(n556) );
  INV_X1 U640 ( .A(KEYINPUT40), .ZN(n555) );
  XNOR2_X1 U641 ( .A(n557), .B(KEYINPUT46), .ZN(n558) );
  AND2_X1 U642 ( .A1(n656), .A2(n674), .ZN(n561) );
  NAND2_X1 U643 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U644 ( .A(KEYINPUT43), .B(KEYINPUT102), .ZN(n563) );
  XNOR2_X1 U645 ( .A(n564), .B(n563), .ZN(n565) );
  AND2_X1 U646 ( .A1(n538), .A2(n565), .ZN(n651) );
  INV_X1 U647 ( .A(n651), .ZN(n566) );
  INV_X1 U648 ( .A(n567), .ZN(n568) );
  NAND2_X1 U649 ( .A1(n568), .A2(KEYINPUT2), .ZN(n569) );
  INV_X1 U650 ( .A(KEYINPUT0), .ZN(n577) );
  INV_X1 U651 ( .A(n570), .ZN(n575) );
  NOR2_X1 U652 ( .A1(G898), .A2(n726), .ZN(n723) );
  NAND2_X1 U653 ( .A1(n723), .A2(G902), .ZN(n572) );
  NAND2_X1 U654 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U655 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U656 ( .A(n596), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n660), .A2(n661), .ZN(n655) );
  NOR2_X1 U658 ( .A1(n579), .A2(n652), .ZN(n580) );
  XNOR2_X2 U659 ( .A(n583), .B(KEYINPUT22), .ZN(n595) );
  INV_X1 U660 ( .A(n660), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n592), .A2(n584), .ZN(n585) );
  NOR2_X1 U662 ( .A1(n585), .A2(n656), .ZN(n586) );
  NOR2_X1 U663 ( .A1(n588), .A2(n660), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n656), .A2(n589), .ZN(n590) );
  OR2_X1 U665 ( .A1(n595), .A2(n590), .ZN(n640) );
  XNOR2_X1 U666 ( .A(n591), .B(KEYINPUT44), .ZN(n608) );
  AND2_X1 U667 ( .A1(n592), .A2(n660), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n593), .A2(n656), .ZN(n594) );
  NOR2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n632) );
  INV_X1 U670 ( .A(n588), .ZN(n602) );
  NOR2_X1 U671 ( .A1(n597), .A2(n602), .ZN(n667) );
  NAND2_X1 U672 ( .A1(n596), .A2(n667), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT31), .ZN(n649) );
  NOR2_X1 U674 ( .A1(n599), .A2(n655), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n596), .A2(n600), .ZN(n601) );
  XNOR2_X1 U676 ( .A(n601), .B(KEYINPUT91), .ZN(n603) );
  AND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n635) );
  NOR2_X1 U678 ( .A1(n649), .A2(n635), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U680 ( .A1(n632), .A2(n606), .ZN(n607) );
  INV_X1 U681 ( .A(KEYINPUT45), .ZN(n609) );
  XOR2_X1 U682 ( .A(KEYINPUT79), .B(n612), .Z(n614) );
  INV_X1 U683 ( .A(KEYINPUT2), .ZN(n613) );
  NOR2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n706), .A2(G472), .ZN(n619) );
  XNOR2_X1 U686 ( .A(KEYINPUT105), .B(KEYINPUT62), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n619), .B(n618), .ZN(n620) );
  NAND2_X1 U689 ( .A1(n620), .A2(n699), .ZN(n622) );
  XNOR2_X1 U690 ( .A(KEYINPUT106), .B(KEYINPUT63), .ZN(n621) );
  XNOR2_X1 U691 ( .A(n622), .B(n621), .ZN(G57) );
  XOR2_X1 U692 ( .A(n623), .B(G131), .Z(G33) );
  NAND2_X1 U693 ( .A1(n706), .A2(G210), .ZN(n628) );
  XNOR2_X1 U694 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT55), .ZN(n626) );
  XNOR2_X1 U696 ( .A(n624), .B(n626), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n628), .B(n627), .ZN(n629) );
  NAND2_X1 U698 ( .A1(n629), .A2(n699), .ZN(n631) );
  XNOR2_X1 U699 ( .A(KEYINPUT83), .B(KEYINPUT56), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n631), .B(n630), .ZN(G51) );
  XNOR2_X1 U701 ( .A(G101), .B(n632), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n633), .B(KEYINPUT107), .ZN(G3) );
  NAND2_X1 U703 ( .A1(n635), .A2(n646), .ZN(n634) );
  XNOR2_X1 U704 ( .A(n634), .B(G104), .ZN(G6) );
  XNOR2_X1 U705 ( .A(KEYINPUT108), .B(KEYINPUT26), .ZN(n639) );
  XOR2_X1 U706 ( .A(G107), .B(KEYINPUT27), .Z(n637) );
  NAND2_X1 U707 ( .A1(n635), .A2(n648), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(G9) );
  XNOR2_X1 U710 ( .A(G110), .B(n640), .ZN(G12) );
  XNOR2_X1 U711 ( .A(G128), .B(n641), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n642), .B(KEYINPUT29), .ZN(G30) );
  XOR2_X1 U713 ( .A(G143), .B(n643), .Z(G45) );
  XOR2_X1 U714 ( .A(G146), .B(KEYINPUT109), .Z(n644) );
  XNOR2_X1 U715 ( .A(n645), .B(n644), .ZN(G48) );
  NAND2_X1 U716 ( .A1(n649), .A2(n646), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n647), .B(G113), .ZN(G15) );
  NAND2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n650), .B(G116), .ZN(G18) );
  XOR2_X1 U720 ( .A(G140), .B(n651), .Z(G42) );
  NOR2_X1 U721 ( .A1(n652), .A2(n673), .ZN(n653) );
  XOR2_X1 U722 ( .A(KEYINPUT118), .B(n653), .Z(n654) );
  NAND2_X1 U723 ( .A1(n726), .A2(n654), .ZN(n691) );
  XNOR2_X1 U724 ( .A(KEYINPUT51), .B(KEYINPUT115), .ZN(n670) );
  XOR2_X1 U725 ( .A(KEYINPUT113), .B(KEYINPUT50), .Z(n658) );
  NAND2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U728 ( .A(KEYINPUT112), .B(n659), .Z(n666) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT49), .B(n662), .Z(n663) );
  NOR2_X1 U731 ( .A1(n663), .A2(n588), .ZN(n664) );
  XNOR2_X1 U732 ( .A(n664), .B(KEYINPUT111), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n668) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U736 ( .A(n671), .B(KEYINPUT114), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n685) );
  OR2_X1 U738 ( .A1(n546), .A2(n674), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n680) );
  NAND2_X1 U740 ( .A1(n354), .A2(n677), .ZN(n679) );
  NAND2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U742 ( .A(KEYINPUT116), .B(n681), .Z(n682) );
  NOR2_X1 U743 ( .A1(n652), .A2(n682), .ZN(n683) );
  XOR2_X1 U744 ( .A(KEYINPUT117), .B(n683), .Z(n684) );
  NOR2_X1 U745 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U746 ( .A(KEYINPUT52), .B(n686), .ZN(n689) );
  NAND2_X1 U747 ( .A1(n687), .A2(G952), .ZN(n688) );
  NOR2_X1 U748 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U749 ( .A1(n691), .A2(n690), .ZN(n692) );
  AND2_X1 U750 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U751 ( .A1(n694), .A2(KEYINPUT2), .ZN(n695) );
  NAND2_X1 U752 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U753 ( .A(KEYINPUT119), .B(n697), .ZN(n698) );
  XNOR2_X1 U754 ( .A(KEYINPUT53), .B(n698), .ZN(G75) );
  INV_X1 U755 ( .A(n699), .ZN(n719) );
  NAND2_X1 U756 ( .A1(n706), .A2(G469), .ZN(n704) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n700) );
  XOR2_X1 U758 ( .A(n700), .B(KEYINPUT121), .Z(n701) );
  XNOR2_X1 U759 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U760 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U761 ( .A1(n719), .A2(n705), .ZN(G54) );
  NAND2_X1 U762 ( .A1(n706), .A2(G475), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X2 U764 ( .A1(n710), .A2(n719), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n711), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U766 ( .A1(n706), .A2(G478), .ZN(n714) );
  XOR2_X1 U767 ( .A(KEYINPUT122), .B(n712), .Z(n713) );
  XNOR2_X1 U768 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U769 ( .A1(n719), .A2(n715), .ZN(G63) );
  NAND2_X1 U770 ( .A1(n706), .A2(G217), .ZN(n717) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U772 ( .A1(n719), .A2(n718), .ZN(G66) );
  XNOR2_X1 U773 ( .A(n720), .B(KEYINPUT123), .ZN(n722) );
  XNOR2_X1 U774 ( .A(n722), .B(n721), .ZN(n724) );
  NOR2_X1 U775 ( .A1(n724), .A2(n723), .ZN(n733) );
  NAND2_X1 U776 ( .A1(n726), .A2(n725), .ZN(n730) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n727) );
  XNOR2_X1 U778 ( .A(KEYINPUT61), .B(n727), .ZN(n728) );
  NAND2_X1 U779 ( .A1(n728), .A2(G898), .ZN(n729) );
  NAND2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n731), .B(KEYINPUT124), .ZN(n732) );
  XNOR2_X1 U782 ( .A(n733), .B(n732), .ZN(G69) );
  XNOR2_X1 U783 ( .A(n734), .B(KEYINPUT125), .ZN(n735) );
  XNOR2_X1 U784 ( .A(n736), .B(n735), .ZN(n741) );
  XNOR2_X1 U785 ( .A(KEYINPUT126), .B(n741), .ZN(n737) );
  XNOR2_X1 U786 ( .A(G227), .B(n737), .ZN(n738) );
  NAND2_X1 U787 ( .A1(G900), .A2(n738), .ZN(n739) );
  NAND2_X1 U788 ( .A1(G953), .A2(n739), .ZN(n740) );
  XOR2_X1 U789 ( .A(KEYINPUT127), .B(n740), .Z(n744) );
  NAND2_X1 U790 ( .A1(n742), .A2(n411), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n744), .A2(n743), .ZN(G72) );
  XOR2_X1 U792 ( .A(n745), .B(G122), .Z(G24) );
  XNOR2_X1 U793 ( .A(G119), .B(n746), .ZN(G21) );
  XOR2_X1 U794 ( .A(n355), .B(G137), .Z(G39) );
endmodule

