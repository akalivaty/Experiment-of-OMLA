//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G107), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  AND3_X1   g010(.A1(new_n196), .A2(KEYINPUT4), .A3(G101), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n195), .A2(new_n191), .A3(new_n198), .A4(new_n193), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT78), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n199), .A2(new_n200), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT4), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(G101), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n197), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT64), .A2(G143), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT64), .A2(G143), .ZN(new_n211));
  OAI211_X1 g025(.A(KEYINPUT65), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n209), .B2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT66), .A3(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT64), .B(G143), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT65), .B1(new_n219), .B2(new_n209), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n208), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g035(.A1(KEYINPUT64), .A2(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT64), .A2(G143), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n222), .A2(KEYINPUT67), .A3(G146), .A4(new_n223), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n210), .A2(new_n211), .A3(new_n209), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n215), .B2(G146), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n224), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n206), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n221), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n205), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n227), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(new_n219), .B2(new_n209), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n219), .B2(new_n209), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n233), .B(new_n224), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n228), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT79), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n190), .A2(G104), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n198), .B1(new_n242), .B2(new_n193), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n194), .A2(KEYINPUT78), .A3(new_n198), .A4(new_n195), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n199), .A2(new_n200), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n210), .A2(new_n211), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n227), .B1(new_n247), .B2(G146), .ZN(new_n248));
  INV_X1    g062(.A(new_n224), .ZN(new_n249));
  OAI211_X1 g063(.A(KEYINPUT79), .B(new_n238), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n241), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT10), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT68), .A2(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G137), .ZN(new_n256));
  OR2_X1    g070(.A1(KEYINPUT68), .A2(KEYINPUT11), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(G137), .ZN(new_n259));
  INV_X1    g073(.A(G137), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G134), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT68), .A2(KEYINPUT11), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(G131), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n265));
  NOR2_X1   g079(.A1(KEYINPUT68), .A2(KEYINPUT11), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n262), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n256), .A2(new_n254), .ZN(new_n268));
  INV_X1    g082(.A(G131), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .A4(new_n259), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n264), .A2(new_n265), .A3(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(KEYINPUT69), .B(G131), .C1(new_n258), .C2(new_n263), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n209), .A2(G143), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n236), .B1(new_n274), .B2(KEYINPUT1), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n212), .A2(new_n217), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n275), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n238), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n233), .B2(new_n224), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n246), .B(KEYINPUT10), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n231), .A2(new_n253), .A3(new_n273), .A4(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(G110), .B(G140), .ZN(new_n285));
  INV_X1    g099(.A(G953), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G227), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n285), .B(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n244), .A2(new_n245), .ZN(new_n290));
  INV_X1    g104(.A(new_n243), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n279), .A2(new_n217), .A3(new_n212), .ZN(new_n293));
  INV_X1    g107(.A(new_n275), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n293), .A2(new_n294), .B1(new_n228), .B2(new_n238), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n246), .A2(new_n250), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n273), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(KEYINPUT12), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT80), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n273), .B1(new_n251), .B2(new_n296), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT12), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT81), .B1(new_n303), .B2(KEYINPUT12), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT81), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT12), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n290), .A2(new_n250), .A3(new_n291), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n310), .A2(new_n241), .B1(new_n295), .B2(new_n292), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n308), .B(new_n309), .C1(new_n311), .C2(new_n273), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n289), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n253), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n283), .B1(new_n205), .B2(new_n230), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n300), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n288), .B1(new_n317), .B2(new_n284), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n187), .B(new_n188), .C1(new_n314), .C2(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n284), .A2(new_n288), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n317), .ZN(new_n321));
  INV_X1    g135(.A(new_n284), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n306), .B2(new_n313), .ZN(new_n323));
  OAI211_X1 g137(.A(G469), .B(new_n321), .C1(new_n323), .C2(new_n288), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n187), .A2(new_n188), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n319), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G221), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT9), .B(G234), .Z(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT77), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n328), .B1(new_n330), .B2(new_n188), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G113), .B(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(new_n192), .ZN(new_n335));
  AND2_X1   g149(.A1(KEYINPUT71), .A2(G237), .ZN(new_n336));
  NOR2_X1   g150(.A1(KEYINPUT71), .A2(G237), .ZN(new_n337));
  OAI211_X1 g151(.A(G214), .B(new_n286), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n247), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT71), .B(G237), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n340), .A2(G143), .A3(G214), .A4(new_n286), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G131), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n341), .A3(new_n269), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G125), .ZN(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G140), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT16), .ZN(new_n350));
  OR3_X1    g164(.A1(new_n348), .A2(KEYINPUT16), .A3(G140), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(G146), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n347), .A2(new_n349), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT19), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT84), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT84), .B1(new_n347), .B2(new_n349), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n355), .B1(new_n358), .B2(new_n354), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n345), .B(new_n352), .C1(G146), .C2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n339), .A2(new_n341), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT18), .A2(G131), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n363), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n339), .A2(new_n341), .A3(new_n361), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n353), .A2(new_n209), .ZN(new_n367));
  OR3_X1    g181(.A1(new_n356), .A2(new_n357), .A3(new_n209), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n364), .A2(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n335), .B1(new_n360), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT17), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n343), .A2(new_n372), .A3(new_n344), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n342), .A2(KEYINPUT17), .A3(G131), .ZN(new_n374));
  INV_X1    g188(.A(new_n352), .ZN(new_n375));
  AOI21_X1  g189(.A(G146), .B1(new_n350), .B2(new_n351), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT86), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n376), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT86), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n352), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n373), .A2(new_n374), .A3(new_n377), .A4(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n370), .A3(new_n335), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT87), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n374), .A2(new_n377), .A3(new_n380), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n369), .B1(new_n384), .B2(new_n373), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n335), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n371), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(G475), .A2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT20), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n371), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n386), .B1(new_n385), .B2(new_n335), .ZN(new_n393));
  AND4_X1   g207(.A1(new_n386), .A2(new_n381), .A3(new_n370), .A4(new_n335), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(new_n389), .ZN(new_n397));
  OAI22_X1  g211(.A1(new_n393), .A2(new_n394), .B1(new_n335), .B2(new_n385), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n188), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n391), .A2(new_n397), .B1(new_n399), .B2(G475), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT88), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n219), .B2(new_n236), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n247), .A2(KEYINPUT88), .A3(G128), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT13), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n215), .A2(G128), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT89), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT13), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT88), .B1(new_n247), .B2(G128), .ZN(new_n408));
  NOR4_X1   g222(.A1(new_n210), .A2(new_n211), .A3(new_n401), .A4(new_n236), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT89), .ZN(new_n411));
  INV_X1    g225(.A(new_n405), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT13), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n406), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G134), .ZN(new_n416));
  AOI211_X1 g230(.A(G134), .B(new_n405), .C1(new_n402), .C2(new_n403), .ZN(new_n417));
  INV_X1    g231(.A(G116), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G122), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n418), .A2(G122), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(new_n190), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n420), .A2(new_n421), .A3(G107), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n416), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n419), .A2(KEYINPUT14), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT90), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n428), .A2(new_n429), .A3(new_n421), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n419), .A2(KEYINPUT14), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n190), .B1(new_n428), .B2(new_n429), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n424), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n402), .A2(new_n403), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n255), .B1(new_n435), .B2(new_n412), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n436), .B2(new_n417), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT91), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n434), .B(new_n439), .C1(new_n417), .C2(new_n436), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n330), .A2(G217), .A3(new_n286), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n427), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT92), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT92), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n427), .A2(new_n441), .A3(new_n446), .A4(new_n443), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n427), .A2(new_n441), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n442), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n188), .ZN(new_n451));
  INV_X1    g265(.A(G478), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT15), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n453), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(new_n188), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(G898), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n188), .B1(G234), .B2(G237), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(G953), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(G234), .A2(G237), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(G952), .A3(new_n286), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n462), .B(KEYINPUT93), .Z(new_n463));
  NAND4_X1  g277(.A1(new_n400), .A2(new_n454), .A3(new_n456), .A4(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n333), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G217), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n466), .B1(G234), .B2(new_n188), .ZN(new_n467));
  NOR2_X1   g281(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT23), .ZN(new_n469));
  INV_X1    g283(.A(G119), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(G128), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n236), .A2(KEYINPUT23), .A3(G119), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n471), .B(new_n472), .C1(G119), .C2(new_n236), .ZN(new_n473));
  XNOR2_X1  g287(.A(G119), .B(G128), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT24), .B(G110), .Z(new_n475));
  AOI22_X1  g289(.A1(new_n473), .A2(G110), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n375), .B2(new_n376), .ZN(new_n477));
  OAI22_X1  g291(.A1(new_n473), .A2(G110), .B1(new_n474), .B2(new_n475), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n352), .A3(new_n367), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT22), .B(G137), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n286), .A2(G221), .A3(G234), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n477), .A2(new_n479), .A3(new_n483), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n468), .B1(new_n487), .B2(G902), .ZN(new_n488));
  NAND2_X1  g302(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n487), .A2(G902), .A3(new_n468), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n467), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n467), .A2(G902), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n493), .B(KEYINPUT76), .Z(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n485), .A2(new_n495), .A3(new_n486), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n470), .A2(G116), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n418), .A2(G119), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT2), .B(G113), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G116), .B(G119), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n504), .A2(KEYINPUT70), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(KEYINPUT70), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n503), .B1(new_n507), .B2(new_n502), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n261), .A2(new_n259), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G131), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n270), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n280), .B2(new_n282), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n271), .A2(new_n221), .A3(new_n229), .A4(new_n272), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n514), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n509), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n340), .A2(G210), .A3(new_n286), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT27), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT26), .B(G101), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n514), .A2(new_n516), .A3(new_n508), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT31), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT72), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n523), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  OAI22_X1  g345(.A1(new_n273), .A2(new_n230), .B1(new_n295), .B2(new_n512), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n509), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n530), .B1(new_n533), .B2(new_n524), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT73), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n524), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n508), .B1(new_n514), .B2(new_n516), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n535), .B(KEYINPUT28), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n529), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n525), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n525), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n528), .A2(new_n541), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT32), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n519), .A2(new_n524), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT29), .B1(new_n551), .B2(new_n529), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT28), .B1(new_n537), .B2(new_n538), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n539), .A3(new_n531), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n552), .B1(new_n555), .B2(new_n529), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT74), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n531), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n524), .A2(KEYINPUT74), .A3(new_n530), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n553), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n523), .A2(KEYINPUT29), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n556), .B(new_n188), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G472), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n546), .A2(KEYINPUT32), .A3(new_n547), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n550), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G214), .B1(G237), .B2(G902), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT82), .ZN(new_n567));
  OAI21_X1  g381(.A(G113), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT5), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n569), .B1(new_n507), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n503), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n246), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n205), .B2(new_n508), .ZN(new_n574));
  XNOR2_X1  g388(.A(G110), .B(G122), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n575), .B(new_n573), .C1(new_n205), .C2(new_n508), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(KEYINPUT6), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n348), .B1(new_n221), .B2(new_n229), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n295), .A2(new_n348), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G224), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(G953), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n583), .B(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT6), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n574), .A2(new_n587), .A3(new_n576), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n579), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n585), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT7), .A4(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n280), .A2(G125), .A3(new_n282), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT7), .ZN(new_n593));
  OAI22_X1  g407(.A1(new_n592), .A2(new_n580), .B1(new_n593), .B2(new_n585), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n292), .A2(new_n571), .A3(new_n572), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n501), .A2(new_n570), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n572), .B1(new_n596), .B2(new_n568), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n246), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n575), .B(KEYINPUT83), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT8), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n595), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n591), .A2(new_n594), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n603), .B2(new_n578), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n589), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(G210), .B1(G237), .B2(G902), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n589), .A2(new_n604), .A3(new_n606), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n567), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n465), .A2(new_n498), .A3(new_n565), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  INV_X1    g426(.A(G472), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(KEYINPUT94), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n546), .B2(new_n188), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n525), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT72), .B1(new_n525), .B2(KEYINPUT31), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n555), .A2(new_n529), .B1(new_n542), .B2(new_n543), .ZN(new_n621));
  AOI21_X1  g435(.A(G902), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n615), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n617), .A2(new_n498), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n333), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n427), .A2(new_n441), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n443), .A2(KEYINPUT95), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n450), .A2(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n452), .A2(G902), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n631), .A2(new_n632), .B1(new_n452), .B2(new_n451), .ZN(new_n633));
  INV_X1    g447(.A(new_n567), .ZN(new_n634));
  INV_X1    g448(.A(new_n609), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n606), .B1(new_n589), .B2(new_n604), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n634), .B(new_n463), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n633), .A2(new_n637), .A3(new_n400), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n624), .A2(new_n625), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NAND3_X1  g455(.A1(new_n617), .A2(new_n623), .A3(new_n498), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n333), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n454), .A2(new_n456), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n400), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n645), .A2(new_n637), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n484), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n480), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n495), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n492), .A2(new_n653), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n610), .A2(new_n617), .A3(new_n623), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n465), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT96), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT97), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n656), .B(new_n659), .ZN(G12));
  NOR2_X1   g474(.A1(new_n286), .A2(G900), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n458), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n662), .A2(KEYINPUT98), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(KEYINPUT98), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n461), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n456), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n455), .B1(new_n450), .B2(new_n188), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n400), .B(new_n665), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n333), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n610), .A2(new_n654), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n669), .A2(new_n565), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n669), .A2(KEYINPUT99), .A3(new_n565), .A4(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(new_n665), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n625), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n608), .A2(new_n609), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT38), .Z(new_n682));
  NOR4_X1   g496(.A1(new_n682), .A2(new_n567), .A3(new_n645), .A4(new_n400), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n546), .A2(KEYINPUT32), .A3(new_n547), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT32), .B1(new_n546), .B2(new_n547), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n551), .A2(new_n523), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n533), .A2(new_n529), .A3(new_n524), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n188), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n654), .B1(new_n687), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n680), .A2(new_n683), .A3(new_n684), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n219), .ZN(G45));
  INV_X1    g509(.A(new_n665), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n391), .A2(new_n397), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n399), .A2(G475), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n450), .A2(new_n626), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n629), .A2(new_n630), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n700), .A3(new_n632), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n451), .A2(new_n452), .ZN(new_n702));
  AOI221_X4 g516(.A(new_n696), .B1(new_n697), .B2(new_n698), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n565), .A2(new_n625), .A3(new_n671), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n209), .ZN(G48));
  INV_X1    g519(.A(KEYINPUT100), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n187), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n306), .A2(new_n313), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n318), .B1(new_n708), .B2(new_n320), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n707), .B1(new_n709), .B2(G902), .ZN(new_n710));
  OAI221_X1 g524(.A(new_n188), .B1(new_n706), .B2(new_n187), .C1(new_n314), .C2(new_n318), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n332), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n565), .A2(new_n638), .A3(new_n713), .A4(new_n498), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT101), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n714), .B(new_n716), .ZN(G15));
  NAND4_X1  g531(.A1(new_n647), .A2(new_n565), .A3(new_n498), .A4(new_n713), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NOR2_X1   g533(.A1(new_n712), .A2(new_n464), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n565), .A2(new_n720), .A3(new_n671), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  INV_X1    g536(.A(new_n463), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n567), .B1(new_n697), .B2(new_n698), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n644), .A2(new_n724), .A3(new_n681), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n644), .A2(new_n724), .A3(new_n681), .A4(KEYINPUT103), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n560), .A2(new_n529), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n526), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n544), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n731), .B1(new_n730), .B2(new_n526), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n547), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n735), .B1(new_n622), .B2(new_n613), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n736), .A2(new_n497), .A3(new_n712), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n729), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  INV_X1    g553(.A(new_n547), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n529), .A2(new_n560), .B1(new_n525), .B2(KEYINPUT31), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n741), .A2(new_n731), .B1(new_n543), .B2(new_n542), .ZN(new_n742));
  INV_X1    g556(.A(new_n734), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n613), .B1(new_n546), .B2(new_n188), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n610), .A2(new_n710), .A3(new_n711), .A4(new_n332), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n703), .A4(new_n654), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT104), .ZN(new_n749));
  INV_X1    g563(.A(new_n654), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n744), .A2(new_n745), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n703), .A4(new_n747), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  AOI21_X1  g569(.A(new_n497), .B1(new_n687), .B2(new_n563), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n635), .A2(new_n636), .A3(new_n567), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n327), .A2(new_n332), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n756), .A2(KEYINPUT42), .A3(new_n703), .A4(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n565), .A2(new_n758), .A3(new_n498), .A4(new_n703), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  INV_X1    g578(.A(new_n668), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n565), .A2(new_n758), .A3(new_n498), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  OR3_X1    g581(.A1(new_n633), .A2(KEYINPUT43), .A3(new_n646), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT43), .B1(new_n633), .B2(new_n646), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n750), .B1(new_n617), .B2(new_n623), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(KEYINPUT44), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT105), .A3(new_n757), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n771), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT105), .B1(new_n772), .B2(new_n757), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT106), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n778), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n776), .A4(new_n773), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n321), .B1(new_n323), .B2(new_n288), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n187), .B1(new_n783), .B2(new_n784), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n326), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n326), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n319), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n332), .A3(new_n678), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n779), .A2(new_n782), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT107), .B(G137), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G39));
  NAND2_X1  g611(.A1(new_n792), .A2(new_n332), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n332), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n701), .A2(new_n702), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n646), .A3(new_n665), .ZN(new_n804));
  INV_X1    g618(.A(new_n757), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n565), .A2(new_n804), .A3(new_n498), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT108), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n802), .A2(new_n809), .A3(new_n806), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  NOR3_X1   g626(.A1(new_n712), .A2(new_n805), .A3(new_n461), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n770), .A2(new_n756), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n815));
  AND2_X1   g629(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n814), .A2(new_n816), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n768), .A2(new_n769), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n461), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n498), .A3(new_n746), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n610), .A2(new_n710), .A3(new_n711), .A4(new_n332), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n550), .A2(new_n564), .A3(new_n692), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n497), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n825), .A2(new_n813), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n633), .A2(new_n400), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(G952), .A3(new_n286), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n817), .A2(new_n818), .A3(new_n823), .A4(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n737), .A2(new_n567), .A3(new_n682), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n820), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n820), .A3(KEYINPUT113), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT114), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n831), .A2(KEYINPUT50), .A3(new_n820), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n834), .A2(new_n840), .A3(new_n835), .A4(new_n836), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n826), .A2(new_n400), .A3(new_n633), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n735), .B(new_n654), .C1(new_n613), .C2(new_n622), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n770), .A2(new_n813), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n710), .A2(new_n711), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n800), .B(new_n801), .C1(new_n332), .C2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n821), .A2(new_n805), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n842), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n830), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n851), .A2(KEYINPUT115), .A3(new_n852), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n704), .B1(new_n674), .B2(new_n675), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n327), .A2(new_n332), .A3(new_n665), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n824), .A2(new_n861), .A3(new_n750), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n727), .A2(new_n728), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n749), .A2(new_n753), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n860), .A2(new_n864), .A3(KEYINPUT52), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT52), .B1(new_n860), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n738), .A2(new_n611), .A3(new_n714), .A4(new_n718), .ZN(new_n868));
  INV_X1    g682(.A(new_n637), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT109), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n666), .B2(new_n667), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n454), .A2(KEYINPUT109), .A3(new_n456), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n871), .A2(new_n872), .A3(new_n400), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n624), .A2(new_n625), .A3(new_n869), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n656), .A3(new_n639), .A4(new_n721), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n758), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n400), .A2(new_n654), .A3(new_n665), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n871), .B2(new_n872), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n565), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n746), .A2(new_n703), .A3(new_n654), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n766), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT110), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT110), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n703), .A2(new_n751), .B1(new_n565), .B2(new_n879), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n885), .B(new_n766), .C1(new_n886), .C2(new_n877), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n876), .A2(new_n763), .A3(new_n884), .A4(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n859), .B1(new_n867), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n884), .A2(new_n763), .A3(new_n887), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n565), .A2(new_n498), .A3(new_n713), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n892), .A2(new_n647), .B1(new_n729), .B2(new_n737), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n611), .A2(new_n714), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n869), .A2(new_n871), .A3(new_n872), .A4(new_n400), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n642), .A2(new_n895), .A3(new_n333), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n565), .A2(new_n720), .A3(new_n671), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n643), .A2(new_n638), .B1(new_n655), .B2(new_n465), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n893), .A2(new_n894), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n891), .A2(new_n900), .A3(new_n859), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT52), .ZN(new_n902));
  INV_X1    g716(.A(new_n704), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n670), .B1(new_n687), .B2(new_n563), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT99), .B1(new_n904), .B2(new_n669), .ZN(new_n905));
  AND4_X1   g719(.A1(KEYINPUT99), .A2(new_n669), .A3(new_n565), .A4(new_n671), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n693), .A2(new_n863), .A3(new_n861), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n844), .A2(new_n804), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n752), .B1(new_n909), .B2(new_n747), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n844), .A2(new_n804), .A3(new_n822), .A4(KEYINPUT104), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n902), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n860), .A2(new_n864), .A3(KEYINPUT52), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(KEYINPUT111), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT111), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n866), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n901), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n889), .A2(new_n890), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n891), .A2(new_n900), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n915), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(KEYINPUT112), .A3(new_n859), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n866), .B2(new_n865), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n859), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT112), .B1(new_n921), .B2(new_n859), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n858), .B(new_n919), .C1(new_n890), .C2(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(G952), .A2(G953), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n847), .A2(KEYINPUT49), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n847), .A2(KEYINPUT49), .ZN(new_n931));
  NOR4_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n646), .A4(new_n633), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n331), .A2(new_n567), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n932), .A2(new_n682), .A3(new_n825), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n929), .A2(new_n934), .ZN(G75));
  AOI21_X1  g749(.A(new_n188), .B1(new_n889), .B2(new_n918), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT56), .B1(new_n936), .B2(G210), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n579), .A2(new_n588), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(new_n586), .Z(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT55), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n937), .A2(KEYINPUT117), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT117), .B1(new_n937), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n937), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT118), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT118), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n937), .A2(new_n947), .A3(new_n941), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n286), .A2(G952), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n944), .A2(new_n949), .A3(new_n951), .ZN(G51));
  NAND2_X1  g766(.A1(new_n889), .A2(new_n918), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n919), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n325), .B(KEYINPUT57), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n318), .B2(new_n314), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n936), .A2(new_n785), .A3(new_n786), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT119), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n950), .B1(new_n958), .B2(new_n960), .ZN(G54));
  NAND3_X1  g775(.A1(new_n936), .A2(KEYINPUT58), .A3(G475), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT120), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n962), .A2(new_n963), .A3(new_n388), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n951), .B1(new_n962), .B2(new_n388), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n962), .B2(new_n388), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G60));
  OAI21_X1  g781(.A(new_n919), .B1(new_n926), .B2(new_n890), .ZN(new_n968));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT59), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n631), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n955), .A2(new_n631), .A3(new_n971), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n951), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(G63));
  XNOR2_X1  g789(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT121), .ZN(new_n977));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT60), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n977), .B1(new_n953), .B2(new_n980), .ZN(new_n981));
  AOI211_X1 g795(.A(KEYINPUT121), .B(new_n979), .C1(new_n889), .C2(new_n918), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n487), .B(KEYINPUT123), .Z(new_n984));
  AOI21_X1  g798(.A(new_n950), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n652), .B(KEYINPUT122), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n981), .B2(new_n982), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n976), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n953), .A2(new_n980), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT121), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n953), .A2(new_n977), .A3(new_n980), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n991), .A3(new_n984), .ZN(new_n992));
  AND4_X1   g806(.A1(new_n951), .A2(new_n992), .A3(new_n987), .A4(new_n976), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n988), .A2(new_n993), .ZN(G66));
  OAI21_X1  g808(.A(G953), .B1(new_n457), .B2(new_n584), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n876), .B2(G953), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n938), .B1(G898), .B2(new_n286), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G69));
  NOR2_X1   g812(.A1(new_n517), .A2(new_n518), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(new_n359), .Z(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n811), .A2(new_n795), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n794), .A2(new_n756), .A3(new_n863), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n860), .A2(new_n754), .ZN(new_n1004));
  AND4_X1   g818(.A1(new_n763), .A2(new_n1003), .A3(new_n1004), .A4(new_n766), .ZN(new_n1005));
  AOI21_X1  g819(.A(G953), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1001), .B1(new_n1006), .B2(new_n661), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n756), .A2(new_n757), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n873), .A2(new_n827), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1008), .A2(new_n679), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1004), .A2(KEYINPUT62), .A3(new_n694), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n694), .A2(new_n860), .A3(new_n754), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT62), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1010), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n811), .A2(new_n1015), .A3(new_n795), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT125), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT125), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n811), .A2(new_n1015), .A3(new_n795), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(G953), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1007), .B1(new_n1020), .B2(new_n1001), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n286), .B1(G227), .B2(G900), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1022), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1007), .B(new_n1024), .C1(new_n1020), .C2(new_n1001), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(G72));
  NAND3_X1  g840(.A1(new_n1002), .A2(new_n876), .A3(new_n1005), .ZN(new_n1027));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n551), .A2(new_n523), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1031), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1033), .A2(new_n688), .A3(new_n1029), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1034), .B(KEYINPUT127), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1032), .B(new_n951), .C1(new_n926), .C2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1017), .A2(new_n876), .A3(new_n1019), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(new_n1029), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n689), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(KEYINPUT126), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT126), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1038), .A2(new_n1041), .A3(new_n689), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1036), .B1(new_n1040), .B2(new_n1042), .ZN(G57));
endmodule


