//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n207), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT64), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n212), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G97), .B(G107), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  AND2_X1   g0046(.A1(new_n246), .A2(new_n218), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n207), .A2(G33), .ZN(new_n249));
  OR2_X1    g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n247), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n202), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n247), .B1(G1), .B2(new_n207), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n256), .B1(new_n257), .B2(new_n202), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  OR2_X1    g0059(.A1(new_n259), .A2(KEYINPUT9), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(KEYINPUT9), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT10), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT66), .ZN(new_n264));
  AND2_X1   g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n218), .ZN(new_n266));
  AND2_X1   g0066(.A1(G1), .A2(G13), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(KEYINPUT66), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n266), .A2(new_n269), .A3(new_n271), .A4(G274), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n266), .A2(new_n269), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(new_n271), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(G226), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n282), .A2(G223), .B1(new_n285), .B2(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n280), .A2(new_n281), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G222), .A3(new_n277), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n265), .A2(new_n218), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n276), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G200), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n276), .A2(new_n291), .A3(G190), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n262), .A2(new_n263), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n260), .A2(new_n294), .A3(new_n261), .ZN(new_n296));
  INV_X1    g0096(.A(new_n293), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT10), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n259), .B1(new_n292), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(G179), .B2(new_n292), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n290), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n282), .A2(G238), .B1(new_n285), .B2(G107), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n287), .A2(G232), .A3(new_n277), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI211_X1 g0107(.A(new_n273), .B(new_n307), .C1(G244), .C2(new_n275), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G20), .A2(G77), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n207), .A2(new_n279), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n310), .B1(new_n248), .B2(new_n311), .C1(new_n249), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n246), .A2(new_n218), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G77), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n255), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n257), .B2(new_n316), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n309), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n308), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n308), .A2(G190), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n324), .B(new_n319), .C1(new_n325), .C2(new_n308), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n303), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n248), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n255), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n328), .B2(new_n257), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n266), .A2(new_n269), .A3(G232), .A4(new_n270), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n272), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(G223), .A2(G1698), .ZN(new_n334));
  INV_X1    g0134(.A(G226), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(G1698), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(new_n287), .B1(G33), .B2(G87), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n333), .B1(new_n304), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n325), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n337), .B2(new_n304), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n335), .A2(G1698), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G223), .B2(G1698), .ZN(new_n343));
  INV_X1    g0143(.A(G87), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n343), .A2(new_n285), .B1(new_n279), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(KEYINPUT72), .A3(new_n290), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n341), .A2(new_n333), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n339), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT69), .ZN(new_n354));
  AND2_X1   g0154(.A1(G58), .A2(G68), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n354), .B(G20), .C1(new_n355), .C2(new_n201), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n251), .A2(G159), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G58), .A2(G68), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n215), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n354), .B1(new_n360), .B2(G20), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT70), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n355), .B2(new_n201), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT69), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT70), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n356), .A4(new_n357), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT7), .B1(new_n287), .B2(G20), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n285), .A2(new_n368), .A3(new_n207), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(G68), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n362), .A2(KEYINPUT16), .A3(new_n366), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n362), .A2(new_n366), .A3(new_n370), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n366), .A2(new_n370), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n356), .A2(new_n357), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n365), .B1(new_n379), .B2(new_n364), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n372), .B(new_n375), .C1(new_n378), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n314), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n331), .B(new_n353), .C1(new_n377), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT17), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n383), .B(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n381), .A2(new_n314), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n373), .A2(new_n376), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n330), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n341), .A2(new_n333), .A3(new_n321), .A4(new_n346), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT73), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n390), .A2(new_n391), .B1(new_n300), .B2(new_n338), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(KEYINPUT73), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT18), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n331), .B1(new_n377), .B2(new_n382), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n390), .A2(new_n391), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n338), .A2(new_n300), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n397), .A2(new_n393), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n385), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(G232), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n404));
  OAI211_X1 g0204(.A(G226), .B(new_n277), .C1(new_n283), .C2(new_n284), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n407), .A2(new_n290), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n266), .A2(new_n269), .A3(G238), .A4(new_n270), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n272), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT13), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n290), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(new_n272), .A4(new_n409), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(KEYINPUT67), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT67), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(KEYINPUT13), .C1(new_n408), .C2(new_n410), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n417), .A3(G169), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n415), .A2(new_n417), .A3(KEYINPUT14), .A4(G169), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n411), .A2(G179), .A3(new_n414), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n249), .A2(new_n316), .B1(new_n207), .B2(G68), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n311), .A2(new_n202), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n314), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT11), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT12), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n255), .B2(new_n214), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n254), .A2(KEYINPUT12), .A3(G68), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n257), .A2(new_n214), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n427), .A2(new_n428), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n429), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n424), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n414), .A2(G190), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n437), .B2(new_n411), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n415), .A2(new_n417), .A3(G200), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT68), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT68), .B1(new_n438), .B2(new_n439), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n327), .A2(new_n403), .A3(new_n436), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G41), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n449), .A3(G274), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT78), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT5), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(G41), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(G41), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n265), .A2(new_n264), .A3(new_n218), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT66), .B1(new_n267), .B2(new_n268), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n456), .A2(new_n459), .A3(KEYINPUT79), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT79), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n462), .A2(new_n454), .A3(new_n453), .A4(new_n447), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n274), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n446), .A2(KEYINPUT5), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n449), .A2(new_n454), .A3(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n467), .A2(new_n266), .A3(new_n269), .ZN(new_n468));
  OAI211_X1 g0268(.A(G250), .B(new_n277), .C1(new_n283), .C2(new_n284), .ZN(new_n469));
  OAI211_X1 g0269(.A(G257), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G294), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(G264), .A2(new_n468), .B1(new_n472), .B2(new_n290), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT84), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT84), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n465), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(G169), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n465), .A2(new_n473), .A3(G179), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n344), .B1(new_n481), .B2(KEYINPUT22), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n287), .A2(new_n207), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(KEYINPUT81), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(KEYINPUT81), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n287), .A2(new_n482), .A3(new_n207), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  INV_X1    g0288(.A(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(G20), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n490), .B(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G116), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n493), .B2(G20), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n488), .B1(G20), .B2(new_n489), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n485), .A2(new_n487), .A3(new_n491), .A4(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n247), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n491), .A2(new_n496), .ZN(new_n500));
  INV_X1    g0300(.A(new_n498), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n500), .A2(new_n487), .A3(new_n485), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n206), .A2(G33), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n247), .A2(new_n254), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT25), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n254), .A2(new_n506), .A3(G107), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n254), .B2(G107), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n505), .A2(G107), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n480), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n510), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n499), .B2(new_n502), .ZN(new_n514));
  AOI21_X1  g0314(.A(G190), .B1(new_n475), .B2(new_n477), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n474), .A2(new_n325), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G238), .B(new_n277), .C1(new_n283), .C2(new_n284), .ZN(new_n519));
  OAI211_X1 g0319(.A(G244), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n520), .A3(new_n493), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n522));
  INV_X1    g0322(.A(G250), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n449), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n521), .A2(new_n290), .B1(new_n459), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G190), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n207), .B(G68), .C1(new_n283), .C2(new_n284), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  INV_X1    g0328(.A(G97), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n249), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n406), .A2(new_n528), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(G20), .ZN(new_n532));
  NOR3_X1   g0332(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n527), .B(new_n530), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(new_n314), .B1(new_n255), .B2(new_n312), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n505), .A2(G87), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n526), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n525), .A2(new_n325), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n525), .A2(new_n321), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n314), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n312), .A2(new_n255), .ZN(new_n541));
  INV_X1    g0341(.A(new_n312), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n505), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n525), .A2(G169), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n537), .A2(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n512), .A2(new_n518), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G116), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n246), .A2(new_n218), .B1(G20), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G283), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n552), .B(new_n207), .C1(G33), .C2(new_n529), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n551), .A2(KEYINPUT20), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT20), .B1(new_n551), .B2(new_n553), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n254), .A2(G116), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n505), .B2(G116), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G264), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n560));
  OAI211_X1 g0360(.A(G257), .B(new_n277), .C1(new_n283), .C2(new_n284), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n280), .A2(G303), .A3(new_n281), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(G270), .A2(new_n468), .B1(new_n563), .B2(new_n290), .ZN(new_n564));
  AND4_X1   g0364(.A1(G179), .A2(new_n559), .A3(new_n465), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n465), .A2(new_n564), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT80), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT80), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n465), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n300), .B1(new_n556), .B2(new_n558), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n565), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n465), .A2(new_n564), .A3(new_n568), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n568), .B1(new_n465), .B2(new_n564), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n352), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n567), .A2(G200), .A3(new_n569), .ZN(new_n577));
  INV_X1    g0377(.A(new_n559), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n574), .A2(new_n575), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(KEYINPUT21), .A3(new_n570), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n573), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n468), .A2(G257), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n465), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n287), .A2(G250), .A3(G1698), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n552), .ZN(new_n586));
  OAI211_X1 g0386(.A(G244), .B(new_n277), .C1(new_n283), .C2(new_n284), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT4), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n586), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT77), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n290), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n282), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n587), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT4), .B1(new_n587), .B2(KEYINPUT76), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n593), .B(new_n595), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n584), .B(new_n321), .C1(new_n594), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n505), .A2(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n255), .A2(new_n529), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n367), .A2(G107), .A3(new_n369), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n251), .A2(G77), .ZN(new_n605));
  XNOR2_X1  g0405(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n242), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n529), .A2(G107), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(new_n606), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n604), .B(new_n605), .C1(new_n609), .C2(new_n207), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n603), .B1(new_n610), .B2(new_n314), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n465), .A2(new_n583), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n304), .B1(new_n614), .B2(KEYINPUT77), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n615), .B2(new_n598), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n600), .B(new_n612), .C1(G169), .C2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n584), .B(G190), .C1(new_n594), .C2(new_n599), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n618), .B(new_n611), .C1(new_n325), .C2(new_n616), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n549), .A2(new_n582), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n445), .A2(new_n621), .ZN(G372));
  AND2_X1   g0422(.A1(new_n438), .A2(new_n439), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n323), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n385), .B1(new_n624), .B2(new_n436), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n299), .B1(new_n625), .B2(new_n402), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n302), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT86), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n573), .A2(new_n629), .A3(new_n581), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n573), .B2(new_n581), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n512), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT85), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n459), .A2(new_n633), .A3(new_n524), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n524), .A2(new_n266), .A3(new_n269), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT85), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n521), .A2(new_n290), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n325), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(G169), .B1(new_n637), .B2(new_n638), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n537), .A2(new_n639), .B1(new_n545), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n518), .A2(new_n617), .A3(new_n619), .A4(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n632), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT87), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n545), .A2(new_n640), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n612), .B1(new_n616), .B2(G169), .ZN(new_n648));
  INV_X1    g0448(.A(new_n600), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n648), .A2(new_n649), .A3(new_n641), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT26), .B1(new_n617), .B2(new_n547), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n646), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n584), .B1(new_n594), .B2(new_n599), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n611), .B1(new_n655), .B2(new_n300), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n656), .A2(new_n642), .A3(new_n651), .A4(new_n600), .ZN(new_n657));
  INV_X1    g0457(.A(new_n647), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n653), .A2(new_n657), .A3(new_n646), .A4(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n645), .B1(new_n654), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n628), .B1(new_n444), .B2(new_n662), .ZN(G369));
  NOR2_X1   g0463(.A1(new_n630), .A2(new_n631), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT88), .Z(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n578), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n582), .B2(new_n671), .ZN(new_n673));
  INV_X1    g0473(.A(new_n477), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n476), .B1(new_n465), .B2(new_n473), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n348), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n511), .B1(new_n676), .B2(new_n516), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n514), .B1(new_n478), .B2(new_n479), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n514), .B2(new_n670), .ZN(new_n680));
  INV_X1    g0480(.A(new_n670), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n673), .A2(G330), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n681), .B1(new_n573), .B2(new_n581), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n679), .A2(new_n685), .B1(new_n678), .B2(new_n670), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(G399));
  NAND2_X1  g0487(.A1(new_n533), .A2(new_n550), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT89), .Z(new_n689));
  INV_X1    g0489(.A(new_n210), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n689), .A2(new_n691), .A3(new_n206), .ZN(new_n692));
  INV_X1    g0492(.A(new_n691), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n692), .A2(KEYINPUT90), .B1(new_n216), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(KEYINPUT90), .B2(new_n692), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n656), .A2(new_n548), .A3(new_n651), .A4(new_n600), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n698), .A2(new_n658), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT26), .B1(new_n617), .B2(new_n641), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n512), .A2(new_n581), .A3(new_n573), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n699), .B(new_n700), .C1(new_n643), .C2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n697), .B1(new_n702), .B2(new_n670), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n653), .A2(new_n658), .A3(new_n657), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT87), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n659), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n681), .B1(new_n706), .B2(new_n645), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n703), .B1(new_n707), .B2(new_n697), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT91), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n566), .A2(new_n321), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n473), .A2(new_n525), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n710), .B1(new_n713), .B2(new_n655), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n616), .A2(KEYINPUT30), .A3(new_n711), .A4(new_n712), .ZN(new_n715));
  AOI21_X1  g0515(.A(G179), .B1(new_n637), .B2(new_n638), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n716), .A2(new_n474), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n580), .A2(new_n717), .A3(new_n655), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n714), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n681), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT31), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n722), .A3(new_n681), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n621), .A2(new_n670), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G330), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n709), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n677), .A2(new_n678), .A3(new_n547), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n573), .A2(new_n579), .A3(new_n581), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n612), .B1(new_n655), .B2(G200), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n600), .A2(new_n656), .B1(new_n729), .B2(new_n618), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n727), .A2(new_n728), .A3(new_n730), .A4(new_n670), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n722), .B1(new_n719), .B2(new_n681), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n719), .A2(new_n722), .A3(new_n681), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT91), .A3(G330), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n726), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n708), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n696), .B1(new_n738), .B2(G1), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT92), .Z(G364));
  AND2_X1   g0540(.A1(new_n207), .A2(G13), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n206), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n691), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n673), .B2(G330), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G330), .B2(new_n673), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n690), .A2(new_n285), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(G355), .B(KEYINPUT93), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n748), .A2(new_n749), .B1(G116), .B2(new_n210), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n690), .A2(new_n287), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n448), .B2(new_n217), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n241), .A2(new_n448), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n218), .B1(G20), .B2(new_n300), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n744), .B1(new_n755), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n207), .A2(new_n321), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n764), .A2(new_n325), .A3(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n766), .A2(new_n316), .B1(new_n768), .B2(new_n214), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n207), .A2(new_n325), .A3(G179), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n348), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n489), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n344), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n769), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n351), .A2(new_n325), .A3(new_n764), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n285), .B1(new_n776), .B2(G50), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n207), .B1(new_n778), .B2(G190), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT95), .Z(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G97), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n778), .A2(G20), .A3(new_n348), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n785));
  XNOR2_X1  g0585(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n351), .A2(G200), .A3(new_n764), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(G58), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n775), .A2(new_n777), .A3(new_n781), .A4(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G303), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n285), .B1(new_n773), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n776), .ZN(new_n792));
  INV_X1    g0592(.A(G326), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n791), .B(new_n794), .C1(G311), .C2(new_n765), .ZN(new_n795));
  INV_X1    g0595(.A(new_n779), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G294), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n787), .A2(G322), .B1(new_n767), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n795), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  INV_X1    g0601(.A(G329), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n771), .A2(new_n801), .B1(new_n802), .B2(new_n782), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT96), .Z(new_n804));
  OAI21_X1  g0604(.A(new_n789), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n762), .B1(new_n805), .B2(new_n759), .ZN(new_n806));
  INV_X1    g0606(.A(new_n758), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n673), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n746), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  OAI21_X1  g0610(.A(new_n326), .B1(new_n319), .B2(new_n670), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n323), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n320), .A2(new_n322), .A3(new_n670), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n707), .B(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n744), .B1(new_n816), .B2(new_n736), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n736), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n768), .A2(new_n801), .ZN(new_n819));
  INV_X1    g0619(.A(new_n782), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n287), .B(new_n819), .C1(G311), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n787), .ZN(new_n822));
  INV_X1    g0622(.A(G294), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n822), .A2(new_n823), .B1(new_n489), .B2(new_n773), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G116), .B2(new_n765), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n771), .A2(new_n344), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n776), .B2(G303), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n821), .A2(new_n825), .A3(new_n781), .A4(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n787), .A2(G143), .B1(G159), .B2(new_n765), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  INV_X1    g0630(.A(G150), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n830), .B2(new_n792), .C1(new_n831), .C2(new_n768), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n285), .B1(new_n820), .B2(G132), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n214), .B2(new_n771), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n773), .A2(new_n202), .B1(new_n213), .B2(new_n779), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n832), .B2(new_n833), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n828), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n759), .ZN(new_n841));
  INV_X1    g0641(.A(new_n744), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n759), .A2(new_n756), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT97), .Z(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n842), .B1(new_n845), .B2(new_n316), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n841), .B(new_n846), .C1(new_n815), .C2(new_n757), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n818), .A2(new_n847), .ZN(G384));
  INV_X1    g0648(.A(KEYINPUT35), .ZN(new_n849));
  OAI211_X1 g0649(.A(G116), .B(new_n219), .C1(new_n609), .C2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n849), .B2(new_n609), .ZN(new_n851));
  XOR2_X1   g0651(.A(KEYINPUT98), .B(KEYINPUT36), .Z(new_n852));
  XNOR2_X1  g0652(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n217), .A2(G77), .A3(new_n359), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n202), .A2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n206), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n376), .A2(new_n314), .A3(new_n371), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n331), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(new_n392), .A3(new_n393), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n383), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT100), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT99), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n860), .A2(new_n864), .A3(new_n669), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n247), .B1(new_n374), .B2(new_n375), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n330), .B1(new_n866), .B2(new_n371), .ZN(new_n867));
  INV_X1    g0667(.A(new_n669), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT99), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT100), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n383), .A2(new_n861), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n863), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n396), .A2(new_n669), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n876), .A3(new_n383), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT101), .B1(new_n388), .B2(new_n394), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT101), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n396), .A2(new_n399), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n874), .A2(KEYINPUT37), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n870), .B1(new_n385), .B2(new_n402), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n858), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n870), .B1(KEYINPUT100), .B2(new_n862), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n876), .B1(new_n887), .B2(new_n873), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n879), .A2(new_n881), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(new_n877), .ZN(new_n890));
  OAI211_X1 g0690(.A(KEYINPUT38), .B(new_n884), .C1(new_n888), .C2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  INV_X1    g0693(.A(new_n435), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(new_n670), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n442), .B2(new_n424), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n623), .A2(new_n895), .ZN(new_n897));
  INV_X1    g0697(.A(new_n423), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n420), .B2(new_n421), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n899), .B2(new_n894), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n734), .A2(new_n893), .A3(new_n815), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n734), .A2(new_n815), .A3(new_n901), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n875), .B(new_n383), .C1(new_n388), .C2(new_n394), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n878), .A2(new_n882), .B1(new_n904), .B2(KEYINPUT37), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n395), .A2(new_n401), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n383), .B(KEYINPUT17), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n875), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n858), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n903), .B1(new_n891), .B2(new_n909), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n892), .A2(new_n902), .B1(new_n910), .B2(new_n893), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT103), .Z(new_n912));
  NAND2_X1  g0712(.A1(new_n445), .A2(new_n734), .ZN(new_n913));
  OAI21_X1  g0713(.A(G330), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n913), .B2(new_n912), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT102), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n661), .A2(new_n697), .A3(new_n670), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n702), .A2(new_n670), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT29), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n916), .B1(new_n920), .B2(new_n445), .ZN(new_n921));
  AOI211_X1 g0721(.A(KEYINPUT102), .B(new_n444), .C1(new_n917), .C2(new_n919), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n628), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n891), .A2(new_n909), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n436), .A2(new_n681), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n886), .A2(KEYINPUT39), .A3(new_n891), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n661), .A2(new_n670), .A3(new_n815), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n813), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n886), .A2(new_n891), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n932), .A3(new_n901), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n402), .A2(new_n868), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n929), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n923), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n915), .A2(new_n937), .B1(new_n206), .B2(new_n741), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n915), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n857), .B1(new_n938), .B2(new_n939), .ZN(G367));
  NAND2_X1  g0740(.A1(new_n751), .A2(new_n237), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n941), .B(new_n760), .C1(new_n210), .C2(new_n312), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n744), .B1(new_n942), .B2(KEYINPUT107), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(KEYINPUT107), .B2(new_n942), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT108), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n771), .A2(new_n529), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n287), .B1(new_n820), .B2(G317), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n766), .B2(new_n801), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n946), .B(new_n948), .C1(G107), .C2(new_n796), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n822), .A2(new_n790), .B1(new_n823), .B2(new_n768), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G311), .B2(new_n776), .ZN(new_n951));
  INV_X1    g0751(.A(new_n773), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(G116), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT46), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n949), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n773), .A2(new_n213), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n771), .A2(new_n316), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(G150), .C2(new_n787), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n780), .A2(G68), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n287), .B1(new_n782), .B2(new_n830), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n765), .B2(G50), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n776), .A2(G143), .B1(G159), .B2(new_n767), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n958), .A2(new_n959), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n955), .A2(KEYINPUT47), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT47), .B1(new_n955), .B2(new_n963), .ZN(new_n965));
  INV_X1    g0765(.A(new_n759), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n945), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n535), .A2(new_n536), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n681), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n642), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n658), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n968), .B1(new_n807), .B2(new_n972), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n617), .B(new_n619), .C1(new_n611), .C2(new_n670), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n656), .A2(new_n600), .A3(new_n681), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n686), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT44), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n686), .A2(new_n980), .A3(new_n976), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n686), .B2(new_n976), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n684), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(new_n684), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n673), .A2(G330), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n679), .A2(new_n685), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n683), .B2(new_n685), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n673), .A3(G330), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(new_n736), .A3(new_n708), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n988), .A2(new_n996), .A3(KEYINPUT105), .ZN(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT105), .B1(new_n988), .B2(new_n996), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n738), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n691), .B(KEYINPUT41), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(KEYINPUT106), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT106), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n737), .B1(new_n997), .B2(new_n998), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n1005), .B2(new_n1001), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n743), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n990), .B1(new_n974), .B2(new_n975), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT42), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n617), .B1(new_n974), .B2(new_n512), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n670), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1009), .A2(new_n1011), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n684), .B1(new_n974), .B2(new_n975), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1014), .B(new_n1015), .Z(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n973), .B1(new_n1007), .B2(new_n1017), .ZN(G387));
  NAND2_X1  g0818(.A1(new_n995), .A2(new_n743), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n234), .A2(new_n448), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1020), .A2(new_n751), .B1(new_n689), .B2(new_n747), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n248), .A2(G50), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT50), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n448), .B1(new_n214), .B2(new_n316), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1024), .B(new_n689), .C1(new_n1023), .C2(new_n1022), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1021), .A2(new_n1025), .B1(G107), .B2(new_n210), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n842), .B1(new_n1026), .B2(new_n760), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n285), .B(new_n946), .C1(G150), .C2(new_n820), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n202), .B2(new_n822), .C1(new_n248), .C2(new_n768), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n780), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1030), .A2(new_n312), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n776), .A2(G159), .B1(G68), .B2(new_n765), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n316), .B2(new_n773), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n771), .A2(new_n550), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n285), .B1(new_n782), .B2(new_n793), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n952), .A2(G294), .B1(new_n796), .B2(G283), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(KEYINPUT109), .B(G322), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G317), .A2(new_n787), .B1(new_n776), .B2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G303), .A2(new_n765), .B1(new_n767), .B2(G311), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1037), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1035), .B(new_n1036), .C1(new_n1044), .C2(KEYINPUT49), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(KEYINPUT49), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1034), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1027), .B1(new_n1047), .B2(new_n966), .C1(new_n683), .C2(new_n807), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n738), .A2(new_n995), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n996), .A2(new_n691), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1019), .B(new_n1048), .C1(new_n1049), .C2(new_n1050), .ZN(G393));
  NAND3_X1  g0851(.A1(new_n986), .A2(new_n743), .A3(new_n987), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n760), .B1(new_n529), .B2(new_n210), .C1(new_n752), .C2(new_n244), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n744), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G311), .A2(new_n787), .B1(new_n776), .B2(G317), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  AOI211_X1 g0856(.A(new_n287), .B(new_n772), .C1(new_n820), .C2(new_n1038), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n801), .C2(new_n773), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n767), .A2(G303), .B1(G116), .B2(new_n796), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n823), .B2(new_n766), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT110), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G150), .A2(new_n776), .B1(new_n787), .B2(G159), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT51), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n285), .B(new_n826), .C1(G143), .C2(new_n820), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n780), .A2(G77), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n952), .A2(G68), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n328), .A2(new_n765), .B1(new_n767), .B2(G50), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1058), .A2(new_n1061), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1054), .B1(new_n1069), .B2(new_n759), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n976), .B2(new_n807), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT111), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n693), .B1(new_n988), .B2(new_n996), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n999), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1072), .B1(new_n999), .B2(new_n1073), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1052), .B(new_n1071), .C1(new_n1074), .C2(new_n1075), .ZN(G390));
  NAND4_X1  g0876(.A1(new_n726), .A2(new_n735), .A3(new_n815), .A4(new_n901), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n701), .A2(new_n643), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n700), .A2(new_n698), .A3(new_n658), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n670), .B(new_n812), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n813), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n901), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n927), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n924), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT39), .B1(new_n891), .B2(new_n909), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n892), .B2(KEYINPUT39), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n927), .B1(new_n931), .B2(new_n901), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1077), .B(new_n1084), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n924), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n813), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n707), .B2(new_n815), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n901), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1083), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n926), .A2(new_n928), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1089), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n734), .A2(G330), .A3(new_n815), .A4(new_n901), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT112), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n721), .A2(new_n723), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n814), .B1(new_n1098), .B2(new_n731), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT112), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1099), .A2(new_n1100), .A3(G330), .A4(new_n901), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1088), .B(new_n743), .C1(new_n1095), .C2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(KEYINPUT113), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n931), .A2(new_n901), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1106), .A2(new_n1083), .B1(new_n926), .B2(new_n928), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1105), .B1(new_n1107), .B2(new_n1089), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT113), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n1088), .A4(new_n743), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1077), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1112), .B(new_n1089), .C1(new_n1094), .C2(new_n1093), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1102), .B1(new_n1114), .B2(new_n1084), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n734), .A2(G330), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n444), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n628), .B(new_n1118), .C1(new_n921), .C2(new_n922), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n734), .A2(G330), .A3(new_n815), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1081), .B1(new_n1092), .B2(new_n1120), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1077), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n726), .A2(new_n735), .A3(new_n815), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1092), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1102), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1122), .B1(new_n1125), .B2(new_n931), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1113), .A2(new_n1115), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT102), .B1(new_n708), .B2(new_n444), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n920), .A2(new_n916), .A3(new_n445), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n627), .B(new_n1117), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1077), .A2(new_n1121), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1105), .B1(new_n1092), .B2(new_n1123), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n1091), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1108), .A2(new_n1130), .A3(new_n1133), .A4(new_n1088), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1127), .A2(new_n1134), .A3(new_n691), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n744), .B1(new_n844), .B2(new_n328), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n822), .A2(new_n550), .B1(new_n529), .B2(new_n766), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n792), .A2(new_n801), .B1(new_n489), .B2(new_n768), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n214), .B2(new_n771), .C1(new_n823), .C2(new_n782), .ZN(new_n1140));
  OR3_X1    g0940(.A1(new_n774), .A2(KEYINPUT114), .A3(new_n287), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT114), .B1(new_n774), .B2(new_n287), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1065), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n768), .A2(new_n830), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n285), .B(new_n1144), .C1(G125), .C2(new_n820), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n787), .A2(G132), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT54), .B(G143), .Z(new_n1147));
  NAND2_X1  g0947(.A1(new_n765), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n771), .A2(new_n202), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n776), .B2(G128), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n773), .A2(new_n831), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n783), .B2(new_n1030), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1140), .A2(new_n1143), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1136), .B1(new_n1155), .B2(new_n759), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1086), .B2(new_n757), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1111), .A2(new_n1135), .A3(new_n1157), .ZN(G378));
  OAI21_X1  g0958(.A(new_n669), .B1(new_n253), .B2(new_n258), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n303), .B(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n756), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n759), .A2(G50), .A3(new_n756), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n792), .A2(new_n550), .B1(new_n529), .B2(new_n768), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n822), .A2(new_n489), .B1(new_n312), .B2(new_n766), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n281), .A2(new_n446), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n284), .B(new_n1167), .C1(new_n820), .C2(G283), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n316), .B2(new_n773), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1165), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n771), .A2(new_n213), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT115), .Z(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n959), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1173), .A2(new_n1174), .B1(new_n202), .B2(new_n1167), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n780), .A2(G150), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n776), .A2(G125), .B1(G137), .B2(new_n765), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G132), .A2(new_n767), .B1(new_n952), .B2(new_n1147), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n787), .A2(G128), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT59), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G33), .B(G41), .C1(new_n820), .C2(G124), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n783), .B2(new_n771), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1175), .B1(new_n1174), .B2(new_n1173), .C1(new_n1181), .C2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n842), .B(new_n1164), .C1(new_n1184), .C2(new_n759), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1163), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1162), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n911), .B2(G330), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n903), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n893), .B1(new_n924), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n902), .B1(new_n886), .B2(new_n891), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1188), .B(G330), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n935), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n935), .ZN(new_n1196));
  OAI21_X1  g0996(.A(G330), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1162), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1198), .A3(new_n1193), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1187), .B1(new_n1200), .B2(new_n743), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1134), .A2(new_n1130), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n691), .B1(new_n1202), .B2(KEYINPUT57), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1088), .B1(new_n1095), .B2(new_n1102), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1130), .B1(new_n1204), .B2(new_n1126), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1200), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1201), .B1(new_n1203), .B2(new_n1208), .ZN(G375));
  XOR2_X1   g1009(.A(new_n742), .B(KEYINPUT116), .Z(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1092), .A2(new_n756), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n844), .A2(G68), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n766), .A2(new_n831), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n285), .B(new_n1214), .C1(G128), .C2(new_n820), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n787), .A2(G137), .B1(new_n767), .B2(new_n1147), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n783), .C2(new_n773), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n776), .A2(G132), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT117), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n1172), .C1(new_n202), .C2(new_n1030), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n768), .A2(new_n550), .B1(new_n529), .B2(new_n773), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G107), .B2(new_n765), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n287), .B(new_n957), .C1(G303), .C2(new_n820), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G283), .A2(new_n787), .B1(new_n776), .B2(G294), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1217), .A2(new_n1220), .B1(new_n1031), .B2(new_n1225), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n842), .B(new_n1213), .C1(new_n1226), .C2(new_n759), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1133), .A2(new_n1211), .B1(new_n1212), .B2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1002), .B1(new_n1126), .B2(new_n1119), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(G381));
  OR2_X1    g1031(.A1(G375), .A2(G378), .ZN(new_n1232));
  OR4_X1    g1032(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G387), .A2(new_n1232), .A3(new_n1233), .A4(G381), .ZN(G407));
  OAI211_X1 g1034(.A(G407), .B(G213), .C1(G343), .C2(new_n1232), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT118), .ZN(G409));
  XNOR2_X1  g1036(.A(G393), .B(new_n809), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT123), .ZN(new_n1239));
  INV_X1    g1039(.A(G390), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G387), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n973), .B(G390), .C1(new_n1007), .C2(new_n1017), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT124), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1239), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AOI211_X1 g1045(.A(KEYINPUT123), .B(KEYINPUT124), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1238), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT106), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1005), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n742), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1016), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G390), .B1(new_n1251), .B2(new_n973), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1242), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1244), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT123), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1243), .A2(new_n1239), .A3(new_n1244), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1237), .A3(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1247), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT120), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1228), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n691), .B1(new_n1126), .B2(new_n1119), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT119), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1261), .B1(new_n1263), .B2(KEYINPUT60), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT119), .B1(new_n1126), .B2(new_n1119), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1260), .B1(new_n1264), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1259), .B1(new_n1268), .B2(G384), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n693), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1263), .A2(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1228), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(G384), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(KEYINPUT120), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1268), .A2(G384), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1269), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT121), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(G213), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(G343), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1205), .A2(new_n1002), .A3(new_n1200), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1187), .B1(new_n1200), .B2(new_n1211), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1282), .B1(new_n1285), .B2(G378), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(G375), .B2(G378), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1269), .A2(new_n1275), .A3(KEYINPUT121), .A4(new_n1276), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1279), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1289), .B(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1281), .A2(G2897), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1279), .A2(new_n1292), .A3(new_n1288), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1287), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1277), .A2(G2897), .A3(new_n1281), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(KEYINPUT125), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1291), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT125), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1258), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT122), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT122), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1293), .A2(new_n1304), .A3(new_n1295), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1294), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1247), .A2(new_n1257), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1289), .B(KEYINPUT63), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1297), .A4(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1301), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT126), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1301), .A2(new_n1312), .A3(new_n1309), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(G405));
  XNOR2_X1  g1114(.A(G375), .B(G378), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1277), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1316), .B(KEYINPUT127), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1279), .A2(new_n1288), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1318), .B2(new_n1315), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(new_n1258), .ZN(G402));
endmodule


