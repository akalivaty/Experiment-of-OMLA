//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n642, new_n643, new_n645, new_n646, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1240, new_n1241, new_n1242;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  OR4_X1    g028(.A1(G235), .A2(G238), .A3(G236), .A4(G237), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n457), .A2(KEYINPUT69), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(KEYINPUT69), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n453), .A2(G2106), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n467), .A2(KEYINPUT70), .A3(G101), .A4(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n466), .A2(G137), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n466), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n465), .A2(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n463), .B2(new_n464), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n487), .B(new_n490), .C1(new_n464), .C2(new_n463), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n463), .B2(new_n464), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n467), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n500), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n492), .A2(new_n499), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G62), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(KEYINPUT73), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n514), .A2(new_n517), .A3(G62), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n511), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT72), .A2(G651), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  AND3_X1   g102(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT6), .B1(KEYINPUT72), .B2(G651), .ZN(new_n529));
  AND2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n526), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n519), .A2(new_n533), .ZN(G166));
  NAND3_X1  g109(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n530), .A2(new_n531), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT74), .ZN(new_n537));
  INV_X1    g112(.A(G63), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n541), .B1(new_n528), .B2(new_n529), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n523), .A2(KEYINPUT75), .A3(new_n524), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(new_n543), .A3(G543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT76), .B(G51), .Z(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n532), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT7), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n548), .A2(G89), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n540), .A2(new_n547), .A3(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n544), .A2(new_n554), .B1(new_n555), .B2(new_n532), .ZN(new_n556));
  NAND2_X1  g131(.A1(G77), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G64), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n537), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n556), .B1(new_n559), .B2(G651), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT77), .ZN(G171));
  AOI22_X1  g136(.A1(new_n545), .A2(G43), .B1(G81), .B2(new_n548), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n514), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(KEYINPUT74), .B1(new_n512), .B2(new_n513), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G56), .ZN(new_n568));
  NAND2_X1  g143(.A1(G68), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n511), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  NAND4_X1  g147(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  INV_X1    g151(.A(G78), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT79), .B1(new_n577), .B2(new_n520), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n579), .A2(G78), .A3(G543), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n514), .A2(G65), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n511), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n580), .ZN(new_n584));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n536), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT80), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n583), .A2(new_n587), .B1(G91), .B2(new_n548), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n523), .A2(new_n524), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n520), .B1(new_n589), .B2(new_n541), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT9), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n590), .A2(new_n591), .A3(G53), .A4(new_n543), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n542), .A2(new_n543), .A3(G53), .A4(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT9), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n595), .B1(new_n592), .B2(new_n594), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n588), .B1(new_n596), .B2(new_n597), .ZN(G299));
  NOR2_X1   g173(.A1(new_n560), .A2(KEYINPUT77), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n600));
  AOI211_X1 g175(.A(new_n600), .B(new_n556), .C1(new_n559), .C2(G651), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n599), .A2(new_n601), .ZN(G301));
  INV_X1    g177(.A(G166), .ZN(G303));
  INV_X1    g178(.A(G74), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n565), .B2(new_n566), .ZN(new_n605));
  INV_X1    g180(.A(G87), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT81), .B1(new_n532), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n589), .A2(new_n514), .A3(new_n608), .A4(G87), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n605), .A2(G651), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n545), .A2(G49), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(G288));
  AOI22_X1  g187(.A1(new_n548), .A2(G86), .B1(G48), .B2(new_n525), .ZN(new_n613));
  OAI21_X1  g188(.A(G61), .B1(new_n530), .B2(new_n531), .ZN(new_n614));
  NAND2_X1  g189(.A1(G73), .A2(G543), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n511), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI211_X1 g193(.A(KEYINPUT82), .B(new_n511), .C1(new_n614), .C2(new_n615), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(new_n618), .B2(new_n619), .ZN(G305));
  AOI22_X1  g195(.A1(new_n545), .A2(G47), .B1(G85), .B2(new_n548), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n567), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n511), .ZN(G290));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n624));
  INV_X1    g199(.A(G92), .ZN(new_n625));
  OAI21_X1  g200(.A(KEYINPUT83), .B1(new_n532), .B2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  NOR3_X1   g202(.A1(new_n532), .A2(KEYINPUT83), .A3(new_n625), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n626), .ZN(new_n631));
  NAND2_X1  g206(.A1(G79), .A2(G543), .ZN(new_n632));
  INV_X1    g207(.A(G66), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n536), .B2(new_n633), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n545), .A2(G54), .B1(G651), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n629), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g213(.A(new_n637), .B1(G171), .B2(G868), .ZN(G321));
  MUX2_X1   g214(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g215(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g216(.A(new_n636), .ZN(new_n642));
  INV_X1    g217(.A(G559), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(G860), .ZN(G148));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G868), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(G868), .B2(new_n571), .ZN(G323));
  XNOR2_X1  g222(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n648));
  XNOR2_X1  g223(.A(G323), .B(new_n648), .ZN(G282));
  NAND2_X1  g224(.A1(new_n466), .A2(G135), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n480), .A2(G123), .ZN(new_n651));
  OR2_X1    g226(.A1(G99), .A2(G2105), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n652), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT12), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT85), .B(KEYINPUT13), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G2100), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(G2100), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n655), .A2(new_n660), .A3(new_n661), .ZN(G156));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2427), .B(G2430), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT15), .B(G2435), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2438), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT14), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n666), .A2(new_n668), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1341), .B(G1348), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  AND3_X1   g249(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n671), .B2(new_n672), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2451), .B(G2454), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2443), .B(G2446), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n677), .A2(new_n681), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n664), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n684), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n663), .A3(new_n682), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n685), .A2(new_n687), .A3(G14), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(KEYINPUT89), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n690));
  NAND4_X1  g265(.A1(new_n685), .A2(new_n687), .A3(new_n690), .A4(G14), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(G401));
  XOR2_X1   g267(.A(G2084), .B(G2090), .Z(new_n693));
  XNOR2_X1  g268(.A(G2072), .B(G2078), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  XNOR2_X1  g270(.A(G2067), .B(G2678), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n693), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(KEYINPUT17), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n697), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT91), .Z(new_n701));
  INV_X1    g276(.A(new_n693), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n695), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT18), .Z(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(new_n696), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n704), .B1(new_n699), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G2096), .B(G2100), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(G227));
  XOR2_X1   g284(.A(G1971), .B(G1976), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT19), .ZN(new_n711));
  XOR2_X1   g286(.A(G1956), .B(G2474), .Z(new_n712));
  XOR2_X1   g287(.A(G1961), .B(G1966), .Z(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n712), .A2(new_n713), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(new_n719), .B(new_n718), .S(new_n711), .Z(new_n720));
  NOR2_X1   g295(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(G1991), .B(G1996), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(G1981), .B(G1986), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(G229));
  NAND2_X1  g304(.A1(G171), .A2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n730), .B(new_n731), .C1(G5), .C2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  NOR2_X1   g308(.A1(G301), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G5), .A2(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(G1961), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n477), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  AND2_X1   g315(.A1(KEYINPUT24), .A2(G34), .ZN(new_n741));
  NOR2_X1   g316(.A1(KEYINPUT24), .A2(G34), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n738), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT96), .Z(new_n744));
  OR3_X1    g319(.A1(new_n739), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n740), .B1(new_n739), .B2(new_n744), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n654), .A2(new_n738), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT30), .B(G28), .ZN(new_n748));
  OR2_X1    g323(.A1(KEYINPUT31), .A2(G11), .ZN(new_n749));
  NAND2_X1  g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n748), .A2(new_n738), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n738), .A2(G33), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n466), .A2(G139), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(G115), .A2(G2104), .ZN(new_n759));
  INV_X1    g334(.A(G127), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n465), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G2105), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n753), .B1(new_n764), .B2(new_n738), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2072), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT99), .B(G2078), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n509), .A2(G29), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n738), .A2(G27), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n768), .A2(new_n769), .A3(new_n767), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n752), .A2(new_n766), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n738), .A2(G32), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n466), .A2(G141), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT26), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n777), .B(new_n779), .C1(G129), .C2(new_n480), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT98), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n776), .A2(KEYINPUT98), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n774), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  INV_X1    g362(.A(G1966), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n733), .A2(G21), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G286), .B2(G16), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n783), .A2(new_n784), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n773), .B1(new_n793), .B2(new_n738), .ZN(new_n794));
  INV_X1    g369(.A(new_n787), .ZN(new_n795));
  INV_X1    g370(.A(new_n791), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n794), .A2(new_n795), .B1(G1966), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n737), .A2(new_n772), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(KEYINPUT100), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n794), .A2(new_n795), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(G1966), .ZN(new_n801));
  AND3_X1   g376(.A1(new_n792), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT100), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n802), .A2(new_n803), .A3(new_n737), .A4(new_n772), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n738), .A2(G35), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n484), .B2(G29), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT29), .ZN(new_n807));
  INV_X1    g382(.A(G2090), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT101), .ZN(new_n810));
  NOR2_X1   g385(.A1(G4), .A2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT94), .Z(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n636), .B2(new_n733), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1348), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n733), .A2(G19), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n571), .B2(new_n733), .ZN(new_n816));
  INV_X1    g391(.A(G1341), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n738), .A2(G26), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT28), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n466), .A2(G140), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n480), .A2(G128), .ZN(new_n823));
  OR2_X1    g398(.A1(G104), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT95), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n821), .B1(new_n827), .B2(G29), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(G2067), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(G2067), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n829), .A2(new_n830), .B1(new_n808), .B2(new_n807), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n810), .A2(new_n814), .A3(new_n818), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n733), .A2(G20), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT23), .Z(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G299), .B2(G16), .ZN(new_n835));
  INV_X1    g410(.A(G1956), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n799), .A2(new_n804), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT34), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n733), .A2(G22), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G166), .B2(new_n733), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G1971), .ZN(new_n843));
  NAND2_X1  g418(.A1(G305), .A2(G16), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT32), .B(G1981), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n733), .A2(G6), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n846), .ZN(new_n848));
  INV_X1    g423(.A(new_n845), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n843), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT92), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n733), .A2(G23), .ZN(new_n853));
  INV_X1    g428(.A(G288), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n854), .B2(new_n733), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT33), .B(G1976), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n851), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n852), .B1(new_n851), .B2(new_n857), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n840), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n851), .A2(new_n857), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT92), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n863), .A2(KEYINPUT34), .A3(new_n858), .ZN(new_n864));
  MUX2_X1   g439(.A(G24), .B(G290), .S(G16), .Z(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(G1986), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(G1986), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n738), .A2(G25), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n466), .A2(G131), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n480), .A2(G119), .ZN(new_n870));
  OR2_X1    g445(.A1(G95), .A2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n868), .B1(new_n874), .B2(new_n738), .ZN(new_n875));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G1991), .Z(new_n876));
  XOR2_X1   g451(.A(new_n875), .B(new_n876), .Z(new_n877));
  NOR3_X1   g452(.A1(new_n866), .A2(new_n867), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n861), .A2(new_n864), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n880));
  NOR2_X1   g455(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n839), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n861), .A2(new_n864), .A3(new_n880), .A4(new_n878), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(G311));
  NAND2_X1  g460(.A1(new_n879), .A2(new_n882), .ZN(new_n886));
  INV_X1    g461(.A(new_n839), .ZN(new_n887));
  AND4_X1   g462(.A1(KEYINPUT102), .A2(new_n886), .A3(new_n884), .A4(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT102), .B1(new_n883), .B2(new_n884), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(G150));
  NAND2_X1  g465(.A1(new_n567), .A2(G67), .ZN(new_n891));
  NAND2_X1  g466(.A1(G80), .A2(G543), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n511), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G55), .ZN(new_n894));
  INV_X1    g469(.A(G93), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n544), .A2(new_n894), .B1(new_n895), .B2(new_n532), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G860), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT37), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n642), .A2(G559), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT38), .ZN(new_n902));
  INV_X1    g477(.A(new_n570), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n891), .A2(new_n892), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G651), .ZN(new_n905));
  INV_X1    g480(.A(new_n896), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n903), .A2(new_n905), .A3(new_n562), .A4(new_n906), .ZN(new_n907));
  OAI22_X1  g482(.A1(new_n570), .A2(new_n563), .B1(new_n893), .B2(new_n896), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n902), .B(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT39), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT103), .Z(new_n913));
  OAI21_X1  g488(.A(new_n898), .B1(new_n911), .B2(KEYINPUT39), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n900), .B1(new_n913), .B2(new_n914), .ZN(G145));
  XNOR2_X1  g490(.A(new_n484), .B(new_n654), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(new_n477), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n785), .A2(new_n827), .ZN(new_n918));
  INV_X1    g493(.A(new_n827), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(new_n783), .A3(new_n784), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n918), .A2(new_n920), .A3(new_n763), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n763), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  INV_X1    g497(.A(new_n491), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT3), .B(G2104), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n490), .B1(new_n924), .B2(new_n487), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT104), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n496), .A2(new_n498), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n489), .A2(new_n929), .A3(new_n491), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n921), .A2(new_n922), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n931), .ZN(new_n933));
  INV_X1    g508(.A(new_n920), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n919), .B1(new_n783), .B2(new_n784), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n764), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n918), .A2(new_n920), .A3(new_n763), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n466), .A2(G142), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n480), .A2(G130), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n467), .A2(G118), .ZN(new_n942));
  OAI21_X1  g517(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n940), .B(new_n941), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(new_n657), .Z(new_n945));
  OR2_X1    g520(.A1(new_n945), .A2(new_n873), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n873), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n917), .B1(new_n939), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n946), .A2(KEYINPUT105), .A3(new_n947), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n932), .B2(new_n938), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n931), .B1(new_n921), .B2(new_n922), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n936), .A2(new_n933), .A3(new_n937), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n952), .A2(new_n953), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT106), .B1(new_n961), .B2(new_n917), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n963));
  INV_X1    g538(.A(new_n917), .ZN(new_n964));
  AOI211_X1 g539(.A(new_n963), .B(new_n964), .C1(new_n955), .C2(new_n960), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n956), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g542(.A(G299), .B(new_n642), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(KEYINPUT41), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(KEYINPUT41), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n909), .B(new_n645), .Z(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n968), .B2(new_n972), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT42), .ZN(new_n975));
  XNOR2_X1  g550(.A(G290), .B(G166), .ZN(new_n976));
  XNOR2_X1  g551(.A(G288), .B(G305), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n976), .B(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n973), .B(new_n979), .C1(new_n968), .C2(new_n972), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n975), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n978), .B1(new_n975), .B2(new_n980), .ZN(new_n982));
  OAI21_X1  g557(.A(G868), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(G868), .B2(new_n897), .ZN(G295));
  OAI21_X1  g559(.A(new_n983), .B1(G868), .B2(new_n897), .ZN(G331));
  NAND2_X1  g560(.A1(new_n909), .A2(G301), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n907), .B(new_n908), .C1(new_n599), .C2(new_n601), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n986), .A2(G168), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(G168), .B1(new_n986), .B2(new_n987), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n969), .B(new_n970), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n989), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n986), .A2(G168), .A3(new_n987), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n968), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT108), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n990), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n978), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n999));
  INV_X1    g574(.A(new_n978), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n990), .A2(new_n993), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G37), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(new_n999), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n994), .A2(new_n978), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1004), .B(KEYINPUT44), .C1(new_n1006), .C2(new_n999), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n999), .B1(new_n998), .B2(new_n1003), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1003), .A2(new_n999), .A3(new_n1005), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n1011));
  OAI21_X1  g586(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(G397));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n931), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n472), .A2(new_n476), .A3(G40), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1996), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n785), .B(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n827), .B(G2067), .Z(new_n1021));
  NAND2_X1  g596(.A1(new_n874), .A2(new_n876), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n874), .A2(new_n876), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(G290), .B(G1986), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1018), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n605), .A2(G651), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n607), .A2(new_n609), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1027), .A2(new_n611), .A3(G1976), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT114), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n472), .A2(new_n476), .A3(G40), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(new_n1013), .A3(new_n931), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n610), .A2(new_n1033), .A3(G1976), .A4(new_n611), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1030), .A2(new_n1032), .A3(G8), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n613), .B(new_n1039), .C1(new_n618), .C2(new_n619), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n525), .A2(G48), .ZN(new_n1041));
  INV_X1    g616(.A(G86), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(new_n532), .ZN(new_n1043));
  OAI21_X1  g618(.A(G1981), .B1(new_n1043), .B2(new_n616), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1040), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1048), .A2(new_n1032), .A3(G8), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1036), .A2(new_n1038), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1035), .A2(KEYINPUT52), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n509), .A2(new_n1013), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(KEYINPUT50), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n489), .A2(new_n491), .B1(new_n927), .B2(new_n500), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1384), .B1(new_n1058), .B2(new_n499), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(KEYINPUT117), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT110), .B(G2090), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1017), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1971), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1015), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1031), .B1(new_n1059), .B2(new_n1067), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n931), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1054), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1072));
  AND2_X1   g647(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1073));
  OAI221_X1 g648(.A(G8), .B1(new_n1072), .B2(new_n1073), .C1(new_n519), .C2(new_n533), .ZN(new_n1074));
  NOR2_X1   g649(.A1(G166), .A2(new_n1054), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(new_n1073), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1052), .B(new_n1053), .C1(new_n1071), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1031), .A2(new_n1063), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1014), .A2(new_n1060), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n509), .A2(KEYINPUT50), .A3(new_n1013), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1017), .B1(new_n1056), .B2(new_n1015), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n931), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1971), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1079), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT50), .B1(new_n931), .B2(new_n1013), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1082), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1031), .B(new_n1063), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1070), .A2(KEYINPUT111), .A3(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1087), .A2(new_n1091), .A3(G8), .A4(new_n1076), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1078), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT126), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1054), .B1(new_n1098), .B2(KEYINPUT111), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1099), .A2(KEYINPUT113), .A3(new_n1076), .A4(new_n1087), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT126), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n1078), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n740), .B(new_n1031), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1031), .B1(new_n1056), .B2(new_n1015), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT45), .B1(new_n931), .B2(new_n1013), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n788), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1108), .A3(G168), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G8), .ZN(new_n1110));
  AOI21_X1  g685(.A(G168), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT51), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1113), .A3(G8), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1116), .A2(G2078), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1031), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1117), .A2(new_n1118), .B1(new_n731), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1118), .A2(G2078), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  OR2_X1    g699(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1125));
  NAND2_X1  g700(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1016), .A2(new_n1085), .A3(new_n1031), .A4(new_n1122), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1120), .A2(new_n1125), .A3(new_n1126), .A4(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1115), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1097), .A2(new_n1104), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(KEYINPUT123), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1032), .A2(G2067), .ZN(new_n1136));
  INV_X1    g711(.A(G1348), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1136), .B1(new_n1119), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1138), .B2(new_n636), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT57), .B(new_n588), .C1(new_n596), .C2(new_n597), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n583), .A2(new_n587), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n548), .A2(G91), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n592), .A2(new_n594), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1140), .A2(new_n1141), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1141), .B1(new_n1140), .B2(new_n1147), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1116), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(G2072), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1152), .A2(new_n836), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1139), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1152), .A2(new_n836), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1160), .A2(new_n1150), .A3(new_n1135), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1138), .A2(new_n636), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1160), .B2(new_n1150), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n927), .B1(new_n492), .B2(KEYINPUT104), .ZN(new_n1166));
  AOI21_X1  g741(.A(G1384), .B1(new_n1166), .B2(new_n930), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1082), .B1(new_n1167), .B2(KEYINPUT50), .ZN(new_n1168));
  AOI21_X1  g743(.A(G1348), .B1(new_n1168), .B2(new_n1031), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1165), .B1(new_n1169), .B2(new_n1136), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1119), .A2(new_n1137), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1136), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1165), .B1(new_n642), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n642), .A2(new_n1173), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1170), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .A4(new_n1176), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1056), .A2(new_n1015), .ZN(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT121), .B(G1996), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1181), .A2(new_n1085), .A3(new_n1031), .A4(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(new_n817), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1032), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1180), .B1(new_n1187), .B2(new_n571), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n903), .A2(new_n562), .ZN(new_n1189));
  AOI211_X1 g764(.A(KEYINPUT59), .B(new_n1189), .C1(new_n1183), .C2(new_n1186), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1179), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1164), .B1(new_n1178), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1162), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1133), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g771(.A(KEYINPUT125), .B(new_n1194), .C1(new_n1162), .C2(new_n1192), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1132), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1115), .A2(KEYINPUT62), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1112), .A2(new_n1200), .A3(new_n1114), .ZN(new_n1201));
  AOI21_X1  g776(.A(G301), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1097), .A2(new_n1104), .A3(new_n1199), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT63), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1207), .A2(G8), .A3(G168), .ZN(new_n1208));
  NOR3_X1   g783(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1099), .A2(new_n1087), .ZN(new_n1210));
  OAI211_X1 g785(.A(new_n1102), .B(new_n1209), .C1(new_n1076), .C2(new_n1210), .ZN(new_n1211));
  AOI211_X1 g786(.A(new_n1208), .B(new_n1077), .C1(new_n1101), .C2(new_n1100), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1211), .B1(new_n1212), .B2(KEYINPUT63), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1102), .A2(new_n1205), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1032), .A2(G8), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1216), .A2(new_n1037), .A3(new_n854), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1040), .B(KEYINPUT116), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1215), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1214), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1204), .A2(new_n1213), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1026), .B1(new_n1198), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1021), .A2(new_n793), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1224));
  OR2_X1    g799(.A1(new_n1224), .A2(KEYINPUT46), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1224), .A2(KEYINPUT46), .ZN(new_n1226));
  AOI22_X1  g801(.A1(new_n1018), .A2(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1227), .B(KEYINPUT47), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1229));
  OAI22_X1  g804(.A1(new_n1229), .A2(new_n1022), .B1(G2067), .B2(new_n827), .ZN(new_n1230));
  AND2_X1   g805(.A1(new_n1230), .A2(new_n1018), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1024), .A2(new_n1018), .ZN(new_n1232));
  XOR2_X1   g807(.A(new_n1232), .B(KEYINPUT127), .Z(new_n1233));
  NOR2_X1   g808(.A1(G290), .A2(G1986), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1018), .A2(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g810(.A(new_n1235), .B(KEYINPUT48), .ZN(new_n1236));
  AOI211_X1 g811(.A(new_n1228), .B(new_n1231), .C1(new_n1233), .C2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1222), .A2(new_n1237), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g813(.A1(G227), .A2(new_n461), .ZN(new_n1240));
  OAI21_X1  g814(.A(new_n1240), .B1(new_n727), .B2(new_n728), .ZN(new_n1241));
  AOI21_X1  g815(.A(new_n1241), .B1(new_n689), .B2(new_n691), .ZN(new_n1242));
  OAI211_X1 g816(.A(new_n966), .B(new_n1242), .C1(new_n1008), .C2(new_n1009), .ZN(G225));
  INV_X1    g817(.A(G225), .ZN(G308));
endmodule


