//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT16), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n191), .A2(KEYINPUT16), .A3(G140), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G146), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(G146), .B1(new_n193), .B2(new_n194), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G237), .ZN(new_n199));
  INV_X1    g013(.A(G953), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G214), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  OR2_X1    g016(.A1(KEYINPUT90), .A2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT90), .A2(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n204), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT17), .A3(G131), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(G131), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n211), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n198), .B(new_n209), .C1(new_n213), .C2(KEYINPUT17), .ZN(new_n214));
  XNOR2_X1  g028(.A(G113), .B(G122), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n215), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT93), .ZN(new_n218));
  XNOR2_X1  g032(.A(G125), .B(G140), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT92), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n190), .A2(new_n192), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT92), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G146), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT64), .B(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n219), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(KEYINPUT91), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G131), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n206), .A2(new_n207), .A3(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n208), .A2(G131), .A3(new_n229), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n218), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AND4_X1   g048(.A1(new_n218), .A2(new_n233), .A3(new_n231), .A4(new_n227), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n214), .B(new_n217), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n233), .A2(new_n231), .A3(new_n227), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT93), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n232), .A2(new_n218), .A3(new_n233), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n217), .B1(new_n241), .B2(new_n214), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n188), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G475), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n219), .B(KEYINPUT19), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n196), .B1(new_n245), .B2(new_n225), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n239), .A2(new_n240), .B1(new_n213), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n236), .B1(new_n247), .B2(new_n217), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT20), .ZN(new_n249));
  NOR2_X1   g063(.A1(G475), .A2(G902), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n249), .B1(new_n248), .B2(new_n250), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n244), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT71), .B(G902), .Z(new_n254));
  INV_X1    g068(.A(G107), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT80), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G107), .ZN(new_n258));
  INV_X1    g072(.A(G122), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G116), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G122), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n256), .A2(new_n258), .A3(new_n260), .A4(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT95), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G143), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n261), .A2(KEYINPUT14), .A3(G122), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n260), .A2(new_n262), .ZN(new_n273));
  OAI211_X1 g087(.A(G107), .B(new_n272), .C1(new_n273), .C2(KEYINPUT14), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n264), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n256), .A2(new_n258), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n273), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n277), .A2(new_n263), .B1(new_n270), .B2(new_n269), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT94), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT13), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n266), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n268), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n266), .A2(new_n280), .ZN(new_n283));
  OAI21_X1  g097(.A(G134), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n278), .A2(new_n279), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n279), .B1(new_n278), .B2(new_n284), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n275), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT9), .B(G234), .Z(new_n288));
  XNOR2_X1  g102(.A(new_n288), .B(KEYINPUT79), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(G217), .A3(new_n200), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n290), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n292), .B(new_n275), .C1(new_n285), .C2(new_n286), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n254), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G478), .ZN(new_n295));
  NOR2_X1   g109(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n294), .B(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n254), .ZN(new_n302));
  AOI211_X1 g116(.A(new_n200), .B(new_n302), .C1(G234), .C2(G237), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT21), .B(G898), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n200), .A2(G952), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(G234), .B2(G237), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n253), .A2(new_n301), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G210), .B1(G237), .B2(G902), .ZN(new_n312));
  OR3_X1    g126(.A1(new_n216), .A2(KEYINPUT82), .A3(G107), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT82), .B1(new_n216), .B2(G107), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT80), .B(G107), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(G104), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G101), .ZN(new_n317));
  XNOR2_X1  g131(.A(G116), .B(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT5), .ZN(new_n319));
  INV_X1    g133(.A(G113), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n261), .A2(G119), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT5), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT2), .B(G113), .Z(new_n324));
  AOI22_X1  g138(.A1(new_n319), .A2(new_n323), .B1(new_n324), .B2(new_n318), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT81), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(G104), .B2(new_n255), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n315), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(G101), .B1(new_n216), .B2(G107), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n326), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n256), .A3(new_n258), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(new_n216), .B2(G107), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n333), .A2(new_n326), .A3(new_n334), .A4(new_n331), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n317), .B(new_n325), .C1(new_n332), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT87), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n216), .A2(G107), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n333), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n341), .B2(G101), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n332), .B2(new_n336), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n339), .A3(G101), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n324), .B1(KEYINPUT68), .B2(new_n318), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT2), .B(G113), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT68), .ZN(new_n347));
  INV_X1    g161(.A(G119), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G116), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n346), .B(new_n347), .C1(new_n321), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n344), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n333), .A2(new_n334), .A3(new_n331), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT81), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n355), .A2(new_n335), .B1(G101), .B2(new_n316), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT87), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n325), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n338), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G110), .B(G122), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n338), .A2(new_n353), .A3(new_n358), .A4(new_n360), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(KEYINPUT6), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT64), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G146), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n367), .A3(G143), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n220), .A2(G143), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n267), .A2(KEYINPUT1), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(KEYINPUT1), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G128), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n220), .A2(G143), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n225), .B2(G143), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT88), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n191), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n267), .B1(new_n368), .B2(KEYINPUT1), .ZN(new_n381));
  INV_X1    g195(.A(new_n375), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n365), .A2(new_n367), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n382), .B1(new_n383), .B2(new_n265), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n380), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT88), .B1(new_n385), .B2(G125), .ZN(new_n386));
  AND2_X1   g200(.A1(KEYINPUT0), .A2(G128), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n368), .A2(new_n370), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT65), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n368), .A2(KEYINPUT65), .A3(new_n370), .A4(new_n387), .ZN(new_n391));
  NOR2_X1   g205(.A1(KEYINPUT0), .A2(G128), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n390), .A2(new_n391), .B1(new_n376), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n379), .B(new_n386), .C1(new_n191), .C2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(G224), .A3(new_n200), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n394), .A2(new_n191), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n200), .A2(G224), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n386), .A4(new_n379), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n359), .A2(new_n401), .A3(new_n361), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n364), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n364), .A2(new_n400), .A3(KEYINPUT89), .A4(new_n402), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT7), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n395), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n360), .B(KEYINPUT8), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n356), .A2(new_n325), .ZN(new_n411));
  INV_X1    g225(.A(new_n337), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n396), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n363), .B1(new_n399), .B2(new_n408), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n188), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n312), .B1(new_n407), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n312), .ZN(new_n419));
  AOI211_X1 g233(.A(new_n419), .B(new_n416), .C1(new_n405), .C2(new_n406), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n187), .B(new_n311), .C1(new_n418), .C2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G221), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n289), .B2(new_n188), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G140), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n200), .A2(G227), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n355), .A2(new_n335), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n317), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n385), .A2(KEYINPUT10), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n356), .A2(KEYINPUT84), .A3(KEYINPUT10), .A4(new_n385), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n390), .A2(new_n391), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n376), .A2(new_n393), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n436), .A2(new_n437), .A3(new_n344), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n439), .B(KEYINPUT1), .C1(new_n265), .C2(G146), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G128), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n375), .B2(KEYINPUT1), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n369), .B1(new_n225), .B2(G143), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n380), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n430), .A2(new_n317), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT10), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n438), .A2(new_n343), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n435), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT11), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n270), .B2(G137), .ZN(new_n451));
  INV_X1    g265(.A(G137), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT11), .A3(G134), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n270), .A2(G137), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G131), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n451), .A2(new_n453), .A3(new_n211), .A4(new_n454), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n449), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n458), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n435), .A2(new_n448), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n428), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT12), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n431), .A2(new_n377), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n463), .B(new_n460), .C1(new_n464), .C2(new_n446), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n446), .B1(new_n385), .B2(new_n356), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT12), .B1(new_n466), .B2(new_n458), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n461), .A2(new_n428), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n469), .B2(KEYINPUT86), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n461), .A2(new_n471), .A3(new_n428), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n462), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(G469), .A3(new_n254), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n461), .B1(new_n465), .B2(new_n467), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n427), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n461), .A2(new_n477), .A3(new_n428), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n459), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n461), .B2(new_n428), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n476), .B(G469), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(G469), .A2(G902), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n424), .B1(new_n474), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n421), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT78), .ZN(new_n486));
  INV_X1    g300(.A(G234), .ZN(new_n487));
  OAI21_X1  g301(.A(G217), .B1(new_n254), .B2(new_n487), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n488), .B(KEYINPUT73), .Z(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n188), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT77), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT22), .B(G137), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n422), .A2(new_n487), .A3(G953), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT74), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n495), .B1(new_n348), .B2(G128), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n267), .A2(KEYINPUT74), .A3(G119), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n348), .A2(G128), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT24), .B(G110), .Z(new_n500));
  NAND3_X1  g314(.A1(new_n267), .A2(KEYINPUT23), .A3(G119), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n348), .A2(G128), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n498), .B(new_n501), .C1(new_n502), .C2(KEYINPUT23), .ZN(new_n503));
  OAI22_X1  g317(.A1(new_n499), .A2(new_n500), .B1(new_n503), .B2(G110), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n195), .A3(new_n226), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n499), .A2(new_n500), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(G110), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n506), .B(new_n507), .C1(new_n196), .C2(new_n197), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n494), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n505), .A2(new_n508), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT75), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n505), .A2(new_n508), .A3(KEYINPUT75), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n509), .B1(new_n514), .B2(new_n494), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n491), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n505), .A2(new_n508), .A3(KEYINPUT75), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT75), .B1(new_n505), .B2(new_n508), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n494), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n509), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n254), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT76), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(KEYINPUT25), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n489), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI22_X1  g338(.A1(new_n515), .A2(new_n254), .B1(new_n522), .B2(KEYINPUT25), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n486), .B(new_n516), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  INV_X1    g341(.A(new_n516), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT78), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT72), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT65), .B1(new_n444), .B2(new_n387), .ZN(new_n533));
  INV_X1    g347(.A(new_n391), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n458), .B(new_n437), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n351), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n270), .A2(G137), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n452), .A2(G134), .ZN(new_n538));
  OAI21_X1  g352(.A(G131), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n457), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n385), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n536), .B1(new_n535), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT28), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT29), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n535), .A2(new_n541), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n351), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n535), .A2(KEYINPUT70), .A3(new_n541), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT28), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n199), .A2(new_n200), .A3(G210), .ZN(new_n551));
  XOR2_X1   g365(.A(new_n551), .B(KEYINPUT27), .Z(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT26), .B(G101), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n545), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n532), .B1(new_n555), .B2(new_n254), .ZN(new_n556));
  INV_X1    g370(.A(new_n554), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n548), .A2(new_n549), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(KEYINPUT28), .ZN(new_n559));
  OAI211_X1 g373(.A(KEYINPUT72), .B(new_n302), .C1(new_n559), .C2(new_n545), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n457), .A2(new_n539), .A3(KEYINPUT66), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT66), .B1(new_n457), .B2(new_n539), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT67), .B1(new_n563), .B2(new_n377), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT67), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n385), .B(new_n565), .C1(new_n562), .C2(new_n561), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n566), .A3(new_n535), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n351), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT69), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT69), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n570), .A3(new_n351), .ZN(new_n571));
  INV_X1    g385(.A(new_n542), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n559), .B1(new_n573), .B2(KEYINPUT28), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT29), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n535), .A2(KEYINPUT30), .A3(new_n541), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT30), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n567), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n542), .B1(new_n579), .B2(new_n351), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n575), .B1(new_n580), .B2(new_n557), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n556), .B(new_n560), .C1(new_n574), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n567), .A2(new_n578), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(new_n351), .A3(new_n576), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n572), .A3(new_n557), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT31), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT31), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n580), .A2(new_n587), .A3(new_n557), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n550), .B1(new_n573), .B2(KEYINPUT28), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n586), .B(new_n588), .C1(new_n589), .C2(new_n557), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT32), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n591), .A2(G472), .A3(G902), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n582), .A2(G472), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(G472), .A2(G902), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n586), .A2(new_n588), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n385), .B1(new_n562), .B2(new_n561), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n596), .A2(KEYINPUT67), .B1(new_n394), .B2(new_n458), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n536), .B1(new_n597), .B2(new_n566), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n572), .B1(new_n598), .B2(new_n570), .ZN(new_n599));
  INV_X1    g413(.A(new_n571), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT28), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n550), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n557), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n594), .B1(new_n595), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n591), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n531), .B1(new_n593), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n485), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  OAI211_X1 g422(.A(new_n530), .B(new_n424), .C1(new_n474), .C2(new_n483), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(G472), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n590), .B2(new_n302), .ZN(new_n612));
  INV_X1    g426(.A(new_n604), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n407), .A2(new_n417), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n419), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n407), .A2(new_n312), .A3(new_n417), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n254), .A2(new_n295), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n291), .A2(new_n293), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(KEYINPUT33), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n291), .B2(new_n293), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n302), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT97), .B(G478), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT98), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n294), .A2(new_n630), .A3(new_n627), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n625), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n253), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n310), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n619), .A2(new_n187), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n615), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT99), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  XNOR2_X1  g453(.A(new_n309), .B(KEYINPUT100), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n187), .B(new_n640), .C1(new_n418), .C2(new_n420), .ZN(new_n641));
  INV_X1    g455(.A(new_n253), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n301), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n615), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT101), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT35), .B(G107), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NOR2_X1   g463(.A1(new_n494), .A2(KEYINPUT36), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n514), .B(new_n650), .Z(new_n651));
  INV_X1    g465(.A(new_n491), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n527), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n612), .A2(new_n613), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n485), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AOI21_X1  g473(.A(new_n655), .B1(new_n593), .B2(new_n605), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n481), .A2(new_n482), .ZN(new_n661));
  INV_X1    g475(.A(G469), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n461), .A2(new_n471), .A3(new_n428), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n471), .B1(new_n461), .B2(new_n428), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n663), .A2(new_n664), .A3(new_n468), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n662), .B(new_n302), .C1(new_n665), .C2(new_n462), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n423), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n303), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n308), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT102), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n253), .A2(new_n300), .A3(new_n672), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n187), .B(new_n673), .C1(new_n418), .C2(new_n420), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n660), .A2(new_n667), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(new_n671), .B(KEYINPUT39), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n667), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT40), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n590), .A2(new_n592), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n580), .A2(new_n554), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n542), .A2(new_n543), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n188), .B1(new_n684), .B2(new_n557), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n605), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT103), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n418), .A2(new_n420), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT38), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n253), .A2(new_n187), .A3(new_n301), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n691), .A2(new_n654), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n680), .A2(new_n689), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  AND3_X1   g509(.A1(new_n253), .A2(new_n632), .A3(new_n671), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n619), .A2(KEYINPUT104), .A3(new_n187), .A4(new_n696), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n187), .B(new_n696), .C1(new_n418), .C2(new_n420), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n697), .A2(new_n660), .A3(new_n700), .A4(new_n667), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  OAI21_X1  g516(.A(G469), .B1(new_n473), .B2(new_n254), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n424), .A3(new_n666), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT105), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n703), .A2(new_n666), .A3(new_n706), .A4(new_n424), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n635), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n606), .A3(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT41), .B(G113), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT106), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n710), .B(new_n712), .ZN(G15));
  NAND3_X1  g527(.A1(new_n708), .A2(new_n606), .A3(new_n644), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  INV_X1    g529(.A(new_n421), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n660), .A2(new_n716), .A3(new_n707), .A4(new_n705), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  INV_X1    g532(.A(new_n692), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n719), .B(new_n640), .C1(new_n418), .C2(new_n420), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n527), .A2(new_n528), .ZN(new_n722));
  INV_X1    g536(.A(new_n544), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n554), .B1(new_n723), .B2(new_n550), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n586), .A2(new_n588), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n725), .A2(new_n594), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n612), .A2(new_n722), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n721), .A2(new_n727), .A3(new_n707), .A4(new_n705), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NAND3_X1  g543(.A1(new_n253), .A2(new_n632), .A3(new_n671), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n612), .A2(new_n726), .A3(new_n655), .A4(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n187), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n690), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n731), .A2(new_n733), .A3(new_n707), .A4(new_n705), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  NAND2_X1  g549(.A1(new_n582), .A2(G472), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n605), .A2(new_n736), .A3(new_n681), .ZN(new_n737));
  INV_X1    g551(.A(new_n722), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n667), .A2(new_n690), .A3(new_n187), .A4(new_n696), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT42), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n617), .A2(new_n187), .A3(new_n618), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n484), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n730), .A2(KEYINPUT42), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n606), .A3(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NOR3_X1   g561(.A1(new_n418), .A2(new_n420), .A3(new_n732), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n737), .A2(new_n530), .A3(new_n748), .A4(new_n667), .ZN(new_n749));
  INV_X1    g563(.A(new_n673), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT107), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n743), .A2(new_n606), .A3(new_n752), .A4(new_n673), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  OAI21_X1  g569(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n662), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n757), .B2(new_n756), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n759), .A2(new_n482), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n666), .B1(new_n760), .B2(KEYINPUT46), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(KEYINPUT46), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n760), .A2(KEYINPUT108), .A3(KEYINPUT46), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n423), .ZN(new_n767));
  INV_X1    g581(.A(new_n632), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT109), .B1(new_n768), .B2(new_n253), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n773), .B(new_n654), .C1(new_n613), .C2(new_n612), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n742), .B1(new_n774), .B2(new_n775), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n678), .A2(new_n767), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n452), .ZN(G39));
  INV_X1    g593(.A(new_n737), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n531), .A3(new_n696), .A4(new_n748), .ZN(new_n781));
  INV_X1    g595(.A(new_n765), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT108), .B1(new_n760), .B2(KEYINPUT46), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(KEYINPUT47), .B(new_n424), .C1(new_n784), .C2(new_n761), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n766), .B2(new_n423), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n781), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n189), .ZN(G42));
  AOI21_X1  g603(.A(new_n722), .B1(new_n593), .B2(new_n605), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n708), .A2(new_n748), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT116), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n708), .A2(new_n794), .A3(new_n748), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n773), .A2(new_n307), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n791), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g613(.A(KEYINPUT117), .B(new_n797), .C1(new_n793), .C2(new_n795), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n790), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT48), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT48), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n803), .B(new_n790), .C1(new_n799), .C2(new_n800), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n773), .A2(new_n307), .A3(new_n727), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n806), .A2(new_n733), .A3(new_n708), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n688), .A2(new_n530), .A3(new_n307), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n795), .B2(new_n793), .ZN(new_n809));
  INV_X1    g623(.A(new_n633), .ZN(new_n810));
  AOI211_X1 g624(.A(new_n306), .B(new_n807), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n737), .A2(new_n705), .A3(new_n530), .A4(new_n707), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n635), .B2(new_n645), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n717), .A2(new_n728), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n485), .B1(new_n606), .B2(new_n656), .ZN(new_n817));
  INV_X1    g631(.A(new_n641), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n300), .B(KEYINPUT110), .Z(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n642), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n633), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n610), .A2(new_n818), .A3(new_n614), .A4(new_n821), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n741), .A2(new_n817), .A3(new_n745), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n737), .A2(new_n667), .A3(new_n654), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n819), .A2(new_n253), .A3(new_n672), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n748), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n751), .B2(new_n753), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT111), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n612), .A2(new_n655), .A3(new_n726), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n829), .B1(new_n831), .B2(new_n740), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n743), .A2(KEYINPUT111), .A3(new_n696), .A4(new_n830), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n816), .A2(new_n823), .A3(new_n828), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n690), .A2(new_n692), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n654), .A2(new_n672), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT112), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n836), .A2(new_n838), .A3(new_n687), .A4(new_n667), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n701), .A2(new_n734), .A3(new_n676), .A4(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT52), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n734), .B2(new_n676), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n835), .B(new_n841), .C1(new_n842), .C2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n817), .A2(new_n822), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n717), .A2(new_n728), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n708), .B(new_n606), .C1(new_n709), .C2(new_n644), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n746), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n827), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n754), .A2(new_n834), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n840), .B(new_n843), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT53), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT54), .B1(new_n846), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n842), .B1(new_n841), .B2(new_n835), .ZN(new_n857));
  INV_X1    g671(.A(new_n852), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n848), .A2(new_n859), .A3(new_n849), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT113), .B1(new_n814), .B2(new_n815), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n741), .A2(new_n817), .A3(new_n745), .A4(new_n822), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n863), .A2(new_n844), .A3(new_n842), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n854), .A2(new_n858), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n857), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n691), .A2(new_n732), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n806), .A2(new_n868), .A3(new_n708), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT50), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n806), .A2(new_n868), .A3(KEYINPUT50), .A4(new_n708), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n253), .A2(new_n632), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n871), .A2(new_n872), .B1(new_n809), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n703), .A2(new_n423), .A3(new_n666), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n785), .A2(new_n787), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n806), .A2(new_n748), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n830), .B1(new_n799), .B2(new_n800), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n874), .A2(new_n878), .A3(new_n879), .A4(KEYINPUT51), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n812), .A2(new_n856), .A3(new_n867), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n785), .A2(new_n787), .A3(KEYINPUT114), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n875), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT114), .B1(new_n785), .B2(new_n787), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n877), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(KEYINPUT115), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n874), .A2(new_n879), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n885), .B2(KEYINPUT115), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT51), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI22_X1  g703(.A1(new_n881), .A2(new_n889), .B1(G952), .B2(G953), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n703), .A2(new_n666), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n891), .A2(KEYINPUT49), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(KEYINPUT49), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n722), .A2(new_n423), .A3(new_n732), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n642), .A3(new_n632), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n688), .A2(new_n691), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n890), .A2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n200), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n302), .B1(new_n857), .B2(new_n865), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n419), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n364), .A2(new_n402), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(new_n400), .Z(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n900), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT56), .B1(new_n902), .B2(KEYINPUT118), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(KEYINPUT118), .B2(new_n902), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(new_n906), .ZN(G51));
  AOI211_X1 g725(.A(new_n302), .B(new_n759), .C1(new_n857), .C2(new_n865), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n482), .B(KEYINPUT57), .Z(new_n913));
  AND3_X1   g727(.A1(new_n857), .A2(new_n865), .A3(new_n866), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n866), .B1(new_n857), .B2(new_n865), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n473), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT119), .B1(new_n918), .B2(new_n899), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  INV_X1    g734(.A(new_n862), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n734), .A2(new_n676), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n842), .B1(new_n922), .B2(KEYINPUT52), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n823), .A3(new_n828), .A4(new_n834), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n921), .A2(new_n841), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT54), .B1(new_n925), .B2(new_n855), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n867), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n473), .B1(new_n927), .B2(new_n913), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n920), .B(new_n900), .C1(new_n928), .C2(new_n912), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n919), .A2(new_n929), .ZN(G54));
  NAND3_X1  g744(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  INV_X1    g745(.A(new_n248), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n931), .A2(KEYINPUT120), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n900), .B1(new_n931), .B2(new_n932), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT120), .B1(new_n931), .B2(new_n932), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G60));
  NOR2_X1   g750(.A1(new_n622), .A2(new_n624), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT121), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n856), .A2(new_n867), .ZN(new_n939));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT59), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n927), .A2(new_n938), .A3(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n899), .A3(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT60), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n857), .B2(new_n865), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n947), .A2(new_n651), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n519), .A2(new_n520), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n900), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(KEYINPUT122), .A3(new_n952), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n952), .A2(KEYINPUT122), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(KEYINPUT122), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n954), .B(new_n955), .C1(new_n948), .C2(new_n950), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n953), .A2(new_n956), .ZN(G66));
  INV_X1    g771(.A(G224), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n304), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n816), .A2(new_n847), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n961), .B2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n904), .B1(G898), .B2(new_n200), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G69));
  AOI21_X1  g778(.A(new_n200), .B1(G227), .B2(G900), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n778), .A2(new_n788), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n767), .A2(new_n678), .A3(new_n836), .A4(new_n790), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n701), .A2(new_n676), .A3(new_n734), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n969), .A2(new_n746), .A3(new_n754), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(G953), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n579), .B(KEYINPUT123), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(new_n245), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(G900), .B2(G953), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n694), .A2(new_n969), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT62), .Z(new_n978));
  XNOR2_X1  g792(.A(new_n821), .B(KEYINPUT125), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n979), .A2(new_n606), .A3(new_n679), .A4(new_n748), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n967), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n981), .A2(new_n200), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n974), .B(KEYINPUT124), .ZN(new_n983));
  OAI221_X1 g797(.A(new_n966), .B1(new_n972), .B2(new_n976), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n972), .A2(new_n976), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n983), .B1(new_n981), .B2(new_n200), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n965), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(G72));
  XNOR2_X1  g802(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n611), .A2(new_n188), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n989), .B(new_n990), .Z(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT127), .Z(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n971), .B2(new_n960), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n580), .A2(new_n554), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n899), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n992), .B1(new_n981), .B2(new_n960), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n682), .ZN(new_n997));
  INV_X1    g811(.A(new_n991), .ZN(new_n998));
  INV_X1    g812(.A(new_n585), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n580), .A2(new_n557), .ZN(new_n1000));
  OAI221_X1 g814(.A(new_n998), .B1(new_n999), .B2(new_n1000), .C1(new_n846), .C2(new_n855), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n995), .A2(new_n997), .A3(new_n1001), .ZN(G57));
endmodule


