

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U321 ( .A(n412), .B(n411), .ZN(n413) );
  INV_X1 U322 ( .A(n421), .ZN(n422) );
  XNOR2_X1 U323 ( .A(n423), .B(n422), .ZN(n424) );
  NOR2_X1 U324 ( .A1(n461), .A2(n449), .ZN(n289) );
  NOR2_X1 U325 ( .A1(n580), .A2(n550), .ZN(n290) );
  XNOR2_X1 U326 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n407) );
  INV_X1 U327 ( .A(KEYINPUT100), .ZN(n467) );
  XNOR2_X1 U328 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U329 ( .A(n408), .B(n407), .ZN(n565) );
  XNOR2_X1 U330 ( .A(n419), .B(n295), .ZN(n296) );
  XNOR2_X1 U331 ( .A(n375), .B(n296), .ZN(n297) );
  AND2_X1 U332 ( .A1(n480), .A2(n290), .ZN(n473) );
  XNOR2_X1 U333 ( .A(n425), .B(n424), .ZN(n429) );
  XNOR2_X1 U334 ( .A(n308), .B(n307), .ZN(n536) );
  INV_X1 U335 ( .A(G43GAT), .ZN(n475) );
  XOR2_X1 U336 ( .A(n461), .B(KEYINPUT28), .Z(n529) );
  XNOR2_X1 U337 ( .A(n453), .B(G190GAT), .ZN(n454) );
  XNOR2_X1 U338 ( .A(n475), .B(KEYINPUT40), .ZN(n476) );
  XNOR2_X1 U339 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n477), .B(n476), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(G99GAT), .B(G85GAT), .Z(n351) );
  XOR2_X1 U342 ( .A(KEYINPUT75), .B(n351), .Z(n292) );
  XOR2_X1 U343 ( .A(G36GAT), .B(G190GAT), .Z(n392) );
  XNOR2_X1 U344 ( .A(G92GAT), .B(n392), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n292), .B(n291), .ZN(n298) );
  XOR2_X1 U346 ( .A(G29GAT), .B(G43GAT), .Z(n294) );
  XNOR2_X1 U347 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n375) );
  XOR2_X1 U349 ( .A(G50GAT), .B(G162GAT), .Z(n419) );
  AND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U351 ( .A(n298), .B(n297), .Z(n300) );
  XNOR2_X1 U352 ( .A(G218GAT), .B(G106GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n308) );
  XOR2_X1 U354 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n302) );
  XNOR2_X1 U355 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U357 ( .A(KEYINPUT74), .B(KEYINPUT64), .Z(n304) );
  XNOR2_X1 U358 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U361 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n310) );
  XNOR2_X1 U362 ( .A(G190GAT), .B(G99GAT), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U364 ( .A(n311), .B(G71GAT), .Z(n313) );
  XOR2_X1 U365 ( .A(G15GAT), .B(G127GAT), .Z(n334) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(n334), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n319) );
  XOR2_X1 U368 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n315) );
  XNOR2_X1 U369 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n395) );
  XOR2_X1 U371 ( .A(G113GAT), .B(n395), .Z(n317) );
  NAND2_X1 U372 ( .A1(G227GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U374 ( .A(n319), .B(n318), .Z(n327) );
  XOR2_X1 U375 ( .A(KEYINPUT82), .B(G134GAT), .Z(n321) );
  XNOR2_X1 U376 ( .A(KEYINPUT81), .B(G120GAT), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U378 ( .A(KEYINPUT0), .B(n322), .Z(n437) );
  XOR2_X1 U379 ( .A(G176GAT), .B(G183GAT), .Z(n324) );
  XNOR2_X1 U380 ( .A(KEYINPUT84), .B(KEYINPUT20), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n437), .B(n325), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n527) );
  XOR2_X1 U384 ( .A(KEYINPUT45), .B(KEYINPUT115), .Z(n349) );
  XNOR2_X1 U385 ( .A(KEYINPUT107), .B(KEYINPUT36), .ZN(n328) );
  XOR2_X1 U386 ( .A(n328), .B(n536), .Z(n580) );
  XOR2_X1 U387 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n330) );
  XNOR2_X1 U388 ( .A(G1GAT), .B(G64GAT), .ZN(n329) );
  XNOR2_X1 U389 ( .A(n330), .B(n329), .ZN(n347) );
  XOR2_X1 U390 ( .A(G78GAT), .B(G211GAT), .Z(n332) );
  XNOR2_X1 U391 ( .A(G22GAT), .B(G155GAT), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U393 ( .A(n334), .B(n333), .Z(n336) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U396 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n338) );
  XNOR2_X1 U397 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U399 ( .A(n340), .B(n339), .Z(n345) );
  XNOR2_X1 U400 ( .A(G8GAT), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n341), .B(KEYINPUT76), .ZN(n391) );
  XOR2_X1 U402 ( .A(G57GAT), .B(KEYINPUT67), .Z(n343) );
  XNOR2_X1 U403 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n391), .B(n350), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U407 ( .A(n347), .B(n346), .Z(n550) );
  INV_X1 U408 ( .A(n550), .ZN(n578) );
  NOR2_X1 U409 ( .A1(n580), .A2(n578), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n367) );
  XOR2_X1 U411 ( .A(KEYINPUT31), .B(n350), .Z(n353) );
  XNOR2_X1 U412 ( .A(G120GAT), .B(n351), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n358) );
  XNOR2_X1 U414 ( .A(G106GAT), .B(G78GAT), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n354), .B(G148GAT), .ZN(n421) );
  XOR2_X1 U416 ( .A(n421), .B(KEYINPUT69), .Z(n356) );
  NAND2_X1 U417 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U419 ( .A(n358), .B(n357), .Z(n366) );
  XOR2_X1 U420 ( .A(G92GAT), .B(G64GAT), .Z(n360) );
  XNOR2_X1 U421 ( .A(G176GAT), .B(KEYINPUT70), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U423 ( .A(G204GAT), .B(n361), .Z(n403) );
  XOR2_X1 U424 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n363) );
  XNOR2_X1 U425 ( .A(KEYINPUT71), .B(KEYINPUT68), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n403), .B(n364), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n575) );
  AND2_X1 U429 ( .A1(n367), .A2(n575), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n368), .B(KEYINPUT116), .ZN(n383) );
  XOR2_X1 U431 ( .A(G8GAT), .B(G197GAT), .Z(n370) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(G15GAT), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U434 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n372) );
  XNOR2_X1 U435 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n382) );
  XOR2_X1 U438 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XOR2_X1 U439 ( .A(n375), .B(n420), .Z(n377) );
  NAND2_X1 U440 ( .A1(G229GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U442 ( .A(G113GAT), .B(G1GAT), .Z(n433) );
  XOR2_X1 U443 ( .A(n378), .B(n433), .Z(n380) );
  XNOR2_X1 U444 ( .A(G50GAT), .B(G36GAT), .ZN(n379) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U446 ( .A(n382), .B(n381), .Z(n541) );
  INV_X1 U447 ( .A(n541), .ZN(n570) );
  NAND2_X1 U448 ( .A1(n383), .A2(n570), .ZN(n389) );
  INV_X1 U449 ( .A(n536), .ZN(n553) );
  XNOR2_X1 U450 ( .A(n575), .B(KEYINPUT41), .ZN(n543) );
  NAND2_X1 U451 ( .A1(n541), .A2(n543), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n384), .B(KEYINPUT46), .ZN(n385) );
  NAND2_X1 U453 ( .A1(n385), .A2(n578), .ZN(n386) );
  NOR2_X1 U454 ( .A1(n553), .A2(n386), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n387), .B(KEYINPUT47), .ZN(n388) );
  NAND2_X1 U456 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n390), .B(KEYINPUT48), .ZN(n526) );
  XOR2_X1 U458 ( .A(n391), .B(KEYINPUT95), .Z(n394) );
  XNOR2_X1 U459 ( .A(n392), .B(KEYINPUT96), .ZN(n393) );
  XNOR2_X1 U460 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U461 ( .A(n395), .B(KEYINPUT94), .Z(n397) );
  NAND2_X1 U462 ( .A1(G226GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U464 ( .A(n399), .B(n398), .Z(n405) );
  XOR2_X1 U465 ( .A(KEYINPUT88), .B(G218GAT), .Z(n401) );
  XNOR2_X1 U466 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U468 ( .A(G197GAT), .B(n402), .Z(n416) );
  XNOR2_X1 U469 ( .A(n416), .B(n403), .ZN(n404) );
  XOR2_X1 U470 ( .A(n405), .B(n404), .Z(n517) );
  INV_X1 U471 ( .A(n517), .ZN(n406) );
  NAND2_X1 U472 ( .A1(n526), .A2(n406), .ZN(n408) );
  XOR2_X1 U473 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n410) );
  XNOR2_X1 U474 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n414) );
  NAND2_X1 U476 ( .A1(G228GAT), .A2(G233GAT), .ZN(n412) );
  INV_X1 U477 ( .A(KEYINPUT91), .ZN(n411) );
  XOR2_X1 U478 ( .A(n415), .B(G204GAT), .Z(n418) );
  XNOR2_X1 U479 ( .A(n416), .B(KEYINPUT23), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n423) );
  XOR2_X1 U482 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n427) );
  XNOR2_X1 U483 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U485 ( .A(KEYINPUT2), .B(n428), .Z(n444) );
  XOR2_X1 U486 ( .A(n429), .B(n444), .Z(n461) );
  XOR2_X1 U487 ( .A(G85GAT), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U488 ( .A(G141GAT), .B(G162GAT), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U490 ( .A(n432), .B(G127GAT), .Z(n435) );
  XNOR2_X1 U491 ( .A(n433), .B(G29GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n448) );
  XOR2_X1 U494 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n439) );
  XNOR2_X1 U495 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U497 ( .A(KEYINPUT93), .B(n440), .Z(n442) );
  NAND2_X1 U498 ( .A1(G225GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U500 ( .A(n443), .B(KEYINPUT5), .Z(n446) );
  XNOR2_X1 U501 ( .A(n444), .B(G57GAT), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n566) );
  INV_X1 U504 ( .A(n566), .ZN(n449) );
  AND2_X1 U505 ( .A1(n565), .A2(n289), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NOR2_X1 U507 ( .A1(n527), .A2(n451), .ZN(n452) );
  XOR2_X1 U508 ( .A(KEYINPUT122), .B(n452), .Z(n561) );
  NOR2_X1 U509 ( .A1(n536), .A2(n561), .ZN(n455) );
  INV_X1 U510 ( .A(KEYINPUT58), .ZN(n453) );
  NAND2_X1 U511 ( .A1(n575), .A2(n541), .ZN(n482) );
  XNOR2_X1 U512 ( .A(n517), .B(KEYINPUT27), .ZN(n464) );
  NOR2_X1 U513 ( .A1(n464), .A2(n566), .ZN(n456) );
  XOR2_X1 U514 ( .A(n456), .B(KEYINPUT97), .Z(n525) );
  AND2_X1 U515 ( .A1(n525), .A2(n529), .ZN(n457) );
  NAND2_X1 U516 ( .A1(n527), .A2(n457), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n458), .B(KEYINPUT98), .ZN(n471) );
  NOR2_X1 U518 ( .A1(n527), .A2(n517), .ZN(n459) );
  NOR2_X1 U519 ( .A1(n461), .A2(n459), .ZN(n460) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n460), .Z(n466) );
  XOR2_X1 U521 ( .A(KEYINPUT99), .B(KEYINPUT26), .Z(n463) );
  NAND2_X1 U522 ( .A1(n461), .A2(n527), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n463), .B(n462), .ZN(n568) );
  NOR2_X1 U524 ( .A1(n568), .A2(n464), .ZN(n465) );
  NOR2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n469), .A2(n566), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n480) );
  XNOR2_X1 U529 ( .A(KEYINPUT108), .B(KEYINPUT37), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n473), .B(n472), .ZN(n514) );
  NOR2_X1 U531 ( .A1(n482), .A2(n514), .ZN(n474) );
  XOR2_X1 U532 ( .A(n474), .B(KEYINPUT38), .Z(n500) );
  NOR2_X1 U533 ( .A1(n527), .A2(n500), .ZN(n477) );
  XOR2_X1 U534 ( .A(KEYINPUT80), .B(KEYINPUT16), .Z(n479) );
  NAND2_X1 U535 ( .A1(n550), .A2(n536), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(n481) );
  NAND2_X1 U537 ( .A1(n481), .A2(n480), .ZN(n504) );
  NOR2_X1 U538 ( .A1(n504), .A2(n482), .ZN(n483) );
  XNOR2_X1 U539 ( .A(n483), .B(KEYINPUT101), .ZN(n492) );
  NOR2_X1 U540 ( .A1(n566), .A2(n492), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT34), .B(n484), .Z(n485) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U543 ( .A1(n517), .A2(n492), .ZN(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  NOR2_X1 U547 ( .A1(n527), .A2(n492), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n491), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n529), .A2(n492), .ZN(n494) );
  XNOR2_X1 U552 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1327GAT) );
  NOR2_X1 U554 ( .A1(n500), .A2(n566), .ZN(n498) );
  XOR2_X1 U555 ( .A(KEYINPUT106), .B(KEYINPUT109), .Z(n496) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n500), .A2(n517), .ZN(n499) );
  XOR2_X1 U560 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  INV_X1 U561 ( .A(G50GAT), .ZN(n502) );
  NOR2_X1 U562 ( .A1(n529), .A2(n500), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U564 ( .A(KEYINPUT110), .B(n503), .ZN(G1331GAT) );
  NAND2_X1 U565 ( .A1(n570), .A2(n543), .ZN(n513) );
  OR2_X1 U566 ( .A1(n513), .A2(n504), .ZN(n510) );
  NOR2_X1 U567 ( .A1(n566), .A2(n510), .ZN(n506) );
  XNOR2_X1 U568 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n507), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n510), .ZN(n508) );
  XOR2_X1 U572 ( .A(G64GAT), .B(n508), .Z(G1333GAT) );
  NOR2_X1 U573 ( .A1(n527), .A2(n510), .ZN(n509) );
  XOR2_X1 U574 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U575 ( .A1(n529), .A2(n510), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U578 ( .A1(n514), .A2(n513), .ZN(n515) );
  XOR2_X1 U579 ( .A(KEYINPUT112), .B(n515), .Z(n521) );
  NOR2_X1 U580 ( .A1(n566), .A2(n521), .ZN(n516) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n516), .Z(G1336GAT) );
  NOR2_X1 U582 ( .A1(n521), .A2(n517), .ZN(n518) );
  XOR2_X1 U583 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n520) );
  NOR2_X1 U585 ( .A1(n527), .A2(n521), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  XNOR2_X1 U587 ( .A(KEYINPUT114), .B(KEYINPUT44), .ZN(n523) );
  NOR2_X1 U588 ( .A1(n529), .A2(n521), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U590 ( .A(G106GAT), .B(n524), .Z(G1339GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n539) );
  NOR2_X1 U592 ( .A1(n527), .A2(n539), .ZN(n528) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n535) );
  NOR2_X1 U594 ( .A1(n570), .A2(n535), .ZN(n530) );
  XOR2_X1 U595 ( .A(G113GAT), .B(n530), .Z(G1340GAT) );
  INV_X1 U596 ( .A(n543), .ZN(n557) );
  NOR2_X1 U597 ( .A1(n557), .A2(n535), .ZN(n532) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U600 ( .A1(n578), .A2(n535), .ZN(n533) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(n533), .Z(n534) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  NOR2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n568), .A2(n539), .ZN(n540) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(n540), .Z(n552) );
  NAND2_X1 U608 ( .A1(n541), .A2(n552), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(G141GAT), .ZN(G1344GAT) );
  NAND2_X1 U610 ( .A1(n543), .A2(n552), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n545) );
  XNOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U621 ( .A1(n561), .A2(n570), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(KEYINPUT123), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(n556), .ZN(G1348GAT) );
  XNOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n559) );
  NOR2_X1 U625 ( .A1(n557), .A2(n561), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G176GAT), .ZN(G1349GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n578), .ZN(n563) );
  XNOR2_X1 U629 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(n564), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n566), .ZN(n567) );
  NOR2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT126), .B(n569), .Z(n581) );
  NOR2_X1 U635 ( .A1(n581), .A2(n570), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n577) );
  NOR2_X1 U641 ( .A1(n575), .A2(n581), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n581), .A2(n578), .ZN(n579) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

