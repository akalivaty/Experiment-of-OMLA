//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  XOR2_X1   g0004(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT65), .ZN(new_n206));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n206), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  NOR2_X1   g0015(.A1(G58), .A2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT66), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n213), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT67), .B(G68), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n210), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n220), .B1(KEYINPUT1), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT16), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(KEYINPUT7), .B1(new_n251), .B2(new_n208), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT7), .ZN(new_n254));
  NOR4_X1   g0054(.A1(new_n249), .A2(new_n250), .A3(new_n254), .A4(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n222), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  OR2_X1    g0058(.A1(KEYINPUT67), .A2(G68), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT67), .A2(G68), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(G20), .B1(new_n261), .B2(new_n216), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G159), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n248), .B1(new_n257), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n214), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT75), .B1(new_n262), .B2(new_n267), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT67), .A2(G68), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT67), .A2(G68), .ZN(new_n276));
  OAI21_X1  g0076(.A(G58), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n208), .B1(new_n277), .B2(new_n217), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT75), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n278), .A2(new_n279), .A3(new_n266), .ZN(new_n280));
  OR2_X1    g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(KEYINPUT74), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT74), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(new_n249), .B2(new_n250), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n285), .A3(new_n208), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n255), .B1(new_n286), .B2(new_n254), .ZN(new_n287));
  INV_X1    g0087(.A(G68), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n274), .A2(new_n280), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n289), .A2(KEYINPUT76), .A3(new_n248), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT76), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n286), .A2(new_n254), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n256), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n279), .B1(new_n278), .B2(new_n266), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n216), .B1(new_n221), .B2(G58), .ZN(new_n295));
  OAI211_X1 g0095(.A(KEYINPUT75), .B(new_n267), .C1(new_n295), .C2(new_n208), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n293), .A2(G68), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n291), .B1(new_n297), .B2(KEYINPUT16), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n273), .B1(new_n290), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT68), .B1(new_n258), .B2(KEYINPUT8), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(KEYINPUT68), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n300), .C1(new_n301), .C2(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n271), .B1(new_n207), .B2(G20), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n306), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G41), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(G1), .A3(G13), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT3), .B(G33), .ZN(new_n314));
  INV_X1    g0114(.A(G223), .ZN(new_n315));
  INV_X1    g0115(.A(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n314), .B(new_n317), .C1(G226), .C2(new_n316), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G87), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n313), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G41), .ZN(new_n322));
  INV_X1    g0122(.A(G45), .ZN(new_n323));
  AOI21_X1  g0123(.A(G1), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n324), .A2(new_n313), .A3(G274), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n324), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(G232), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(G190), .B2(new_n329), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n299), .A2(new_n311), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT17), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT71), .B(G179), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n321), .A2(new_n337), .A3(new_n328), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT77), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n327), .A2(G232), .ZN(new_n340));
  INV_X1    g0140(.A(new_n325), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(G169), .B1(new_n342), .B2(new_n320), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n338), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n339), .B1(new_n338), .B2(new_n343), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT76), .B1(new_n289), .B2(new_n248), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n297), .A2(new_n291), .A3(KEYINPUT16), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n272), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n346), .B1(new_n349), .B2(new_n310), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT18), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT18), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(new_n346), .C1(new_n349), .C2(new_n310), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n299), .A2(KEYINPUT17), .A3(new_n311), .A4(new_n332), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n335), .A2(new_n351), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n309), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT72), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT72), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n309), .A2(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n271), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(G68), .C1(G1), .C2(new_n208), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT12), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n309), .B2(G68), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(KEYINPUT12), .A3(new_n222), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n208), .A2(G33), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT70), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G77), .ZN(new_n370));
  INV_X1    g0170(.A(G50), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n370), .B1(new_n208), .B2(new_n221), .C1(new_n371), .C2(new_n264), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n372), .A2(KEYINPUT11), .A3(new_n271), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT11), .B1(new_n372), .B2(new_n271), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n366), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n314), .A2(G232), .A3(G1698), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n314), .A2(G226), .A3(new_n316), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G97), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n326), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n325), .B1(G238), .B2(new_n327), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT13), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT13), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n385), .A3(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT14), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n388), .A3(G169), .ZN(new_n389));
  INV_X1    g0189(.A(G179), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(new_n387), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n387), .B2(G169), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n376), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n387), .A2(G200), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n375), .B(new_n394), .C1(new_n395), .C2(new_n387), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n314), .A2(G232), .A3(new_n316), .ZN(new_n397));
  INV_X1    g0197(.A(G107), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n314), .A2(G1698), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n397), .B1(new_n398), .B2(new_n314), .C1(new_n399), .C2(new_n223), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n326), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n325), .B1(G244), .B2(new_n327), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G200), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n401), .A2(G190), .A3(new_n402), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n361), .B(G77), .C1(G1), .C2(new_n208), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G20), .A2(G77), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT15), .B(G87), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n407), .B1(new_n408), .B2(new_n367), .C1(new_n264), .C2(new_n301), .ZN(new_n409));
  INV_X1    g0209(.A(G77), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n409), .A2(new_n271), .B1(new_n360), .B2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n404), .A2(new_n405), .A3(new_n406), .A4(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G169), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n403), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n406), .A2(new_n411), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(new_n415), .C1(new_n337), .C2(new_n403), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n393), .A2(new_n396), .A3(new_n412), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n271), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n303), .A2(new_n305), .A3(new_n369), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n371), .A2(new_n258), .A3(new_n288), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(G20), .B1(G150), .B2(new_n263), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n307), .A2(G50), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G50), .B2(new_n309), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT9), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n314), .A2(G222), .A3(new_n316), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n428), .B1(new_n410), .B2(new_n314), .C1(new_n399), .C2(new_n315), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n326), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n325), .B1(G226), .B2(new_n327), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n330), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n430), .A2(new_n431), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n432), .B1(G190), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n427), .A2(KEYINPUT73), .A3(KEYINPUT10), .A4(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n425), .A2(new_n426), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n422), .A2(KEYINPUT9), .A3(new_n424), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n439));
  OR2_X1    g0239(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n433), .A2(new_n336), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n442), .B1(G169), .B2(new_n433), .C1(new_n422), .C2(new_n424), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n435), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n355), .A2(new_n417), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n323), .A2(G1), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(G264), .A3(new_n313), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT84), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n326), .B1(new_n447), .B2(new_n446), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT84), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(G264), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n446), .A2(G274), .A3(new_n313), .A4(new_n447), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n314), .A2(G257), .A3(G1698), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n314), .A2(G250), .A3(new_n316), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G294), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n456), .B1(new_n460), .B2(new_n326), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n330), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n395), .A3(new_n449), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n356), .A2(KEYINPUT25), .A3(new_n398), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT83), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT25), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n309), .B2(G107), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n469), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n207), .A2(G33), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n418), .A2(new_n472), .A3(new_n309), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n470), .A2(new_n471), .B1(G107), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n208), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT22), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n314), .A2(new_n478), .A3(new_n208), .A4(G87), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n398), .A2(KEYINPUT23), .A3(G20), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT23), .B1(new_n398), .B2(G20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G116), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n481), .A2(new_n482), .B1(G20), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT24), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n480), .A2(new_n488), .A3(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT82), .B1(new_n490), .B2(new_n271), .ZN(new_n491));
  AOI211_X1 g0291(.A(KEYINPUT24), .B(new_n484), .C1(new_n477), .C2(new_n479), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n488), .B1(new_n480), .B2(new_n485), .ZN(new_n493));
  OAI211_X1 g0293(.A(KEYINPUT82), .B(new_n271), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n465), .B(new_n475), .C1(new_n491), .C2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT85), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n461), .A2(new_n449), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G169), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n390), .B2(new_n462), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n475), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n271), .B1(new_n492), .B2(new_n493), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT82), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n505), .B2(new_n494), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n496), .B(new_n497), .C1(new_n501), .C2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n475), .B1(new_n491), .B2(new_n495), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n500), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n497), .B1(new_n510), .B2(new_n496), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n314), .A2(new_n208), .A3(G68), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT19), .ZN(new_n514));
  INV_X1    g0314(.A(G97), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n514), .B1(new_n367), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n518));
  INV_X1    g0318(.A(G87), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n208), .A2(new_n518), .B1(new_n202), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n271), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n360), .A2(new_n408), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n474), .A2(G87), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G250), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n323), .B2(G1), .ZN(new_n526));
  INV_X1    g0326(.A(G274), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n207), .A2(new_n527), .A3(G45), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n313), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(G238), .B(new_n316), .C1(new_n249), .C2(new_n250), .ZN(new_n531));
  OAI21_X1  g0331(.A(G244), .B1(new_n249), .B2(new_n250), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(new_n483), .C1(new_n532), .C2(new_n316), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n533), .B2(new_n326), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n534), .A2(new_n330), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(G190), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n524), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n521), .B(new_n522), .C1(new_n473), .C2(new_n408), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n533), .A2(new_n326), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n413), .B1(new_n539), .B2(new_n529), .ZN(new_n540));
  AOI211_X1 g0340(.A(new_n336), .B(new_n530), .C1(new_n533), .C2(new_n326), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(KEYINPUT4), .A2(G244), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n316), .B(new_n545), .C1(new_n249), .C2(new_n250), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G283), .ZN(new_n547));
  INV_X1    g0347(.A(G244), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n281), .B2(new_n282), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n546), .B(new_n547), .C1(new_n549), .C2(KEYINPUT4), .ZN(new_n550));
  OAI21_X1  g0350(.A(G250), .B1(new_n249), .B2(new_n250), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n316), .B1(new_n551), .B2(KEYINPUT4), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n326), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n448), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n326), .A2(new_n527), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n451), .A2(G257), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n553), .A2(new_n556), .A3(new_n336), .ZN(new_n557));
  AOI21_X1  g0357(.A(G169), .B1(new_n553), .B2(new_n556), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT78), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n264), .A2(new_n410), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g0362(.A(G97), .B(G107), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT6), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n515), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n563), .A2(new_n564), .B1(new_n398), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n560), .B(new_n562), .C1(new_n566), .C2(new_n208), .ZN(new_n567));
  AND2_X1   g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n564), .B1(new_n568), .B2(new_n202), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n398), .A2(KEYINPUT6), .A3(G97), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n208), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT78), .B1(new_n571), .B2(new_n561), .ZN(new_n572));
  OAI21_X1  g0372(.A(G107), .B1(new_n252), .B2(new_n255), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n567), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n271), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n309), .A2(G97), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n473), .B2(new_n515), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT79), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n559), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n553), .A2(new_n556), .A3(new_n336), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n448), .A2(G257), .A3(new_n313), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n455), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n525), .B1(new_n281), .B2(new_n282), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  OAI21_X1  g0387(.A(G1698), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n532), .A2(new_n587), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n588), .A2(new_n547), .A3(new_n546), .A4(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n585), .B1(new_n590), .B2(new_n326), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n583), .B1(new_n591), .B2(G169), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n578), .B1(new_n574), .B2(new_n271), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT79), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n553), .A2(new_n556), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G200), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n593), .B(new_n596), .C1(new_n395), .C2(new_n595), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n544), .A2(new_n582), .A3(new_n594), .A4(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n456), .B1(G270), .B2(new_n451), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n314), .A2(G264), .A3(G1698), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n314), .A2(G257), .A3(new_n316), .ZN(new_n601));
  INV_X1    g0401(.A(G303), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n600), .B(new_n601), .C1(new_n602), .C2(new_n314), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n326), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n357), .A2(new_n359), .ZN(new_n606));
  INV_X1    g0406(.A(G116), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n207), .B2(G33), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n418), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n547), .B(new_n208), .C1(G33), .C2(new_n515), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(G20), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n271), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT80), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(KEYINPUT20), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n357), .A2(new_n607), .A3(new_n359), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(KEYINPUT20), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n612), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n609), .A2(new_n616), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n605), .A2(KEYINPUT21), .A3(new_n620), .A4(G169), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n413), .B1(new_n599), .B2(new_n604), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT81), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT21), .A4(new_n620), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(new_n620), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n599), .A2(new_n604), .A3(G179), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n627), .A2(new_n628), .B1(new_n630), .B2(new_n620), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n620), .B1(new_n605), .B2(G200), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n395), .B2(new_n605), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n626), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n598), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n445), .A2(new_n512), .A3(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n393), .A2(new_n416), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n335), .A2(new_n637), .A3(new_n354), .A4(new_n396), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n351), .A2(new_n353), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n441), .B(new_n435), .C1(new_n638), .C2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(new_n443), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT86), .B1(new_n540), .B2(new_n541), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n539), .A2(new_n337), .A3(new_n529), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT86), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n644), .B(new_n645), .C1(new_n413), .C2(new_n534), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n538), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n592), .A2(new_n593), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n534), .A2(new_n330), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(KEYINPUT87), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT87), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n534), .A2(new_n652), .A3(new_n330), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n536), .B(new_n524), .C1(new_n651), .C2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n648), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n581), .B1(new_n559), .B2(new_n580), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT79), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n544), .B(KEYINPUT26), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n626), .B(new_n631), .C1(new_n506), .C2(new_n501), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n524), .A2(new_n536), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n535), .A2(new_n652), .ZN(new_n664));
  INV_X1    g0464(.A(new_n653), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n506), .B2(new_n465), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n582), .A2(new_n594), .A3(new_n597), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n662), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n661), .A2(new_n669), .A3(new_n648), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n445), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n642), .A2(new_n671), .ZN(G369));
  NAND3_X1  g0472(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n509), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n510), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n512), .A2(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n626), .A2(new_n631), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n620), .A2(new_n678), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT88), .Z(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(new_n633), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n682), .B2(new_n684), .ZN(new_n686));
  XOR2_X1   g0486(.A(KEYINPUT89), .B(G330), .Z(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n681), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n682), .A2(new_n678), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n512), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n510), .B2(new_n678), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT90), .Z(G399));
  INV_X1    g0495(.A(new_n211), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n218), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  INV_X1    g0502(.A(new_n678), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT29), .B1(new_n670), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n655), .A2(new_n656), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n544), .B1(new_n658), .B2(new_n659), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT92), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n656), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n543), .B1(new_n582), .B2(new_n594), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT92), .B1(new_n709), .B2(KEYINPUT26), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n705), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n648), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n496), .A2(new_n654), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n582), .A2(new_n594), .A3(new_n597), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n712), .B1(new_n715), .B2(new_n662), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n678), .B1(new_n711), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n704), .B1(KEYINPUT29), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n635), .B(new_n703), .C1(new_n508), .C2(new_n511), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n460), .A2(new_n326), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n591), .A2(new_n721), .A3(new_n454), .A4(new_n534), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n722), .B2(new_n629), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n454), .A2(new_n721), .A3(new_n534), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n630), .A2(new_n724), .A3(KEYINPUT30), .A4(new_n591), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n462), .A2(new_n595), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n534), .A2(new_n337), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT91), .B1(new_n605), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n605), .A2(new_n728), .A3(KEYINPUT91), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n727), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT31), .B(new_n678), .C1(new_n726), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n605), .A2(new_n728), .A3(KEYINPUT91), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n729), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n723), .B(new_n725), .C1(new_n736), .C2(new_n727), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT31), .B1(new_n737), .B2(new_n678), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n687), .B1(new_n719), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n718), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n702), .B1(new_n741), .B2(G1), .ZN(G364));
  INV_X1    g0542(.A(G13), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n207), .B1(new_n744), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n697), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n214), .B1(G20), .B2(new_n413), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n208), .A2(new_n395), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n330), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n208), .A2(G190), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G303), .A2(new_n754), .B1(new_n758), .B2(G329), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n755), .A2(new_n752), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n314), .B1(new_n761), .B2(G283), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n756), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n759), .B(new_n762), .C1(new_n763), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n336), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n751), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n208), .A2(new_n330), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n337), .A2(G190), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n770), .A2(G322), .B1(new_n773), .B2(G326), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n337), .A2(new_n395), .A3(new_n771), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT33), .B(G317), .Z(new_n776));
  OAI21_X1  g0576(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT97), .ZN(new_n778));
  AND3_X1   g0578(.A1(new_n768), .A2(new_n778), .A3(new_n755), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(new_n768), .B2(new_n755), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n767), .B(new_n777), .C1(G311), .C2(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n782), .A2(G77), .B1(G50), .B2(new_n773), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n769), .B(KEYINPUT96), .Z(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n258), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT98), .Z(new_n787));
  NAND2_X1  g0587(.A1(new_n754), .A2(G87), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n788), .B(new_n314), .C1(new_n398), .C2(new_n760), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n757), .A2(KEYINPUT32), .A3(new_n265), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G97), .B2(new_n765), .ZN(new_n791));
  OAI21_X1  g0591(.A(KEYINPUT32), .B1(new_n757), .B2(new_n265), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n775), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n789), .B(new_n793), .C1(G68), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n783), .B1(new_n796), .B2(KEYINPUT99), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT99), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n787), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n750), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n750), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT95), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n696), .A2(new_n251), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G355), .B1(new_n607), .B2(new_n696), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT94), .Z(new_n809));
  NAND2_X1  g0609(.A1(new_n283), .A2(new_n285), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n696), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n219), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(G45), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n243), .A2(new_n323), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n809), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n748), .B(new_n800), .C1(new_n806), .C2(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT100), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(KEYINPUT100), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(new_n686), .C2(new_n804), .ZN(new_n819));
  INV_X1    g0619(.A(new_n689), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n747), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n688), .B2(new_n686), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT93), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n819), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT101), .ZN(G396));
  NAND2_X1  g0627(.A1(new_n670), .A2(new_n703), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT102), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n416), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n415), .A2(new_n678), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n416), .A2(new_n829), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n830), .A2(new_n412), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n416), .A2(new_n703), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n828), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n830), .A2(new_n832), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n838), .A2(new_n412), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n839), .A2(new_n670), .A3(new_n703), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n740), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT103), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(new_n748), .C1(new_n740), .C2(new_n841), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G137), .A2(new_n773), .B1(new_n794), .B2(G150), .ZN(new_n845));
  INV_X1    g0645(.A(G143), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n265), .B2(new_n781), .C1(new_n785), .C2(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT34), .Z(new_n848));
  AOI22_X1  g0648(.A1(G50), .A2(new_n754), .B1(new_n758), .B2(G132), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n761), .A2(G68), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n765), .A2(G58), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n849), .A2(new_n810), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n314), .B1(new_n754), .B2(G107), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n765), .A2(G97), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n758), .A2(G311), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n761), .A2(G87), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n770), .A2(G294), .B1(new_n794), .B2(G283), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n602), .B2(new_n772), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n858), .B(new_n860), .C1(G116), .C2(new_n782), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n749), .B1(new_n853), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n749), .A2(new_n801), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n748), .B1(new_n410), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n862), .B(new_n864), .C1(new_n835), .C2(new_n802), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n844), .A2(new_n865), .ZN(G384));
  NAND2_X1  g0666(.A1(new_n215), .A2(G116), .ZN(new_n867));
  INV_X1    g0667(.A(new_n566), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(KEYINPUT35), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(KEYINPUT35), .B2(new_n868), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT36), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n261), .A2(new_n218), .A3(new_n410), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n288), .A2(G50), .ZN(new_n873));
  OAI211_X1 g0673(.A(G1), .B(new_n743), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT104), .ZN(new_n876));
  INV_X1    g0676(.A(new_n676), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n271), .B1(new_n297), .B2(KEYINPUT16), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n348), .B2(new_n347), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n877), .B1(new_n879), .B2(new_n310), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n346), .B1(new_n879), .B2(new_n310), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(new_n333), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n877), .B1(new_n349), .B2(new_n310), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n333), .A2(new_n350), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n880), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n355), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n393), .A2(new_n396), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n375), .A2(new_n703), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n393), .B(new_n396), .C1(new_n375), .C2(new_n703), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n838), .A2(new_n678), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT105), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n901), .B2(new_n840), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n893), .A2(new_n902), .B1(new_n640), .B2(new_n676), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n904));
  INV_X1    g0704(.A(new_n884), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n355), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n333), .A2(new_n350), .A3(new_n884), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n886), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT106), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n892), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT106), .A4(KEYINPUT38), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n904), .B1(new_n914), .B2(KEYINPUT39), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n393), .A2(new_n678), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n903), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT107), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n718), .B2(new_n445), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n711), .A2(new_n716), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(KEYINPUT29), .A3(new_n703), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT29), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n828), .A2(new_n922), .ZN(new_n923));
  AND4_X1   g0723(.A1(new_n918), .A2(new_n921), .A3(new_n923), .A4(new_n445), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n642), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n917), .B(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT40), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n890), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n719), .A2(new_n739), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT108), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n719), .A2(new_n739), .A3(KEYINPUT108), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n836), .B1(new_n897), .B2(new_n896), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n910), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n886), .A2(new_n883), .B1(new_n355), .B2(new_n888), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT106), .B1(new_n938), .B2(KEYINPUT38), .ZN(new_n939));
  AND4_X1   g0739(.A1(KEYINPUT106), .A2(new_n887), .A3(new_n889), .A4(KEYINPUT38), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n935), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n936), .B1(new_n943), .B2(KEYINPUT40), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n932), .A2(new_n445), .A3(new_n933), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n926), .B1(new_n946), .B2(new_n687), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n207), .B2(new_n744), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n926), .A2(new_n946), .A3(new_n687), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n876), .B1(new_n948), .B2(new_n949), .ZN(G367));
  NAND2_X1  g0750(.A1(new_n648), .A2(new_n654), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n524), .A2(new_n703), .ZN(new_n952));
  MUX2_X1   g0752(.A(new_n648), .B(new_n951), .S(new_n952), .Z(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n668), .B1(new_n593), .B2(new_n703), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT109), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n649), .A2(new_n678), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n692), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT42), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n680), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n658), .A2(new_n659), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n678), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n955), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n690), .A2(new_n959), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n968), .B(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n697), .B(KEYINPUT41), .Z(new_n972));
  INV_X1    g0772(.A(new_n690), .ZN(new_n973));
  INV_X1    g0773(.A(new_n959), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n693), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT44), .Z(new_n976));
  NOR2_X1   g0776(.A1(new_n974), .A2(new_n693), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT45), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n973), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n681), .B1(new_n682), .B2(new_n678), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n692), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n820), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n741), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n976), .A2(new_n973), .A3(new_n978), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n980), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n972), .B1(new_n987), .B2(new_n741), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n971), .B1(new_n988), .B2(new_n746), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n806), .B1(new_n211), .B2(new_n408), .ZN(new_n990));
  INV_X1    g0790(.A(new_n811), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n239), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n747), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT110), .Z(new_n994));
  INV_X1    g0794(.A(G150), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n769), .A2(new_n995), .B1(new_n775), .B2(new_n265), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G143), .B2(new_n773), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n760), .A2(new_n410), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G58), .B2(new_n754), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n765), .A2(G68), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n251), .B1(new_n758), .B2(G137), .ZN(new_n1001));
  AND3_X1   g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n997), .B(new_n1002), .C1(new_n371), .C2(new_n781), .ZN(new_n1003));
  INV_X1    g0803(.A(G283), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n785), .A2(new_n602), .B1(new_n781), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n754), .A2(G116), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT46), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1006), .A2(new_n1007), .B1(new_n398), .B2(new_n766), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n1007), .B2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n773), .A2(G311), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n794), .A2(G294), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n760), .A2(new_n515), .B1(new_n757), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1013), .A2(new_n810), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1003), .B1(new_n1005), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT47), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n750), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n994), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n954), .B2(new_n804), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT111), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n989), .A2(new_n1023), .ZN(G387));
  INV_X1    g0824(.A(new_n699), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n807), .A2(new_n1025), .B1(new_n398), .B2(new_n696), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n236), .A2(new_n323), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n301), .A2(G50), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT50), .Z(new_n1029));
  OAI211_X1 g0829(.A(new_n699), .B(new_n323), .C1(new_n288), .C2(new_n410), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n811), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1026), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n748), .B1(new_n1032), .B2(new_n806), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n754), .A2(G77), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n515), .B2(new_n760), .C1(new_n995), .C2(new_n757), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n769), .A2(new_n371), .B1(new_n772), .B2(new_n265), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n810), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n766), .A2(new_n408), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n288), .B2(new_n781), .C1(new_n306), .C2(new_n775), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT112), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G311), .A2(new_n794), .B1(new_n773), .B2(G322), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n602), .B2(new_n781), .C1(new_n785), .C2(new_n1012), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n754), .A2(G294), .B1(new_n765), .B2(G283), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT49), .Z(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT113), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n758), .A2(G326), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1037), .B(new_n1051), .C1(new_n607), .C2(new_n760), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n1049), .B2(KEYINPUT113), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1041), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1033), .B1(new_n1054), .B2(new_n750), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n681), .B2(new_n803), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n983), .B2(new_n746), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n983), .A2(new_n741), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n984), .A2(new_n697), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(G393));
  NAND3_X1  g0860(.A1(new_n980), .A2(new_n746), .A3(new_n986), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n806), .B1(new_n515), .B2(new_n211), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n991), .A2(new_n246), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n747), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n810), .B1(new_n766), .B2(new_n410), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n857), .B1(new_n846), .B2(new_n757), .C1(new_n222), .C2(new_n753), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G50), .C2(new_n794), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n769), .A2(new_n265), .B1(new_n772), .B2(new_n995), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(new_n301), .C2(new_n781), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n775), .A2(new_n602), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G283), .A2(new_n754), .B1(new_n758), .B2(G322), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1072), .B(new_n251), .C1(new_n398), .C2(new_n760), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(G116), .C2(new_n765), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n763), .B2(new_n781), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n770), .A2(G311), .B1(new_n773), .B2(G317), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1070), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1064), .B1(new_n1078), .B2(new_n749), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n959), .B2(new_n804), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1061), .A2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n987), .A2(new_n697), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n986), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n984), .B1(new_n1083), .B2(new_n979), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G390));
  NAND4_X1  g0886(.A1(new_n930), .A2(new_n688), .A3(new_n835), .A4(new_n898), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n900), .B1(new_n717), .B2(new_n839), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(new_n899), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n941), .A2(new_n1089), .A3(new_n916), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT39), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n928), .A2(new_n890), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n941), .B2(new_n1091), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n916), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n902), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1087), .B(new_n1090), .C1(new_n1093), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1095), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n914), .A2(new_n1094), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n915), .A2(new_n1097), .B1(new_n1098), .B2(new_n1089), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n932), .A2(new_n934), .A3(G330), .A4(new_n933), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1096), .B(new_n746), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n306), .A2(new_n863), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n781), .A2(new_n515), .B1(new_n398), .B2(new_n775), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n758), .A2(G294), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n788), .A2(new_n850), .A3(new_n1106), .A4(new_n251), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n769), .A2(new_n607), .B1(new_n772), .B2(new_n1004), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(G77), .C2(new_n765), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1104), .A2(new_n1105), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT117), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n251), .B1(new_n761), .B2(G50), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n758), .A2(G125), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(new_n265), .C2(new_n766), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n753), .A2(new_n995), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT115), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1115), .B1(KEYINPUT53), .B2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n782), .A2(new_n1120), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1117), .A2(KEYINPUT53), .ZN(new_n1122));
  INV_X1    g0922(.A(G132), .ZN(new_n1123));
  INV_X1    g0923(.A(G128), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n769), .A2(new_n1123), .B1(new_n772), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G137), .B2(new_n794), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1112), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n748), .B(new_n1102), .C1(new_n1129), .C2(new_n749), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT118), .Z(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1093), .B2(new_n802), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1101), .A2(KEYINPUT119), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT119), .B1(new_n1101), .B2(new_n1132), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n901), .A2(new_n840), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n740), .A2(new_n835), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n899), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1100), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n932), .A2(G330), .A3(new_n835), .A4(new_n933), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n899), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1088), .A2(new_n1087), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1136), .A2(new_n1139), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n932), .A2(new_n445), .A3(G330), .A4(new_n933), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n642), .B(new_n1144), .C1(new_n919), .C2(new_n924), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1146), .B(new_n1096), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1147), .A2(new_n697), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT114), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1090), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1100), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1149), .B(new_n1146), .C1(new_n1152), .C2(new_n1096), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1146), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT114), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1148), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1135), .A2(new_n1157), .ZN(G378));
  INV_X1    g0958(.A(KEYINPUT123), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n425), .A2(new_n676), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n444), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n435), .A2(new_n441), .A3(new_n443), .A4(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1164), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1159), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(KEYINPUT123), .A3(new_n1165), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n802), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n748), .B1(new_n371), .B2(new_n863), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n770), .A2(G107), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT121), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n408), .B2(new_n781), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n761), .A2(G58), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT120), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n515), .B2(new_n775), .C1(new_n607), .C2(new_n772), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1037), .A2(new_n322), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1034), .B(new_n1000), .C1(new_n1004), .C2(new_n757), .ZN(new_n1180));
  NOR4_X1   g0980(.A1(new_n1175), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1179), .B(new_n371), .C1(G33), .C2(G41), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n770), .A2(G128), .B1(new_n773), .B2(G125), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n754), .A2(new_n1120), .B1(new_n765), .B2(G150), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n1123), .C2(new_n775), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G137), .B2(new_n782), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT122), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G33), .B(G41), .C1(new_n758), .C2(G124), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n265), .B2(new_n760), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1190), .B2(KEYINPUT59), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1185), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1172), .B1(new_n1195), .B2(new_n750), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1171), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n917), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1169), .A2(new_n1165), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT124), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(KEYINPUT40), .B1(new_n914), .B2(new_n935), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n942), .A2(new_n893), .A3(new_n927), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1201), .B1(new_n1204), .B2(G330), .ZN(new_n1205));
  INV_X1    g1005(.A(G330), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1169), .A2(KEYINPUT123), .A3(KEYINPUT124), .A4(new_n1165), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1168), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1206), .B(new_n1209), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1198), .B1(new_n1205), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n927), .B1(new_n941), .B2(new_n942), .ZN(new_n1212));
  OAI211_X1 g1012(.A(G330), .B(new_n1208), .C1(new_n1212), .C2(new_n936), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1206), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n917), .C1(new_n1214), .C2(new_n1201), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1197), .B1(new_n1216), .B2(new_n746), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1145), .B(KEYINPUT125), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1147), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1215), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n944), .A2(new_n1206), .B1(new_n1200), .B2(new_n1199), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n917), .B1(new_n1221), .B2(new_n1213), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1219), .B(KEYINPUT57), .C1(new_n1220), .C2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n697), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1211), .A2(new_n1215), .B1(new_n1147), .B2(new_n1218), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT57), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1217), .B1(new_n1224), .B2(new_n1226), .ZN(G375));
  NOR2_X1   g1027(.A1(new_n1146), .A2(new_n972), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1143), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1145), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1177), .B1(new_n1123), .B2(new_n772), .C1(new_n775), .C2(new_n1119), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n766), .A2(new_n371), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n753), .A2(new_n265), .B1(new_n757), .B2(new_n1124), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1232), .A2(new_n1037), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(G137), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1235), .B1(new_n1236), .B2(new_n785), .C1(new_n995), .C2(new_n781), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n607), .A2(new_n775), .B1(new_n772), .B2(new_n763), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G283), .B2(new_n770), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n753), .A2(new_n515), .B1(new_n757), .B2(new_n602), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1038), .A2(new_n1240), .A3(new_n314), .A4(new_n998), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1239), .B(new_n1241), .C1(new_n398), .C2(new_n781), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n750), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n748), .B(new_n1243), .C1(new_n288), .C2(new_n863), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n802), .B2(new_n898), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1143), .B2(new_n745), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1231), .A2(new_n1247), .ZN(G381));
  NAND3_X1  g1048(.A1(new_n989), .A2(new_n1085), .A3(new_n1023), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G375), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1101), .A2(new_n1132), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1157), .A2(new_n1252), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1251), .A3(new_n1253), .A4(new_n1254), .ZN(G407));
  INV_X1    g1055(.A(G213), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(G343), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1251), .A2(new_n1253), .A3(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(G407), .A2(G213), .A3(new_n1258), .ZN(G409));
  OAI211_X1 g1059(.A(G378), .B(new_n1217), .C1(new_n1226), .C2(new_n1224), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1217), .B1(new_n972), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1253), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1257), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT126), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1155), .B(new_n697), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1247), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT127), .B1(new_n844), .B2(new_n865), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(G384), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1272), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n1247), .B1(G384), .B2(new_n1274), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(G2897), .A3(new_n1257), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1257), .A2(G2897), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1276), .A2(new_n1277), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT61), .B1(new_n1266), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1266), .B2(new_n1278), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G396), .B(G393), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1085), .B1(new_n989), .B2(new_n1023), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1250), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(G390), .ZN(new_n1290));
  XOR2_X1   g1090(.A(G396), .B(G393), .Z(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1249), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1257), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1278), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(KEYINPUT63), .A3(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1284), .A2(new_n1286), .A3(new_n1293), .A4(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT62), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1294), .A2(new_n1298), .A3(new_n1295), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1294), .B2(new_n1282), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1298), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1299), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1297), .B1(new_n1303), .B2(new_n1293), .ZN(G405));
  AND2_X1   g1104(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1305));
  AND2_X1   g1105(.A1(G375), .A2(new_n1253), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1260), .ZN(new_n1307));
  OR3_X1    g1107(.A1(new_n1306), .A2(new_n1307), .A3(new_n1295), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1295), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1305), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1305), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(G402));
endmodule


