// Benchmark "locked_c3540" written by ABC on Sat Dec 16 11:14:46 2023

module locked_c3540 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41,
    G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132,
    G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226,
    G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311,
    G317, G322, G326, G329, G330, G343, G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13,
    G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124,
    G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213,
    G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283,
    G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n137, new_n138, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n163, new_n165, new_n166, new_n167,
    new_n168, new_n169, new_n170, new_n171, new_n173, new_n174, new_n175,
    new_n176, new_n177, new_n178, new_n179, new_n181, new_n182, new_n183,
    new_n184, new_n185, new_n186, new_n187, new_n188, new_n189, new_n190,
    new_n191, new_n192, new_n193, new_n194, new_n195, new_n196, new_n197,
    new_n198, new_n199, new_n200, new_n201, new_n202, new_n203, new_n204,
    new_n205, new_n206, new_n207, new_n208, new_n209, new_n210, new_n211,
    new_n212, new_n213, new_n214, new_n215, new_n216, new_n217, new_n218,
    new_n219, new_n220, new_n221, new_n222, new_n223, new_n224, new_n225,
    new_n226, new_n227, new_n228, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n303, new_n304, new_n305, new_n306, new_n307, new_n308, new_n309,
    new_n310, new_n311, new_n312, new_n313, new_n314, new_n315, new_n316,
    new_n317, new_n318, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n409, new_n410, new_n411, new_n412, new_n413, new_n414,
    new_n415, new_n416, new_n417, new_n418, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n425, new_n426, new_n427, new_n428,
    new_n429, new_n430, new_n431, new_n432, new_n433, new_n434, new_n435,
    new_n436, new_n437, new_n438, new_n439, new_n440, new_n441, new_n442,
    new_n443, new_n444, new_n445, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n451, new_n452, new_n453, new_n454, new_n455, new_n456,
    new_n457, new_n458, new_n459, new_n460, new_n461, new_n462, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009;
  NOR3_X1   g000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n137));
  INV_X1    g001(.A(G77), .ZN(new_n138));
  AND2_X1   g002(.A1(new_n137), .A2(new_n138), .ZN(G353));
  OAI21_X1  g003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g004(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n141));
  NAND2_X1  g005(.A1(G77), .A2(G244), .ZN(new_n142));
  INV_X1    g006(.A(G68), .ZN(new_n143));
  INV_X1    g007(.A(G238), .ZN(new_n144));
  OAI211_X1 g008(.A(new_n141), .B(new_n142), .C1(new_n143), .C2(new_n144), .ZN(new_n145));
  AOI21_X1  g009(.A(new_n145), .B1(G50), .B2(G226), .ZN(new_n146));
  NAND2_X1  g010(.A1(G107), .A2(G264), .ZN(new_n147));
  NAND2_X1  g011(.A1(G116), .A2(G270), .ZN(new_n148));
  NAND2_X1  g012(.A1(G87), .A2(G250), .ZN(new_n149));
  NAND4_X1  g013(.A1(new_n146), .A2(new_n147), .A3(new_n148), .A4(new_n149), .ZN(new_n150));
  NAND2_X1  g014(.A1(G1), .A2(G20), .ZN(new_n151));
  NAND2_X1  g015(.A1(new_n150), .A2(new_n151), .ZN(new_n152));
  NAND2_X1  g016(.A1(G1), .A2(G13), .ZN(new_n153));
  INV_X1    g017(.A(new_n153), .ZN(new_n154));
  NOR2_X1   g018(.A1(new_n154), .A2(new_n151), .ZN(new_n155));
  OAI211_X1 g019(.A(new_n155), .B(G250), .C1(G257), .C2(G264), .ZN(new_n156));
  INV_X1    g020(.A(new_n156), .ZN(new_n157));
  OAI22_X1  g021(.A1(new_n152), .A2(KEYINPUT1), .B1(KEYINPUT0), .B2(new_n157), .ZN(new_n158));
  AND2_X1   g022(.A1(new_n152), .A2(KEYINPUT1), .ZN(new_n159));
  AND2_X1   g023(.A1(new_n157), .A2(KEYINPUT0), .ZN(new_n160));
  OAI21_X1  g024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n161));
  INV_X1    g025(.A(G20), .ZN(new_n162));
  NOR3_X1   g026(.A1(new_n161), .A2(new_n162), .A3(new_n153), .ZN(new_n163));
  NOR4_X1   g027(.A1(new_n158), .A2(new_n159), .A3(new_n160), .A4(new_n163), .ZN(G361));
  XOR2_X1   g028(.A(G264), .B(G270), .Z(new_n165));
  XNOR2_X1  g029(.A(new_n165), .B(G250), .ZN(new_n166));
  XNOR2_X1  g030(.A(new_n166), .B(G257), .ZN(new_n167));
  XNOR2_X1  g031(.A(G238), .B(G244), .ZN(new_n168));
  XNOR2_X1  g032(.A(new_n168), .B(G232), .ZN(new_n169));
  XNOR2_X1  g033(.A(KEYINPUT2), .B(G226), .ZN(new_n170));
  XNOR2_X1  g034(.A(new_n169), .B(new_n170), .ZN(new_n171));
  XNOR2_X1  g035(.A(new_n167), .B(new_n171), .ZN(G358));
  XNOR2_X1  g036(.A(G87), .B(G97), .ZN(new_n173));
  INV_X1    g037(.A(G107), .ZN(new_n174));
  XNOR2_X1  g038(.A(new_n173), .B(new_n174), .ZN(new_n175));
  XNOR2_X1  g039(.A(new_n175), .B(G116), .ZN(new_n176));
  XOR2_X1   g040(.A(G68), .B(G77), .Z(new_n177));
  XNOR2_X1  g041(.A(G50), .B(G58), .ZN(new_n178));
  XNOR2_X1  g042(.A(new_n177), .B(new_n178), .ZN(new_n179));
  XNOR2_X1  g043(.A(new_n176), .B(new_n179), .ZN(G351));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G33), .ZN(new_n181));
  INV_X1    g045(.A(G1698), .ZN(new_n182));
  NAND3_X1  g046(.A1(new_n181), .A2(G226), .A3(new_n182), .ZN(new_n183));
  NAND2_X1  g047(.A1(G33), .A2(G97), .ZN(new_n184));
  NAND2_X1  g048(.A1(new_n181), .A2(G1698), .ZN(new_n185));
  INV_X1    g049(.A(G232), .ZN(new_n186));
  OAI211_X1 g050(.A(new_n183), .B(new_n184), .C1(new_n185), .C2(new_n186), .ZN(new_n187));
  AOI21_X1  g051(.A(new_n153), .B1(G33), .B2(G41), .ZN(new_n188));
  NAND2_X1  g052(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g053(.A(KEYINPUT13), .ZN(new_n190));
  INV_X1    g054(.A(G41), .ZN(new_n191));
  INV_X1    g055(.A(G45), .ZN(new_n192));
  AOI21_X1  g056(.A(G1), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g057(.A1(new_n193), .A2(G274), .ZN(new_n194));
  INV_X1    g058(.A(new_n194), .ZN(new_n195));
  NOR2_X1   g059(.A1(new_n188), .A2(new_n193), .ZN(new_n196));
  AOI21_X1  g060(.A(new_n195), .B1(new_n196), .B2(G238), .ZN(new_n197));
  NAND3_X1  g061(.A1(new_n189), .A2(new_n190), .A3(new_n197), .ZN(new_n198));
  INV_X1    g062(.A(new_n198), .ZN(new_n199));
  AOI21_X1  g063(.A(new_n190), .B1(new_n189), .B2(new_n197), .ZN(new_n200));
  OAI21_X1  g064(.A(G169), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g065(.A1(new_n201), .A2(KEYINPUT14), .ZN(new_n202));
  INV_X1    g066(.A(new_n200), .ZN(new_n203));
  NAND2_X1  g067(.A1(new_n203), .A2(new_n198), .ZN(new_n204));
  INV_X1    g068(.A(KEYINPUT14), .ZN(new_n205));
  NAND3_X1  g069(.A1(new_n204), .A2(new_n205), .A3(G169), .ZN(new_n206));
  NAND3_X1  g070(.A1(new_n203), .A2(G179), .A3(new_n198), .ZN(new_n207));
  NAND3_X1  g071(.A1(new_n202), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g072(.A1(new_n143), .A2(G20), .ZN(new_n209));
  NAND2_X1  g073(.A1(new_n162), .A2(G33), .ZN(new_n210));
  NOR2_X1   g074(.A1(G20), .A2(G33), .ZN(new_n211));
  INV_X1    g075(.A(new_n211), .ZN(new_n212));
  INV_X1    g076(.A(G50), .ZN(new_n213));
  OAI221_X1 g077(.A(new_n209), .B1(new_n210), .B2(new_n138), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND3_X1  g078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n215));
  NAND2_X1  g079(.A1(new_n215), .A2(new_n153), .ZN(new_n216));
  NAND2_X1  g080(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g081(.A(new_n217), .B(KEYINPUT11), .ZN(new_n218));
  INV_X1    g082(.A(new_n216), .ZN(new_n219));
  OAI21_X1  g083(.A(new_n219), .B1(G1), .B2(new_n162), .ZN(new_n220));
  INV_X1    g084(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g085(.A1(new_n221), .A2(G68), .ZN(new_n222));
  INV_X1    g086(.A(G13), .ZN(new_n223));
  NOR2_X1   g087(.A1(new_n223), .A2(G1), .ZN(new_n224));
  INV_X1    g088(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g089(.A1(new_n225), .A2(new_n209), .ZN(new_n226));
  XOR2_X1   g090(.A(new_n226), .B(KEYINPUT12), .Z(new_n227));
  NAND3_X1  g091(.A1(new_n218), .A2(new_n222), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g092(.A1(new_n208), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g093(.A1(new_n204), .A2(G200), .ZN(new_n230));
  INV_X1    g094(.A(new_n228), .ZN(new_n231));
  NAND3_X1  g095(.A1(new_n203), .A2(G190), .A3(new_n198), .ZN(new_n232));
  AND3_X1   g096(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g097(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g098(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  INV_X1    g099(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g100(.A1(new_n181), .A2(G223), .A3(G1698), .ZN(new_n237));
  NAND2_X1  g101(.A1(new_n181), .A2(new_n182), .ZN(new_n238));
  INV_X1    g102(.A(G222), .ZN(new_n239));
  OAI221_X1 g103(.A(new_n237), .B1(new_n138), .B2(new_n181), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g104(.A1(new_n240), .A2(new_n188), .ZN(new_n241));
  AOI21_X1  g105(.A(new_n195), .B1(new_n196), .B2(G226), .ZN(new_n242));
  AND2_X1   g106(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g107(.A(KEYINPUT9), .ZN(new_n244));
  NAND2_X1  g108(.A1(new_n211), .A2(G150), .ZN(new_n245));
  XNOR2_X1  g109(.A(KEYINPUT8), .B(G58), .ZN(new_n246));
  OAI221_X1 g110(.A(new_n245), .B1(new_n137), .B2(new_n162), .C1(new_n246), .C2(new_n210), .ZN(new_n247));
  NOR3_X1   g111(.A1(new_n223), .A2(new_n162), .A3(G1), .ZN(new_n248));
  AOI22_X1  g112(.A1(new_n247), .A2(new_n216), .B1(new_n213), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g113(.A(new_n249), .B1(new_n213), .B2(new_n220), .ZN(new_n250));
  AOI22_X1  g114(.A1(new_n243), .A2(G190), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  INV_X1    g115(.A(G200), .ZN(new_n252));
  OAI221_X1 g116(.A(new_n251), .B1(new_n244), .B2(new_n250), .C1(new_n252), .C2(new_n243), .ZN(new_n253));
  XNOR2_X1  g117(.A(new_n253), .B(KEYINPUT10), .ZN(new_n254));
  OAI21_X1  g118(.A(new_n250), .B1(new_n243), .B2(G169), .ZN(new_n255));
  INV_X1    g119(.A(G179), .ZN(new_n256));
  AOI21_X1  g120(.A(new_n255), .B1(new_n256), .B2(new_n243), .ZN(new_n257));
  INV_X1    g121(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g122(.A1(new_n236), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  INV_X1    g123(.A(G33), .ZN(new_n260));
  NAND2_X1  g124(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g126(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND2_X1  g127(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g128(.A(KEYINPUT7), .B1(new_n264), .B2(new_n162), .ZN(new_n265));
  INV_X1    g129(.A(KEYINPUT7), .ZN(new_n266));
  AOI211_X1 g130(.A(new_n266), .B(G20), .C1(new_n261), .C2(new_n263), .ZN(new_n267));
  OAI21_X1  g131(.A(G68), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g132(.A(G58), .ZN(new_n269));
  NOR2_X1   g133(.A1(new_n269), .A2(new_n143), .ZN(new_n270));
  NOR2_X1   g134(.A1(G58), .A2(G68), .ZN(new_n271));
  OAI21_X1  g135(.A(G20), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g136(.A1(new_n211), .A2(G159), .ZN(new_n273));
  NAND2_X1  g137(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g138(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g139(.A1(new_n268), .A2(KEYINPUT16), .A3(new_n275), .ZN(new_n276));
  INV_X1    g140(.A(KEYINPUT16), .ZN(new_n277));
  OAI21_X1  g141(.A(new_n266), .B1(new_n181), .B2(G20), .ZN(new_n278));
  NOR2_X1   g142(.A1(new_n262), .A2(G33), .ZN(new_n279));
  NOR2_X1   g143(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n280));
  OAI211_X1 g144(.A(KEYINPUT7), .B(new_n162), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AOI21_X1  g145(.A(new_n143), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g146(.A(new_n277), .B1(new_n282), .B2(new_n274), .ZN(new_n283));
  NAND3_X1  g147(.A1(new_n276), .A2(new_n283), .A3(new_n216), .ZN(new_n284));
  INV_X1    g148(.A(new_n246), .ZN(new_n285));
  NAND2_X1  g149(.A1(new_n221), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g150(.A1(new_n246), .A2(new_n248), .ZN(new_n287));
  NAND3_X1  g151(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND4_X1  g152(.A1(new_n261), .A2(new_n263), .A3(G226), .A4(G1698), .ZN(new_n289));
  NAND4_X1  g153(.A1(new_n261), .A2(new_n263), .A3(G223), .A4(new_n182), .ZN(new_n290));
  INV_X1    g154(.A(G87), .ZN(new_n291));
  OAI211_X1 g155(.A(new_n289), .B(new_n290), .C1(new_n260), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g156(.A1(new_n292), .A2(new_n188), .ZN(new_n293));
  NAND2_X1  g157(.A1(new_n196), .A2(G232), .ZN(new_n294));
  NAND3_X1  g158(.A1(new_n293), .A2(new_n194), .A3(new_n294), .ZN(new_n295));
  INV_X1    g159(.A(G169), .ZN(new_n296));
  NAND2_X1  g160(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g161(.A1(new_n295), .A2(G179), .ZN(new_n298));
  NAND3_X1  g162(.A1(new_n288), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g163(.A(KEYINPUT18), .ZN(new_n300));
  NAND2_X1  g164(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g165(.A1(new_n288), .A2(KEYINPUT18), .A3(new_n297), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g166(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND3_X1   g167(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n304));
  INV_X1    g168(.A(KEYINPUT17), .ZN(new_n305));
  INV_X1    g169(.A(G190), .ZN(new_n306));
  NOR2_X1   g170(.A1(new_n295), .A2(new_n306), .ZN(new_n307));
  INV_X1    g171(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g172(.A1(new_n295), .A2(G200), .ZN(new_n309));
  NAND4_X1  g173(.A1(new_n304), .A2(new_n305), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  NAND4_X1  g174(.A1(new_n284), .A2(new_n309), .A3(new_n286), .A4(new_n287), .ZN(new_n311));
  OAI21_X1  g175(.A(KEYINPUT17), .B1(new_n311), .B2(new_n307), .ZN(new_n312));
  NAND2_X1  g176(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g177(.A1(G20), .A2(G77), .ZN(new_n314));
  XNOR2_X1  g178(.A(KEYINPUT15), .B(G87), .ZN(new_n315));
  OAI221_X1 g179(.A(new_n314), .B1(new_n315), .B2(new_n210), .C1(new_n212), .C2(new_n246), .ZN(new_n316));
  AOI22_X1  g180(.A1(new_n316), .A2(new_n216), .B1(new_n138), .B2(new_n248), .ZN(new_n317));
  NAND2_X1  g181(.A1(new_n221), .A2(G77), .ZN(new_n318));
  NAND2_X1  g182(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI22_X1  g183(.A1(new_n186), .A2(new_n238), .B1(new_n185), .B2(new_n144), .ZN(new_n320));
  NOR2_X1   g184(.A1(new_n181), .A2(new_n174), .ZN(new_n321));
  OAI21_X1  g185(.A(new_n188), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g186(.A(new_n195), .B1(new_n196), .B2(G244), .ZN(new_n323));
  NAND2_X1  g187(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g188(.A1(new_n324), .A2(new_n256), .ZN(new_n325));
  AOI21_X1  g189(.A(new_n296), .B1(new_n322), .B2(new_n323), .ZN(new_n326));
  OAI21_X1  g190(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g191(.A1(new_n324), .A2(G200), .ZN(new_n328));
  INV_X1    g192(.A(new_n319), .ZN(new_n329));
  OAI211_X1 g193(.A(new_n328), .B(new_n329), .C1(new_n306), .C2(new_n324), .ZN(new_n330));
  NAND4_X1  g194(.A1(new_n303), .A2(new_n313), .A3(new_n327), .A4(new_n330), .ZN(new_n331));
  NOR2_X1   g195(.A1(new_n259), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g196(.A1(new_n261), .A2(new_n263), .A3(new_n162), .A4(G87), .ZN(new_n333));
  NAND2_X1  g197(.A1(new_n333), .A2(KEYINPUT22), .ZN(new_n334));
  INV_X1    g198(.A(KEYINPUT22), .ZN(new_n335));
  NAND4_X1  g199(.A1(new_n181), .A2(new_n335), .A3(new_n162), .A4(G87), .ZN(new_n336));
  NAND2_X1  g200(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g201(.A1(new_n162), .A2(G33), .A3(G116), .ZN(new_n338));
  NAND2_X1  g202(.A1(new_n174), .A2(G20), .ZN(new_n339));
  XOR2_X1   g203(.A(new_n339), .B(KEYINPUT23), .Z(new_n340));
  NAND3_X1  g204(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g205(.A(KEYINPUT24), .ZN(new_n342));
  NAND2_X1  g206(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g207(.A1(new_n337), .A2(KEYINPUT24), .A3(new_n338), .A4(new_n340), .ZN(new_n344));
  NAND3_X1  g208(.A1(new_n343), .A2(new_n216), .A3(new_n344), .ZN(new_n345));
  INV_X1    g209(.A(G1), .ZN(new_n346));
  NAND2_X1  g210(.A1(new_n346), .A2(G33), .ZN(new_n347));
  NAND3_X1  g211(.A1(new_n347), .A2(new_n153), .A3(new_n215), .ZN(new_n348));
  NOR2_X1   g212(.A1(new_n348), .A2(new_n248), .ZN(new_n349));
  NAND2_X1  g213(.A1(new_n349), .A2(G107), .ZN(new_n350));
  NOR2_X1   g214(.A1(new_n225), .A2(new_n339), .ZN(new_n351));
  XNOR2_X1  g215(.A(new_n351), .B(KEYINPUT25), .ZN(new_n352));
  NAND3_X1  g216(.A1(new_n345), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g217(.A1(new_n181), .A2(G250), .A3(new_n182), .ZN(new_n354));
  NAND3_X1  g218(.A1(new_n181), .A2(G257), .A3(G1698), .ZN(new_n355));
  NAND2_X1  g219(.A1(G33), .A2(G294), .ZN(new_n356));
  NAND3_X1  g220(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g221(.A1(new_n357), .A2(new_n188), .ZN(new_n358));
  NAND2_X1  g222(.A1(new_n346), .A2(G45), .ZN(new_n359));
  INV_X1    g223(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g224(.A1(new_n360), .A2(G274), .ZN(new_n361));
  INV_X1    g225(.A(new_n361), .ZN(new_n362));
  XNOR2_X1  g226(.A(KEYINPUT5), .B(G41), .ZN(new_n363));
  NAND2_X1  g227(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g228(.A(new_n188), .B1(new_n363), .B2(new_n360), .ZN(new_n365));
  NAND2_X1  g229(.A1(new_n365), .A2(G264), .ZN(new_n366));
  NAND3_X1  g230(.A1(new_n358), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g231(.A1(new_n367), .A2(G169), .ZN(new_n368));
  OAI21_X1  g232(.A(new_n368), .B1(new_n256), .B2(new_n367), .ZN(new_n369));
  NAND2_X1  g233(.A1(new_n353), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g234(.A1(new_n367), .A2(new_n306), .ZN(new_n371));
  NAND2_X1  g235(.A1(new_n367), .A2(G200), .ZN(new_n372));
  NAND4_X1  g236(.A1(new_n345), .A2(new_n372), .A3(new_n350), .A4(new_n352), .ZN(new_n373));
  OAI21_X1  g237(.A(new_n370), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g238(.A1(new_n315), .A2(new_n248), .ZN(new_n375));
  NAND4_X1  g239(.A1(new_n261), .A2(new_n263), .A3(new_n162), .A4(G68), .ZN(new_n376));
  INV_X1    g240(.A(KEYINPUT19), .ZN(new_n377));
  INV_X1    g241(.A(G97), .ZN(new_n378));
  OAI21_X1  g242(.A(new_n377), .B1(new_n210), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g243(.A1(new_n291), .A2(new_n378), .A3(new_n174), .ZN(new_n380));
  NAND2_X1  g244(.A1(new_n380), .A2(G20), .ZN(new_n381));
  NAND4_X1  g245(.A1(new_n162), .A2(KEYINPUT19), .A3(G33), .A4(G97), .ZN(new_n382));
  NAND4_X1  g246(.A1(new_n376), .A2(new_n379), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  AOI21_X1  g247(.A(new_n375), .B1(new_n383), .B2(new_n216), .ZN(new_n384));
  INV_X1    g248(.A(new_n349), .ZN(new_n385));
  OAI21_X1  g249(.A(new_n384), .B1(new_n385), .B2(new_n315), .ZN(new_n386));
  NAND4_X1  g250(.A1(new_n261), .A2(new_n263), .A3(G238), .A4(new_n182), .ZN(new_n387));
  NAND4_X1  g251(.A1(new_n261), .A2(new_n263), .A3(G244), .A4(G1698), .ZN(new_n388));
  INV_X1    g252(.A(G116), .ZN(new_n389));
  OAI211_X1 g253(.A(new_n387), .B(new_n388), .C1(new_n260), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g254(.A1(new_n390), .A2(new_n188), .ZN(new_n391));
  NOR2_X1   g255(.A1(new_n260), .A2(new_n191), .ZN(new_n392));
  OAI211_X1 g256(.A(new_n359), .B(G250), .C1(new_n392), .C2(new_n153), .ZN(new_n393));
  NAND4_X1  g257(.A1(new_n391), .A2(new_n256), .A3(new_n361), .A4(new_n393), .ZN(new_n394));
  INV_X1    g258(.A(new_n393), .ZN(new_n395));
  AOI211_X1 g259(.A(new_n362), .B(new_n395), .C1(new_n390), .C2(new_n188), .ZN(new_n396));
  OAI211_X1 g260(.A(new_n386), .B(new_n394), .C1(new_n396), .C2(G169), .ZN(new_n397));
  NOR3_X1   g261(.A1(new_n348), .A2(new_n248), .A3(new_n291), .ZN(new_n398));
  AOI211_X1 g262(.A(new_n375), .B(new_n398), .C1(new_n216), .C2(new_n383), .ZN(new_n399));
  NAND4_X1  g263(.A1(new_n391), .A2(G190), .A3(new_n361), .A4(new_n393), .ZN(new_n400));
  OAI211_X1 g264(.A(new_n399), .B(new_n400), .C1(new_n396), .C2(new_n252), .ZN(new_n401));
  AND2_X1   g265(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g266(.A1(new_n261), .A2(new_n263), .A3(G244), .A4(new_n182), .ZN(new_n403));
  INV_X1    g267(.A(KEYINPUT4), .ZN(new_n404));
  NAND2_X1  g268(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g269(.A1(new_n181), .A2(KEYINPUT4), .A3(G244), .A4(new_n182), .ZN(new_n406));
  NAND2_X1  g270(.A1(G33), .A2(G283), .ZN(new_n407));
  NAND3_X1  g271(.A1(new_n181), .A2(G250), .A3(G1698), .ZN(new_n408));
  NAND4_X1  g272(.A1(new_n405), .A2(new_n406), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g273(.A1(new_n409), .A2(new_n188), .ZN(new_n410));
  NAND2_X1  g274(.A1(new_n365), .A2(G257), .ZN(new_n411));
  AND2_X1   g275(.A1(new_n411), .A2(new_n364), .ZN(new_n412));
  NAND3_X1  g276(.A1(new_n410), .A2(G190), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g277(.A1(new_n412), .A2(new_n410), .ZN(new_n414));
  NAND2_X1  g278(.A1(new_n414), .A2(G200), .ZN(new_n415));
  NAND2_X1  g279(.A1(new_n224), .A2(G20), .ZN(new_n416));
  NOR2_X1   g280(.A1(new_n416), .A2(G97), .ZN(new_n417));
  INV_X1    g281(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g282(.A1(new_n385), .A2(new_n378), .ZN(new_n419));
  OAI21_X1  g283(.A(G107), .B1(new_n265), .B2(new_n267), .ZN(new_n420));
  NAND3_X1  g284(.A1(new_n174), .A2(KEYINPUT6), .A3(G97), .ZN(new_n421));
  NOR2_X1   g285(.A1(new_n378), .A2(new_n174), .ZN(new_n422));
  NOR2_X1   g286(.A1(G97), .A2(G107), .ZN(new_n423));
  NOR2_X1   g287(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g288(.A(new_n421), .B1(new_n424), .B2(KEYINPUT6), .ZN(new_n425));
  NAND2_X1  g289(.A1(new_n425), .A2(G20), .ZN(new_n426));
  NAND2_X1  g290(.A1(new_n211), .A2(G77), .ZN(new_n427));
  NAND3_X1  g291(.A1(new_n420), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g292(.A(new_n419), .B1(new_n428), .B2(new_n216), .ZN(new_n429));
  NAND4_X1  g293(.A1(new_n413), .A2(new_n415), .A3(new_n418), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g294(.A1(new_n428), .A2(new_n216), .ZN(new_n431));
  INV_X1    g295(.A(new_n419), .ZN(new_n432));
  NAND3_X1  g296(.A1(new_n431), .A2(new_n418), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g297(.A1(new_n414), .A2(new_n296), .ZN(new_n434));
  NAND3_X1  g298(.A1(new_n412), .A2(new_n256), .A3(new_n410), .ZN(new_n435));
  NAND3_X1  g299(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g300(.A1(new_n402), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g301(.A1(new_n261), .A2(new_n263), .A3(G264), .A4(G1698), .ZN(new_n438));
  NAND4_X1  g302(.A1(new_n261), .A2(new_n263), .A3(G257), .A4(new_n182), .ZN(new_n439));
  INV_X1    g303(.A(G303), .ZN(new_n440));
  OAI211_X1 g304(.A(new_n438), .B(new_n439), .C1(new_n440), .C2(new_n181), .ZN(new_n441));
  NAND2_X1  g305(.A1(new_n441), .A2(new_n188), .ZN(new_n442));
  NAND2_X1  g306(.A1(new_n365), .A2(G270), .ZN(new_n443));
  NAND3_X1  g307(.A1(new_n442), .A2(new_n443), .A3(new_n364), .ZN(new_n444));
  NAND2_X1  g308(.A1(new_n444), .A2(G200), .ZN(new_n445));
  NAND2_X1  g309(.A1(new_n349), .A2(G116), .ZN(new_n446));
  NAND2_X1  g310(.A1(new_n248), .A2(new_n389), .ZN(new_n447));
  AOI22_X1  g311(.A1(new_n215), .A2(new_n153), .B1(G20), .B2(new_n389), .ZN(new_n448));
  OAI211_X1 g312(.A(new_n407), .B(new_n162), .C1(G33), .C2(new_n378), .ZN(new_n449));
  AND3_X1   g313(.A1(new_n448), .A2(KEYINPUT20), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g314(.A(KEYINPUT20), .B1(new_n448), .B2(new_n449), .ZN(new_n451));
  OAI211_X1 g315(.A(new_n446), .B(new_n447), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g316(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g317(.A(new_n445), .B(new_n453), .C1(new_n306), .C2(new_n444), .ZN(new_n454));
  INV_X1    g318(.A(new_n444), .ZN(new_n455));
  NAND3_X1  g319(.A1(new_n455), .A2(G179), .A3(new_n452), .ZN(new_n456));
  NAND4_X1  g320(.A1(new_n444), .A2(KEYINPUT21), .A3(G169), .A4(new_n452), .ZN(new_n457));
  NAND3_X1  g321(.A1(new_n444), .A2(G169), .A3(new_n452), .ZN(new_n458));
  INV_X1    g322(.A(KEYINPUT21), .ZN(new_n459));
  NAND2_X1  g323(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g324(.A1(new_n454), .A2(new_n456), .A3(new_n457), .A4(new_n460), .ZN(new_n461));
  NOR3_X1   g325(.A1(new_n374), .A2(new_n437), .A3(new_n461), .ZN(new_n462));
  AND2_X1   g326(.A1(new_n332), .A2(new_n462), .ZN(G372));
  NAND3_X1  g327(.A1(new_n460), .A2(new_n456), .A3(new_n457), .ZN(new_n464));
  OAI21_X1  g328(.A(new_n464), .B1(new_n371), .B2(new_n373), .ZN(new_n465));
  NAND2_X1  g329(.A1(new_n465), .A2(new_n370), .ZN(new_n466));
  INV_X1    g330(.A(new_n437), .ZN(new_n467));
  NAND2_X1  g331(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n469));
  AND3_X1   g333(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n470));
  AOI21_X1  g334(.A(new_n469), .B1(new_n470), .B2(new_n402), .ZN(new_n471));
  NAND2_X1  g335(.A1(new_n397), .A2(new_n401), .ZN(new_n472));
  NOR3_X1   g336(.A1(new_n436), .A2(new_n472), .A3(KEYINPUT26), .ZN(new_n473));
  NOR2_X1   g337(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g338(.A1(new_n468), .A2(new_n474), .A3(new_n397), .ZN(new_n475));
  NAND2_X1  g339(.A1(new_n332), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g340(.A1(new_n234), .A2(new_n313), .ZN(new_n477));
  INV_X1    g341(.A(new_n327), .ZN(new_n478));
  AOI21_X1  g342(.A(new_n478), .B1(new_n208), .B2(new_n228), .ZN(new_n479));
  OAI21_X1  g343(.A(new_n303), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g344(.A1(new_n480), .A2(new_n254), .ZN(new_n481));
  NAND2_X1  g345(.A1(new_n481), .A2(new_n258), .ZN(new_n482));
  INV_X1    g346(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g347(.A1(new_n476), .A2(new_n483), .ZN(G369));
  OR3_X1    g348(.A1(new_n225), .A2(KEYINPUT27), .A3(G20), .ZN(new_n485));
  OAI21_X1  g349(.A(KEYINPUT27), .B1(new_n225), .B2(G20), .ZN(new_n486));
  NAND3_X1  g350(.A1(new_n485), .A2(G213), .A3(new_n486), .ZN(new_n487));
  INV_X1    g351(.A(G343), .ZN(new_n488));
  NOR2_X1   g352(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g353(.A1(new_n353), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g354(.A1(new_n374), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g355(.A1(new_n490), .A2(new_n369), .ZN(new_n492));
  AND2_X1   g356(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g357(.A(new_n489), .ZN(new_n494));
  NAND2_X1  g358(.A1(new_n464), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g359(.A1(new_n494), .A2(new_n453), .ZN(new_n496));
  INV_X1    g360(.A(new_n496), .ZN(new_n497));
  OR2_X1    g361(.A1(new_n464), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g362(.A1(new_n461), .A2(new_n497), .ZN(new_n499));
  NAND2_X1  g363(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g364(.A(G330), .ZN(new_n501));
  NOR2_X1   g365(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g366(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g367(.A(new_n493), .B1(new_n495), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g368(.A1(new_n370), .A2(new_n489), .ZN(new_n505));
  OR2_X1    g369(.A1(new_n504), .A2(new_n505), .ZN(G399));
  INV_X1    g370(.A(new_n155), .ZN(new_n507));
  NOR2_X1   g371(.A1(new_n507), .A2(G41), .ZN(new_n508));
  INV_X1    g372(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g373(.A1(new_n380), .A2(G116), .ZN(new_n510));
  NAND3_X1  g374(.A1(new_n509), .A2(G1), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g375(.A(new_n511), .B1(new_n161), .B2(new_n509), .ZN(new_n512));
  XNOR2_X1  g376(.A(new_n512), .B(KEYINPUT28), .ZN(new_n513));
  INV_X1    g377(.A(new_n367), .ZN(new_n514));
  NAND4_X1  g378(.A1(new_n514), .A2(new_n410), .A3(new_n412), .A4(new_n396), .ZN(new_n515));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n516));
  NAND2_X1  g380(.A1(new_n455), .A2(G179), .ZN(new_n517));
  OR3_X1    g381(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g382(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n519));
  NOR3_X1   g383(.A1(new_n455), .A2(new_n396), .A3(G179), .ZN(new_n520));
  NAND3_X1  g384(.A1(new_n520), .A2(new_n367), .A3(new_n414), .ZN(new_n521));
  NAND3_X1  g385(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n523));
  NAND3_X1  g387(.A1(new_n522), .A2(new_n523), .A3(new_n489), .ZN(new_n524));
  INV_X1    g388(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g389(.A(new_n523), .B1(new_n462), .B2(new_n494), .ZN(new_n526));
  NAND2_X1  g390(.A1(new_n522), .A2(new_n489), .ZN(new_n527));
  AOI21_X1  g391(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g392(.A1(new_n528), .A2(G330), .ZN(new_n529));
  INV_X1    g393(.A(new_n397), .ZN(new_n530));
  AOI21_X1  g394(.A(new_n530), .B1(new_n466), .B2(new_n467), .ZN(new_n531));
  AOI21_X1  g395(.A(new_n489), .B1(new_n531), .B2(new_n474), .ZN(new_n532));
  AND2_X1   g396(.A1(new_n532), .A2(KEYINPUT29), .ZN(new_n533));
  NOR2_X1   g397(.A1(new_n532), .A2(KEYINPUT29), .ZN(new_n534));
  OAI21_X1  g398(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g399(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g400(.A(new_n513), .B1(new_n536), .B2(G1), .ZN(G364));
  AOI21_X1  g401(.A(new_n153), .B1(G20), .B2(new_n296), .ZN(new_n538));
  NOR2_X1   g402(.A1(new_n162), .A2(new_n252), .ZN(new_n539));
  INV_X1    g403(.A(new_n539), .ZN(new_n540));
  NOR3_X1   g404(.A1(new_n540), .A2(G179), .A3(G190), .ZN(new_n541));
  INV_X1    g405(.A(new_n541), .ZN(new_n542));
  INV_X1    g406(.A(G283), .ZN(new_n543));
  NOR2_X1   g407(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g408(.A1(new_n540), .A2(new_n306), .A3(G179), .ZN(new_n545));
  AOI21_X1  g409(.A(new_n181), .B1(new_n545), .B2(G303), .ZN(new_n546));
  NAND2_X1  g410(.A1(G20), .A2(G179), .ZN(new_n547));
  INV_X1    g411(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g412(.A1(new_n548), .A2(G200), .ZN(new_n549));
  NOR2_X1   g413(.A1(new_n549), .A2(G190), .ZN(new_n550));
  INV_X1    g414(.A(G317), .ZN(new_n551));
  OR2_X1    g415(.A1(new_n551), .A2(KEYINPUT33), .ZN(new_n552));
  NAND2_X1  g416(.A1(new_n551), .A2(KEYINPUT33), .ZN(new_n553));
  NAND3_X1  g417(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g418(.A(G294), .ZN(new_n555));
  NOR2_X1   g419(.A1(new_n539), .A2(new_n548), .ZN(new_n556));
  NAND2_X1  g420(.A1(new_n306), .A2(G20), .ZN(new_n557));
  NAND2_X1  g421(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g422(.A(new_n546), .B(new_n554), .C1(new_n555), .C2(new_n558), .ZN(new_n559));
  NOR3_X1   g423(.A1(new_n539), .A2(new_n548), .A3(new_n557), .ZN(new_n560));
  AOI211_X1 g424(.A(new_n544), .B(new_n559), .C1(G329), .C2(new_n560), .ZN(new_n561));
  INV_X1    g425(.A(G311), .ZN(new_n562));
  NOR3_X1   g426(.A1(new_n547), .A2(G190), .A3(G200), .ZN(new_n563));
  INV_X1    g427(.A(new_n563), .ZN(new_n564));
  INV_X1    g428(.A(G326), .ZN(new_n565));
  NOR2_X1   g429(.A1(new_n549), .A2(new_n306), .ZN(new_n566));
  INV_X1    g430(.A(new_n566), .ZN(new_n567));
  OAI221_X1 g431(.A(new_n561), .B1(new_n562), .B2(new_n564), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  NOR3_X1   g432(.A1(new_n547), .A2(new_n306), .A3(G200), .ZN(new_n569));
  AOI21_X1  g433(.A(new_n568), .B1(G322), .B2(new_n569), .ZN(new_n570));
  INV_X1    g434(.A(new_n550), .ZN(new_n571));
  OAI22_X1  g435(.A1(new_n542), .A2(new_n174), .B1(new_n571), .B2(new_n143), .ZN(new_n572));
  NAND2_X1  g436(.A1(new_n560), .A2(G159), .ZN(new_n573));
  XNOR2_X1  g437(.A(new_n573), .B(KEYINPUT32), .ZN(new_n574));
  AOI211_X1 g438(.A(new_n572), .B(new_n574), .C1(G87), .C2(new_n545), .ZN(new_n575));
  OAI21_X1  g439(.A(new_n575), .B1(new_n213), .B2(new_n567), .ZN(new_n576));
  INV_X1    g440(.A(new_n569), .ZN(new_n577));
  NOR2_X1   g441(.A1(new_n577), .A2(new_n269), .ZN(new_n578));
  OAI21_X1  g442(.A(new_n181), .B1(new_n564), .B2(new_n138), .ZN(new_n579));
  NOR2_X1   g443(.A1(new_n558), .A2(new_n378), .ZN(new_n580));
  NOR4_X1   g444(.A1(new_n576), .A2(new_n578), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  OAI21_X1  g445(.A(new_n538), .B1(new_n570), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g446(.A1(new_n507), .A2(new_n181), .ZN(new_n583));
  OR2_X1    g447(.A1(new_n161), .A2(G45), .ZN(new_n584));
  OAI211_X1 g448(.A(new_n583), .B(new_n584), .C1(new_n179), .C2(new_n192), .ZN(new_n585));
  INV_X1    g449(.A(G355), .ZN(new_n586));
  NAND2_X1  g450(.A1(new_n155), .A2(new_n181), .ZN(new_n587));
  OAI221_X1 g451(.A(new_n585), .B1(G116), .B2(new_n155), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NOR2_X1   g452(.A1(G13), .A2(G33), .ZN(new_n589));
  INV_X1    g453(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g454(.A1(new_n590), .A2(G20), .ZN(new_n591));
  NOR2_X1   g455(.A1(new_n591), .A2(new_n538), .ZN(new_n592));
  NAND2_X1  g456(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g457(.A1(new_n223), .A2(G20), .ZN(new_n594));
  NAND2_X1  g458(.A1(new_n594), .A2(G45), .ZN(new_n595));
  NAND3_X1  g459(.A1(new_n509), .A2(G1), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g460(.A(new_n596), .B1(new_n500), .B2(new_n591), .ZN(new_n597));
  NAND3_X1  g461(.A1(new_n582), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g462(.A(new_n500), .B(new_n501), .ZN(new_n599));
  INV_X1    g463(.A(new_n596), .ZN(new_n600));
  OAI21_X1  g464(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(G396));
  OAI211_X1 g465(.A(new_n327), .B(new_n330), .C1(new_n329), .C2(new_n494), .ZN(new_n602));
  OAI211_X1 g466(.A(new_n319), .B(new_n489), .C1(new_n325), .C2(new_n326), .ZN(new_n603));
  NAND2_X1  g467(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g468(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g469(.A1(new_n529), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g470(.A1(new_n374), .A2(new_n437), .ZN(new_n607));
  INV_X1    g471(.A(new_n461), .ZN(new_n608));
  NAND3_X1  g472(.A1(new_n607), .A2(new_n608), .A3(new_n494), .ZN(new_n609));
  NAND3_X1  g473(.A1(new_n609), .A2(KEYINPUT31), .A3(new_n527), .ZN(new_n610));
  NAND4_X1  g474(.A1(new_n610), .A2(G330), .A3(new_n524), .A4(new_n604), .ZN(new_n611));
  NAND2_X1  g475(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g476(.A(new_n612), .B(new_n532), .ZN(new_n613));
  NAND2_X1  g477(.A1(new_n605), .A2(new_n589), .ZN(new_n614));
  INV_X1    g478(.A(new_n538), .ZN(new_n615));
  OAI221_X1 g479(.A(new_n264), .B1(new_n378), .B2(new_n558), .C1(new_n542), .C2(new_n291), .ZN(new_n616));
  NOR2_X1   g480(.A1(new_n564), .A2(new_n389), .ZN(new_n617));
  OAI22_X1  g481(.A1(new_n571), .A2(new_n543), .B1(new_n567), .B2(new_n440), .ZN(new_n618));
  INV_X1    g482(.A(new_n545), .ZN(new_n619));
  NOR2_X1   g483(.A1(new_n619), .A2(new_n174), .ZN(new_n620));
  NOR4_X1   g484(.A1(new_n616), .A2(new_n617), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  INV_X1    g485(.A(new_n560), .ZN(new_n622));
  OAI221_X1 g486(.A(new_n621), .B1(new_n555), .B2(new_n577), .C1(new_n562), .C2(new_n622), .ZN(new_n623));
  AOI22_X1  g487(.A1(G143), .A2(new_n569), .B1(new_n563), .B2(G159), .ZN(new_n624));
  INV_X1    g488(.A(G137), .ZN(new_n625));
  INV_X1    g489(.A(G150), .ZN(new_n626));
  OAI221_X1 g490(.A(new_n624), .B1(new_n567), .B2(new_n625), .C1(new_n626), .C2(new_n571), .ZN(new_n627));
  XNOR2_X1  g491(.A(new_n627), .B(KEYINPUT34), .ZN(new_n628));
  AOI22_X1  g492(.A1(G50), .A2(new_n545), .B1(new_n541), .B2(G68), .ZN(new_n629));
  INV_X1    g493(.A(G132), .ZN(new_n630));
  OAI211_X1 g494(.A(new_n629), .B(new_n181), .C1(new_n630), .C2(new_n622), .ZN(new_n631));
  INV_X1    g495(.A(new_n558), .ZN(new_n632));
  AOI21_X1  g496(.A(new_n631), .B1(G58), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g497(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g498(.A(new_n615), .B1(new_n623), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g499(.A1(new_n538), .A2(new_n589), .ZN(new_n636));
  AOI211_X1 g500(.A(new_n596), .B(new_n635), .C1(new_n138), .C2(new_n636), .ZN(new_n637));
  AOI22_X1  g501(.A1(new_n613), .A2(new_n596), .B1(new_n614), .B2(new_n637), .ZN(new_n638));
  INV_X1    g502(.A(new_n638), .ZN(G384));
  NAND2_X1  g503(.A1(new_n303), .A2(new_n313), .ZN(new_n640));
  INV_X1    g504(.A(new_n487), .ZN(new_n641));
  NAND2_X1  g505(.A1(new_n288), .A2(new_n641), .ZN(new_n642));
  INV_X1    g506(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g507(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g508(.A(KEYINPUT37), .ZN(new_n645));
  OAI22_X1  g509(.A1(new_n304), .A2(new_n487), .B1(new_n311), .B2(new_n307), .ZN(new_n646));
  AND3_X1   g510(.A1(new_n288), .A2(new_n297), .A3(new_n298), .ZN(new_n647));
  OAI21_X1  g511(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g512(.A1(new_n304), .A2(new_n308), .A3(new_n309), .ZN(new_n649));
  NAND4_X1  g513(.A1(new_n649), .A2(KEYINPUT37), .A3(new_n299), .A4(new_n642), .ZN(new_n650));
  AND2_X1   g514(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g515(.A1(new_n644), .A2(new_n651), .A3(KEYINPUT38), .ZN(new_n652));
  INV_X1    g516(.A(KEYINPUT38), .ZN(new_n653));
  AOI21_X1  g517(.A(new_n642), .B1(new_n303), .B2(new_n313), .ZN(new_n654));
  NAND2_X1  g518(.A1(new_n648), .A2(new_n650), .ZN(new_n655));
  OAI21_X1  g519(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g520(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g521(.A1(new_n228), .A2(new_n489), .ZN(new_n658));
  NAND3_X1  g522(.A1(new_n229), .A2(new_n234), .A3(new_n658), .ZN(new_n659));
  OAI211_X1 g523(.A(new_n228), .B(new_n489), .C1(new_n233), .C2(new_n208), .ZN(new_n660));
  AND2_X1   g524(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g525(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g526(.A1(new_n657), .A2(new_n528), .A3(new_n662), .A4(new_n604), .ZN(new_n663));
  INV_X1    g527(.A(KEYINPUT40), .ZN(new_n664));
  NAND2_X1  g528(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g529(.A(new_n661), .B1(new_n656), .B2(new_n652), .ZN(new_n666));
  NAND4_X1  g530(.A1(new_n666), .A2(KEYINPUT40), .A3(new_n528), .A4(new_n604), .ZN(new_n667));
  NAND2_X1  g531(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g532(.A1(new_n332), .A2(new_n528), .ZN(new_n669));
  XOR2_X1   g533(.A(new_n668), .B(new_n669), .Z(new_n670));
  NAND2_X1  g534(.A1(new_n670), .A2(G330), .ZN(new_n671));
  NOR2_X1   g535(.A1(new_n303), .A2(new_n641), .ZN(new_n672));
  INV_X1    g536(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g537(.A1(new_n657), .A2(new_n662), .ZN(new_n674));
  AOI21_X1  g538(.A(new_n605), .B1(new_n531), .B2(new_n474), .ZN(new_n675));
  OAI21_X1  g539(.A(new_n494), .B1(new_n675), .B2(new_n478), .ZN(new_n676));
  OAI21_X1  g540(.A(new_n673), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g541(.A1(new_n229), .A2(new_n489), .ZN(new_n678));
  INV_X1    g542(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g543(.A(KEYINPUT38), .B1(new_n644), .B2(new_n651), .ZN(new_n680));
  NOR3_X1   g544(.A1(new_n654), .A2(new_n655), .A3(new_n653), .ZN(new_n681));
  OAI21_X1  g545(.A(KEYINPUT39), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g546(.A(KEYINPUT39), .ZN(new_n683));
  NAND3_X1  g547(.A1(new_n652), .A2(new_n683), .A3(new_n656), .ZN(new_n684));
  AOI21_X1  g548(.A(new_n679), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g549(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g550(.A1(new_n533), .A2(new_n534), .ZN(new_n687));
  INV_X1    g551(.A(new_n332), .ZN(new_n688));
  OAI21_X1  g552(.A(new_n483), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g553(.A(new_n686), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g554(.A(new_n671), .B(new_n690), .ZN(new_n691));
  OAI21_X1  g555(.A(new_n691), .B1(new_n346), .B2(new_n594), .ZN(new_n692));
  AOI211_X1 g556(.A(new_n162), .B(new_n153), .C1(new_n425), .C2(KEYINPUT35), .ZN(new_n693));
  OAI211_X1 g557(.A(new_n693), .B(G116), .C1(KEYINPUT35), .C2(new_n425), .ZN(new_n694));
  XNOR2_X1  g558(.A(new_n694), .B(KEYINPUT36), .ZN(new_n695));
  OAI21_X1  g559(.A(G77), .B1(new_n269), .B2(new_n143), .ZN(new_n696));
  OAI22_X1  g560(.A1(new_n696), .A2(new_n161), .B1(G50), .B2(new_n143), .ZN(new_n697));
  NAND3_X1  g561(.A1(new_n697), .A2(G1), .A3(new_n223), .ZN(new_n698));
  NAND3_X1  g562(.A1(new_n692), .A2(new_n695), .A3(new_n698), .ZN(G367));
  XOR2_X1   g563(.A(new_n508), .B(KEYINPUT41), .Z(new_n700));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n701));
  NOR2_X1   g565(.A1(new_n493), .A2(new_n495), .ZN(new_n702));
  NOR2_X1   g566(.A1(new_n702), .A2(new_n505), .ZN(new_n703));
  NAND2_X1  g567(.A1(new_n433), .A2(new_n489), .ZN(new_n704));
  NAND2_X1  g568(.A1(new_n430), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g569(.A1(new_n705), .A2(new_n436), .ZN(new_n706));
  OAI21_X1  g570(.A(new_n706), .B1(new_n436), .B2(new_n489), .ZN(new_n707));
  INV_X1    g571(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g572(.A(new_n701), .B1(new_n703), .B2(new_n708), .ZN(new_n709));
  NOR4_X1   g573(.A1(new_n702), .A2(KEYINPUT45), .A3(new_n505), .A4(new_n707), .ZN(new_n710));
  NOR2_X1   g574(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n712));
  OAI21_X1  g576(.A(new_n712), .B1(new_n703), .B2(new_n708), .ZN(new_n713));
  OAI211_X1 g577(.A(KEYINPUT44), .B(new_n707), .C1(new_n702), .C2(new_n505), .ZN(new_n714));
  NAND2_X1  g578(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g579(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g580(.A1(new_n491), .A2(new_n492), .ZN(new_n717));
  AOI211_X1 g581(.A(new_n502), .B(new_n717), .C1(new_n464), .C2(new_n494), .ZN(new_n718));
  NOR2_X1   g582(.A1(new_n718), .A2(new_n504), .ZN(new_n719));
  NAND2_X1  g583(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g584(.A(new_n700), .B1(new_n720), .B2(new_n536), .ZN(new_n721));
  OR2_X1    g585(.A1(new_n494), .A2(new_n399), .ZN(new_n722));
  NOR2_X1   g586(.A1(new_n530), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g587(.A(new_n723), .B1(new_n472), .B2(new_n722), .ZN(new_n724));
  INV_X1    g588(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g589(.A(KEYINPUT42), .B1(new_n370), .B2(new_n489), .ZN(new_n726));
  OAI211_X1 g590(.A(new_n708), .B(new_n726), .C1(new_n702), .C2(new_n505), .ZN(new_n727));
  NAND4_X1  g591(.A1(new_n717), .A2(new_n464), .A3(new_n494), .A4(new_n706), .ZN(new_n728));
  AOI22_X1  g592(.A1(new_n728), .A2(KEYINPUT42), .B1(new_n470), .B2(new_n494), .ZN(new_n729));
  NAND2_X1  g593(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n731));
  OAI21_X1  g595(.A(new_n725), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g596(.A(KEYINPUT43), .B1(new_n727), .B2(new_n729), .ZN(new_n733));
  NOR2_X1   g597(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g598(.A(new_n730), .ZN(new_n735));
  NOR3_X1   g599(.A1(new_n735), .A2(KEYINPUT43), .A3(new_n725), .ZN(new_n736));
  NOR2_X1   g600(.A1(new_n493), .A2(new_n503), .ZN(new_n737));
  INV_X1    g601(.A(new_n737), .ZN(new_n738));
  OAI22_X1  g602(.A1(new_n734), .A2(new_n736), .B1(new_n738), .B2(new_n707), .ZN(new_n739));
  NAND2_X1  g603(.A1(new_n735), .A2(KEYINPUT43), .ZN(new_n740));
  INV_X1    g604(.A(new_n733), .ZN(new_n741));
  NAND3_X1  g605(.A1(new_n740), .A2(new_n725), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g606(.A1(new_n738), .A2(new_n707), .ZN(new_n743));
  NAND2_X1  g607(.A1(new_n732), .A2(new_n733), .ZN(new_n744));
  NAND3_X1  g608(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g609(.A1(new_n721), .A2(new_n739), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g610(.A1(new_n595), .A2(G1), .ZN(new_n747));
  NAND3_X1  g611(.A1(new_n739), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g612(.A(new_n583), .ZN(new_n749));
  OAI221_X1 g613(.A(new_n592), .B1(new_n155), .B2(new_n315), .C1(new_n167), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g614(.A(new_n596), .B1(new_n725), .B2(new_n591), .ZN(new_n751));
  NAND2_X1  g615(.A1(new_n560), .A2(G137), .ZN(new_n752));
  AOI21_X1  g616(.A(new_n264), .B1(G150), .B2(new_n569), .ZN(new_n753));
  OAI221_X1 g617(.A(new_n753), .B1(new_n143), .B2(new_n558), .C1(new_n619), .C2(new_n269), .ZN(new_n754));
  NOR2_X1   g618(.A1(new_n542), .A2(new_n138), .ZN(new_n755));
  AOI21_X1  g619(.A(new_n755), .B1(G143), .B2(new_n566), .ZN(new_n756));
  INV_X1    g620(.A(G159), .ZN(new_n757));
  OAI21_X1  g621(.A(new_n756), .B1(new_n757), .B2(new_n571), .ZN(new_n758));
  AOI211_X1 g622(.A(new_n754), .B(new_n758), .C1(G50), .C2(new_n563), .ZN(new_n759));
  NOR2_X1   g623(.A1(new_n558), .A2(new_n174), .ZN(new_n760));
  NAND2_X1  g624(.A1(new_n545), .A2(G116), .ZN(new_n761));
  XNOR2_X1  g625(.A(new_n761), .B(KEYINPUT46), .ZN(new_n762));
  NAND2_X1  g626(.A1(new_n563), .A2(G283), .ZN(new_n763));
  AOI22_X1  g627(.A1(new_n541), .A2(G97), .B1(new_n550), .B2(G294), .ZN(new_n764));
  AOI21_X1  g628(.A(new_n181), .B1(G303), .B2(new_n569), .ZN(new_n765));
  NAND4_X1  g629(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  AOI211_X1 g630(.A(new_n760), .B(new_n766), .C1(G311), .C2(new_n566), .ZN(new_n767));
  NAND2_X1  g631(.A1(new_n560), .A2(G317), .ZN(new_n768));
  AOI22_X1  g632(.A1(new_n752), .A2(new_n759), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g633(.A(new_n769), .B(KEYINPUT47), .ZN(new_n770));
  OAI211_X1 g634(.A(new_n750), .B(new_n751), .C1(new_n770), .C2(new_n615), .ZN(new_n771));
  NAND3_X1  g635(.A1(new_n746), .A2(new_n748), .A3(new_n771), .ZN(G387));
  NOR2_X1   g636(.A1(new_n558), .A2(new_n315), .ZN(new_n773));
  AOI21_X1  g637(.A(new_n773), .B1(G159), .B2(new_n566), .ZN(new_n774));
  OAI21_X1  g638(.A(new_n774), .B1(new_n626), .B2(new_n622), .ZN(new_n775));
  AOI21_X1  g639(.A(new_n775), .B1(G68), .B2(new_n563), .ZN(new_n776));
  NAND2_X1  g640(.A1(new_n545), .A2(G77), .ZN(new_n777));
  AOI22_X1  g641(.A1(new_n541), .A2(G97), .B1(G50), .B2(new_n569), .ZN(new_n778));
  AOI21_X1  g642(.A(new_n264), .B1(new_n550), .B2(new_n285), .ZN(new_n779));
  NAND4_X1  g643(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  AOI22_X1  g644(.A1(new_n550), .A2(G311), .B1(G317), .B2(new_n569), .ZN(new_n781));
  INV_X1    g645(.A(G322), .ZN(new_n782));
  OAI221_X1 g646(.A(new_n781), .B1(new_n440), .B2(new_n564), .C1(new_n782), .C2(new_n567), .ZN(new_n783));
  XNOR2_X1  g647(.A(new_n783), .B(KEYINPUT48), .ZN(new_n784));
  OAI221_X1 g648(.A(new_n784), .B1(new_n543), .B2(new_n558), .C1(new_n555), .C2(new_n619), .ZN(new_n785));
  XOR2_X1   g649(.A(new_n785), .B(KEYINPUT49), .Z(new_n786));
  OAI221_X1 g650(.A(new_n264), .B1(new_n622), .B2(new_n565), .C1(new_n542), .C2(new_n389), .ZN(new_n787));
  OAI21_X1  g651(.A(new_n780), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g652(.A(new_n596), .B1(new_n788), .B2(new_n538), .ZN(new_n789));
  INV_X1    g653(.A(new_n591), .ZN(new_n790));
  OAI21_X1  g654(.A(new_n789), .B1(new_n717), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g655(.A1(new_n246), .A2(KEYINPUT50), .A3(G50), .ZN(new_n792));
  NOR3_X1   g656(.A1(new_n792), .A2(G116), .A3(new_n380), .ZN(new_n793));
  NAND2_X1  g657(.A1(G68), .A2(G77), .ZN(new_n794));
  OAI21_X1  g658(.A(KEYINPUT50), .B1(new_n246), .B2(G50), .ZN(new_n795));
  NAND4_X1  g659(.A1(new_n793), .A2(new_n192), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  OAI211_X1 g660(.A(new_n583), .B(new_n796), .C1(new_n171), .C2(new_n192), .ZN(new_n797));
  OAI221_X1 g661(.A(new_n797), .B1(G107), .B2(new_n155), .C1(new_n510), .C2(new_n587), .ZN(new_n798));
  AOI21_X1  g662(.A(new_n791), .B1(new_n592), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g663(.A(new_n799), .B1(new_n747), .B2(new_n719), .ZN(new_n800));
  NAND2_X1  g664(.A1(new_n536), .A2(new_n719), .ZN(new_n801));
  NAND2_X1  g665(.A1(new_n801), .A2(new_n508), .ZN(new_n802));
  NOR2_X1   g666(.A1(new_n536), .A2(new_n719), .ZN(new_n803));
  OAI21_X1  g667(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(G393));
  NAND2_X1  g668(.A1(new_n716), .A2(new_n737), .ZN(new_n805));
  NAND3_X1  g669(.A1(new_n711), .A2(new_n738), .A3(new_n715), .ZN(new_n806));
  NAND4_X1  g670(.A1(new_n805), .A2(new_n536), .A3(new_n719), .A4(new_n806), .ZN(new_n807));
  AND3_X1   g671(.A1(new_n711), .A2(new_n738), .A3(new_n715), .ZN(new_n808));
  AOI21_X1  g672(.A(new_n738), .B1(new_n711), .B2(new_n715), .ZN(new_n809));
  OAI21_X1  g673(.A(new_n801), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g674(.A1(new_n807), .A2(new_n810), .A3(new_n508), .ZN(new_n811));
  OAI22_X1  g675(.A1(new_n567), .A2(new_n551), .B1(new_n562), .B2(new_n577), .ZN(new_n812));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n813));
  OAI221_X1 g677(.A(new_n264), .B1(new_n174), .B2(new_n542), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AND2_X1   g678(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NOR2_X1   g679(.A1(new_n571), .A2(new_n440), .ZN(new_n816));
  OAI22_X1  g680(.A1(new_n622), .A2(new_n782), .B1(new_n555), .B2(new_n564), .ZN(new_n817));
  NOR4_X1   g681(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  OAI221_X1 g682(.A(new_n818), .B1(new_n389), .B2(new_n558), .C1(new_n543), .C2(new_n619), .ZN(new_n819));
  NOR2_X1   g683(.A1(new_n558), .A2(new_n138), .ZN(new_n820));
  AOI22_X1  g684(.A1(new_n566), .A2(G150), .B1(G159), .B2(new_n569), .ZN(new_n821));
  XNOR2_X1  g685(.A(new_n821), .B(KEYINPUT51), .ZN(new_n822));
  OAI22_X1  g686(.A1(new_n542), .A2(new_n291), .B1(new_n619), .B2(new_n143), .ZN(new_n823));
  NOR3_X1   g687(.A1(new_n822), .A2(new_n264), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g688(.A1(new_n285), .A2(new_n563), .ZN(new_n825));
  NAND2_X1  g689(.A1(new_n560), .A2(G143), .ZN(new_n826));
  NAND2_X1  g690(.A1(new_n550), .A2(G50), .ZN(new_n827));
  NAND4_X1  g691(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g692(.A(new_n819), .B1(new_n820), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g693(.A1(new_n829), .A2(new_n538), .ZN(new_n830));
  OAI221_X1 g694(.A(new_n592), .B1(new_n378), .B2(new_n155), .C1(new_n176), .C2(new_n749), .ZN(new_n831));
  NAND2_X1  g695(.A1(new_n707), .A2(new_n591), .ZN(new_n832));
  AND4_X1   g696(.A1(new_n600), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g697(.A1(new_n808), .A2(new_n809), .ZN(new_n834));
  AOI21_X1  g698(.A(new_n833), .B1(new_n834), .B2(new_n747), .ZN(new_n835));
  NAND2_X1  g699(.A1(new_n811), .A2(new_n835), .ZN(G390));
  OAI211_X1 g700(.A(new_n679), .B(new_n657), .C1(new_n676), .C2(new_n235), .ZN(new_n837));
  NAND2_X1  g701(.A1(new_n475), .A2(new_n604), .ZN(new_n838));
  AOI21_X1  g702(.A(new_n489), .B1(new_n838), .B2(new_n327), .ZN(new_n839));
  AOI21_X1  g703(.A(new_n678), .B1(new_n839), .B2(new_n236), .ZN(new_n840));
  NAND2_X1  g704(.A1(new_n682), .A2(new_n684), .ZN(new_n841));
  OAI21_X1  g705(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g706(.A1(new_n611), .A2(new_n661), .ZN(new_n843));
  AND2_X1   g707(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g708(.A1(new_n611), .A2(new_n661), .ZN(new_n845));
  OAI211_X1 g709(.A(new_n837), .B(new_n845), .C1(new_n840), .C2(new_n841), .ZN(new_n846));
  INV_X1    g710(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g711(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g712(.A(new_n482), .B1(new_n535), .B2(new_n332), .ZN(new_n849));
  NAND2_X1  g713(.A1(new_n611), .A2(new_n661), .ZN(new_n850));
  INV_X1    g714(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g715(.A(new_n839), .B1(new_n851), .B2(new_n843), .ZN(new_n852));
  NAND3_X1  g716(.A1(new_n845), .A2(new_n676), .A3(new_n850), .ZN(new_n853));
  NAND2_X1  g717(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g718(.A1(new_n848), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g719(.A1(new_n854), .A2(new_n849), .ZN(new_n856));
  OAI21_X1  g720(.A(new_n856), .B1(new_n844), .B2(new_n847), .ZN(new_n857));
  NAND3_X1  g721(.A1(new_n855), .A2(new_n508), .A3(new_n857), .ZN(new_n858));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n859));
  OAI21_X1  g723(.A(new_n859), .B1(new_n619), .B2(new_n626), .ZN(new_n860));
  NAND3_X1  g724(.A1(new_n545), .A2(KEYINPUT53), .A3(G150), .ZN(new_n861));
  AOI21_X1  g725(.A(new_n264), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g726(.A1(new_n541), .A2(G50), .ZN(new_n863));
  NAND2_X1  g727(.A1(new_n566), .A2(G128), .ZN(new_n864));
  AOI22_X1  g728(.A1(new_n632), .A2(G159), .B1(G132), .B2(new_n569), .ZN(new_n865));
  NAND4_X1  g729(.A1(new_n862), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  XNOR2_X1  g730(.A(KEYINPUT54), .B(G143), .ZN(new_n867));
  NOR2_X1   g731(.A1(new_n564), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g732(.A1(new_n571), .A2(new_n625), .ZN(new_n869));
  INV_X1    g733(.A(G125), .ZN(new_n870));
  NOR2_X1   g734(.A1(new_n622), .A2(new_n870), .ZN(new_n871));
  NOR4_X1   g735(.A1(new_n866), .A2(new_n868), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g736(.A1(new_n622), .A2(new_n555), .ZN(new_n873));
  AOI21_X1  g737(.A(new_n820), .B1(G68), .B2(new_n541), .ZN(new_n874));
  NAND2_X1  g738(.A1(new_n566), .A2(G283), .ZN(new_n875));
  AOI22_X1  g739(.A1(new_n545), .A2(G87), .B1(new_n550), .B2(G107), .ZN(new_n876));
  AOI21_X1  g740(.A(new_n181), .B1(G97), .B2(new_n563), .ZN(new_n877));
  NAND4_X1  g741(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI211_X1 g742(.A(new_n873), .B(new_n878), .C1(G116), .C2(new_n569), .ZN(new_n879));
  OAI21_X1  g743(.A(new_n538), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g744(.A(new_n880), .B1(new_n841), .B2(new_n590), .ZN(new_n881));
  AOI21_X1  g745(.A(new_n881), .B1(new_n246), .B2(new_n636), .ZN(new_n882));
  AOI22_X1  g746(.A1(new_n848), .A2(new_n747), .B1(new_n600), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g747(.A1(new_n858), .A2(new_n883), .ZN(G378));
  NAND2_X1  g748(.A1(new_n842), .A2(new_n843), .ZN(new_n885));
  NAND3_X1  g749(.A1(new_n885), .A2(new_n854), .A3(new_n846), .ZN(new_n886));
  NAND2_X1  g750(.A1(new_n886), .A2(new_n849), .ZN(new_n887));
  NAND3_X1  g751(.A1(new_n665), .A2(G330), .A3(new_n667), .ZN(new_n888));
  NAND2_X1  g752(.A1(new_n888), .A2(new_n686), .ZN(new_n889));
  AND3_X1   g753(.A1(new_n652), .A2(new_n683), .A3(new_n656), .ZN(new_n890));
  AOI21_X1  g754(.A(new_n683), .B1(new_n652), .B2(new_n656), .ZN(new_n891));
  OAI21_X1  g755(.A(new_n678), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g756(.A(new_n672), .B1(new_n666), .B2(new_n839), .ZN(new_n893));
  NAND2_X1  g757(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g758(.A1(new_n894), .A2(G330), .A3(new_n665), .A4(new_n667), .ZN(new_n895));
  NAND2_X1  g759(.A1(new_n254), .A2(new_n258), .ZN(new_n896));
  NAND2_X1  g760(.A1(new_n250), .A2(new_n641), .ZN(new_n897));
  XNOR2_X1  g761(.A(new_n896), .B(new_n897), .ZN(new_n898));
  XOR2_X1   g762(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n899));
  XNOR2_X1  g763(.A(new_n898), .B(new_n899), .ZN(new_n900));
  AND3_X1   g764(.A1(new_n889), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g765(.A(new_n900), .B1(new_n889), .B2(new_n895), .ZN(new_n902));
  OAI21_X1  g766(.A(new_n887), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g767(.A(KEYINPUT57), .ZN(new_n904));
  NAND2_X1  g768(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g769(.A(new_n887), .B(KEYINPUT57), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  NAND3_X1  g770(.A1(new_n905), .A2(new_n508), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g771(.A(new_n747), .B1(new_n901), .B2(new_n902), .ZN(new_n908));
  AOI21_X1  g772(.A(new_n596), .B1(new_n900), .B2(new_n589), .ZN(new_n909));
  NAND2_X1  g773(.A1(new_n264), .A2(new_n191), .ZN(new_n910));
  OAI211_X1 g774(.A(new_n910), .B(new_n213), .C1(G33), .C2(G41), .ZN(new_n911));
  AOI22_X1  g775(.A1(new_n632), .A2(G150), .B1(G132), .B2(new_n550), .ZN(new_n912));
  INV_X1    g776(.A(G128), .ZN(new_n913));
  OAI21_X1  g777(.A(new_n912), .B1(new_n913), .B2(new_n577), .ZN(new_n914));
  INV_X1    g778(.A(new_n867), .ZN(new_n915));
  AOI21_X1  g779(.A(new_n914), .B1(new_n545), .B2(new_n915), .ZN(new_n916));
  OAI221_X1 g780(.A(new_n916), .B1(new_n870), .B2(new_n567), .C1(new_n625), .C2(new_n564), .ZN(new_n917));
  XOR2_X1   g781(.A(new_n917), .B(KEYINPUT59), .Z(new_n918));
  NAND2_X1  g782(.A1(new_n560), .A2(G124), .ZN(new_n919));
  NAND4_X1  g783(.A1(new_n918), .A2(new_n260), .A3(new_n191), .A4(new_n919), .ZN(new_n920));
  NOR2_X1   g784(.A1(new_n542), .A2(new_n757), .ZN(new_n921));
  OAI21_X1  g785(.A(new_n911), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g786(.A1(new_n542), .A2(new_n269), .ZN(new_n923));
  OAI221_X1 g787(.A(new_n777), .B1(new_n564), .B2(new_n315), .C1(new_n378), .C2(new_n571), .ZN(new_n924));
  AOI211_X1 g788(.A(new_n923), .B(new_n924), .C1(G283), .C2(new_n560), .ZN(new_n925));
  NOR2_X1   g789(.A1(new_n558), .A2(new_n143), .ZN(new_n926));
  AOI211_X1 g790(.A(new_n910), .B(new_n926), .C1(G116), .C2(new_n566), .ZN(new_n927));
  OAI211_X1 g791(.A(new_n925), .B(new_n927), .C1(new_n174), .C2(new_n577), .ZN(new_n928));
  XOR2_X1   g792(.A(new_n928), .B(KEYINPUT58), .Z(new_n929));
  OAI21_X1  g793(.A(new_n538), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g794(.A1(new_n636), .A2(new_n213), .ZN(new_n931));
  NAND3_X1  g795(.A1(new_n909), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g796(.A1(new_n908), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g797(.A1(new_n907), .A2(new_n933), .ZN(G375));
  NAND2_X1  g798(.A1(new_n661), .A2(new_n589), .ZN(new_n935));
  OAI221_X1 g799(.A(new_n181), .B1(new_n558), .B2(new_n213), .C1(new_n913), .C2(new_n622), .ZN(new_n936));
  OAI22_X1  g800(.A1(new_n542), .A2(new_n269), .B1(new_n567), .B2(new_n630), .ZN(new_n937));
  NOR2_X1   g801(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g802(.A(new_n938), .B1(new_n625), .B2(new_n577), .ZN(new_n939));
  AOI21_X1  g803(.A(new_n939), .B1(new_n550), .B2(new_n915), .ZN(new_n940));
  OAI221_X1 g804(.A(new_n940), .B1(new_n626), .B2(new_n564), .C1(new_n757), .C2(new_n619), .ZN(new_n941));
  OAI22_X1  g805(.A1(new_n571), .A2(new_n389), .B1(new_n543), .B2(new_n577), .ZN(new_n942));
  OAI21_X1  g806(.A(new_n264), .B1(new_n564), .B2(new_n174), .ZN(new_n943));
  OR4_X1    g807(.A1(new_n755), .A2(new_n942), .A3(new_n773), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g808(.A(new_n944), .B1(G294), .B2(new_n566), .ZN(new_n945));
  OAI221_X1 g809(.A(new_n945), .B1(new_n378), .B2(new_n619), .C1(new_n440), .C2(new_n622), .ZN(new_n946));
  AOI21_X1  g810(.A(new_n615), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  AOI211_X1 g811(.A(new_n596), .B(new_n947), .C1(new_n143), .C2(new_n636), .ZN(new_n948));
  AOI22_X1  g812(.A1(new_n854), .A2(new_n747), .B1(new_n935), .B2(new_n948), .ZN(new_n949));
  INV_X1    g813(.A(new_n700), .ZN(new_n950));
  NAND2_X1  g814(.A1(new_n856), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g815(.A1(new_n854), .A2(new_n849), .ZN(new_n952));
  OAI21_X1  g816(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G381));
  NOR4_X1   g817(.A1(G375), .A2(G396), .A3(G393), .A4(G378), .ZN(new_n954));
  OR2_X1    g818(.A1(G387), .A2(G390), .ZN(new_n955));
  NOR3_X1   g819(.A1(new_n955), .A2(G384), .A3(G381), .ZN(new_n956));
  NAND2_X1  g820(.A1(new_n954), .A2(new_n956), .ZN(G407));
  AND2_X1   g821(.A1(new_n858), .A2(new_n883), .ZN(new_n958));
  NAND4_X1  g822(.A1(new_n907), .A2(new_n958), .A3(new_n488), .A4(new_n933), .ZN(new_n959));
  NAND3_X1  g823(.A1(G407), .A2(G213), .A3(new_n959), .ZN(G409));
  INV_X1    g824(.A(KEYINPUT60), .ZN(new_n961));
  OAI21_X1  g825(.A(new_n961), .B1(new_n854), .B2(new_n849), .ZN(new_n962));
  INV_X1    g826(.A(new_n849), .ZN(new_n963));
  NAND4_X1  g827(.A1(new_n963), .A2(KEYINPUT60), .A3(new_n852), .A4(new_n853), .ZN(new_n964));
  NAND4_X1  g828(.A1(new_n962), .A2(new_n964), .A3(new_n508), .A4(new_n856), .ZN(new_n965));
  NAND3_X1  g829(.A1(new_n965), .A2(new_n638), .A3(new_n949), .ZN(new_n966));
  INV_X1    g830(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g831(.A(new_n638), .B1(new_n965), .B2(new_n949), .ZN(new_n968));
  NOR2_X1   g832(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g833(.A1(new_n488), .A2(G213), .ZN(new_n970));
  INV_X1    g834(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g835(.A1(new_n907), .A2(G378), .A3(new_n933), .ZN(new_n972));
  OAI211_X1 g836(.A(new_n908), .B(new_n932), .C1(new_n903), .C2(new_n700), .ZN(new_n973));
  NAND2_X1  g837(.A1(new_n958), .A2(new_n973), .ZN(new_n974));
  AOI211_X1 g838(.A(new_n969), .B(new_n971), .C1(new_n972), .C2(new_n974), .ZN(new_n975));
  INV_X1    g839(.A(KEYINPUT62), .ZN(new_n976));
  AOI21_X1  g840(.A(KEYINPUT61), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g841(.A1(new_n971), .A2(G2897), .ZN(new_n978));
  OR2_X1    g842(.A1(new_n969), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g843(.A1(new_n972), .A2(new_n974), .ZN(new_n980));
  NAND2_X1  g844(.A1(new_n980), .A2(new_n970), .ZN(new_n981));
  OAI21_X1  g845(.A(KEYINPUT62), .B1(new_n981), .B2(new_n969), .ZN(new_n982));
  NAND3_X1  g846(.A1(new_n981), .A2(new_n969), .A3(new_n978), .ZN(new_n983));
  NAND4_X1  g847(.A1(new_n977), .A2(new_n979), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g848(.A1(G387), .A2(G390), .ZN(new_n985));
  INV_X1    g849(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g850(.A1(G387), .A2(G390), .ZN(new_n987));
  XOR2_X1   g851(.A(G393), .B(G396), .Z(new_n988));
  NOR3_X1   g852(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  XNOR2_X1  g853(.A(G393), .B(G396), .ZN(new_n990));
  AOI21_X1  g854(.A(new_n990), .B1(new_n955), .B2(new_n985), .ZN(new_n991));
  NOR2_X1   g855(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g856(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g857(.A1(new_n984), .A2(new_n993), .ZN(new_n994));
  INV_X1    g858(.A(new_n969), .ZN(new_n995));
  NAND4_X1  g859(.A1(new_n980), .A2(KEYINPUT63), .A3(new_n995), .A4(new_n970), .ZN(new_n996));
  NAND2_X1  g860(.A1(new_n996), .A2(new_n992), .ZN(new_n997));
  AOI21_X1  g861(.A(new_n971), .B1(new_n972), .B2(new_n974), .ZN(new_n998));
  AOI21_X1  g862(.A(KEYINPUT63), .B1(new_n998), .B2(new_n995), .ZN(new_n999));
  NOR2_X1   g863(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g864(.A(KEYINPUT61), .ZN(new_n1001));
  NAND4_X1  g865(.A1(new_n1000), .A2(new_n1001), .A3(new_n979), .A4(new_n983), .ZN(new_n1002));
  NAND2_X1  g866(.A1(new_n994), .A2(new_n1002), .ZN(G405));
  NAND2_X1  g867(.A1(G375), .A2(new_n958), .ZN(new_n1004));
  NAND2_X1  g868(.A1(new_n1004), .A2(new_n972), .ZN(new_n1005));
  OR2_X1    g869(.A1(new_n992), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g870(.A1(new_n992), .A2(new_n1005), .ZN(new_n1007));
  AND3_X1   g871(.A1(new_n1006), .A2(new_n969), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g872(.A(new_n969), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1009));
  NOR2_X1   g873(.A1(new_n1008), .A2(new_n1009), .ZN(G402));
endmodule


