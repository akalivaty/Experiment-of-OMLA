

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783;

  BUF_X1 U367 ( .A(n633), .Z(n693) );
  AND2_X1 U368 ( .A1(n374), .A2(n373), .ZN(n372) );
  OR2_X1 U369 ( .A1(n547), .A2(KEYINPUT0), .ZN(n374) );
  XNOR2_X1 U370 ( .A(n458), .B(n459), .ZN(n462) );
  XNOR2_X1 U371 ( .A(n498), .B(KEYINPUT10), .ZN(n516) );
  BUF_X1 U372 ( .A(G128), .Z(n345) );
  INV_X1 U373 ( .A(G953), .ZN(n757) );
  AND2_X2 U374 ( .A1(n388), .A2(n355), .ZN(n391) );
  OR2_X2 U375 ( .A1(n703), .A2(G902), .ZN(n424) );
  XNOR2_X2 U376 ( .A(n466), .B(n483), .ZN(n703) );
  XNOR2_X1 U377 ( .A(G107), .B(G116), .ZN(n524) );
  XNOR2_X1 U378 ( .A(n596), .B(n595), .ZN(n683) );
  XNOR2_X2 U379 ( .A(n426), .B(n349), .ZN(n454) );
  XNOR2_X2 U380 ( .A(n506), .B(n350), .ZN(n381) );
  AND2_X1 U381 ( .A1(n368), .A2(n357), .ZN(n366) );
  XNOR2_X1 U382 ( .A(n375), .B(KEYINPUT22), .ZN(n559) );
  INV_X1 U383 ( .A(n618), .ZN(n567) );
  INV_X1 U384 ( .A(G134), .ZN(n456) );
  INV_X1 U385 ( .A(KEYINPUT39), .ZN(n397) );
  NOR2_X1 U386 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U387 ( .A1(n366), .A2(n369), .ZN(n365) );
  INV_X1 U388 ( .A(n559), .ZN(n419) );
  NOR2_X1 U389 ( .A1(n537), .A2(n717), .ZN(n398) );
  NAND2_X2 U390 ( .A1(n372), .A2(n370), .ZN(n625) );
  XNOR2_X1 U391 ( .A(KEYINPUT91), .B(G110), .ZN(n489) );
  XNOR2_X1 U392 ( .A(G104), .B(G122), .ZN(n514) );
  INV_X1 U393 ( .A(n646), .ZN(n411) );
  XNOR2_X2 U394 ( .A(n609), .B(G146), .ZN(n483) );
  NOR2_X1 U395 ( .A1(n384), .A2(n627), .ZN(n379) );
  NAND2_X1 U396 ( .A1(n367), .A2(n365), .ZN(n642) );
  NAND2_X1 U397 ( .A1(n392), .A2(KEYINPUT34), .ZN(n387) );
  NAND2_X1 U398 ( .A1(n625), .A2(n347), .ZN(n375) );
  NOR2_X1 U399 ( .A1(n628), .A2(n386), .ZN(n629) );
  NOR2_X1 U400 ( .A1(n626), .A2(KEYINPUT100), .ZN(n385) );
  AND2_X1 U401 ( .A1(n639), .A2(n641), .ZN(n369) );
  AND2_X1 U402 ( .A1(n733), .A2(n718), .ZN(n487) );
  INV_X1 U403 ( .A(KEYINPUT110), .ZN(n468) );
  INV_X1 U404 ( .A(G902), .ZN(n533) );
  XNOR2_X1 U405 ( .A(n360), .B(n442), .ZN(n656) );
  XNOR2_X1 U406 ( .A(n608), .B(n441), .ZN(n360) );
  NAND2_X1 U407 ( .A1(n411), .A2(n660), .ZN(n715) );
  AND2_X1 U408 ( .A1(n541), .A2(n733), .ZN(n741) );
  NOR2_X1 U409 ( .A1(n579), .A2(n417), .ZN(n416) );
  NOR2_X1 U410 ( .A1(n383), .A2(n723), .ZN(n382) );
  NOR2_X1 U411 ( .A1(n766), .A2(KEYINPUT100), .ZN(n383) );
  INV_X1 U412 ( .A(KEYINPUT46), .ZN(n428) );
  NAND2_X1 U413 ( .A1(n407), .A2(n405), .ZN(n404) );
  NAND2_X1 U414 ( .A1(n657), .A2(KEYINPUT64), .ZN(n407) );
  NAND2_X1 U415 ( .A1(n409), .A2(n406), .ZN(n405) );
  NAND2_X1 U416 ( .A1(KEYINPUT2), .A2(KEYINPUT64), .ZN(n406) );
  NOR2_X1 U417 ( .A1(G953), .A2(G237), .ZN(n507) );
  NAND2_X1 U418 ( .A1(G953), .A2(G902), .ZN(n542) );
  XNOR2_X1 U419 ( .A(G137), .B(G116), .ZN(n478) );
  XNOR2_X1 U420 ( .A(G119), .B(G113), .ZN(n363) );
  XNOR2_X1 U421 ( .A(KEYINPUT24), .B(KEYINPUT82), .ZN(n435) );
  XNOR2_X1 U422 ( .A(G110), .B(KEYINPUT94), .ZN(n436) );
  XNOR2_X1 U423 ( .A(KEYINPUT23), .B(KEYINPUT73), .ZN(n433) );
  XNOR2_X1 U424 ( .A(G119), .B(KEYINPUT93), .ZN(n425) );
  XNOR2_X1 U425 ( .A(G140), .B(G113), .ZN(n511) );
  XOR2_X1 U426 ( .A(G131), .B(G143), .Z(n512) );
  INV_X1 U427 ( .A(G140), .ZN(n443) );
  XNOR2_X1 U428 ( .A(KEYINPUT92), .B(KEYINPUT78), .ZN(n495) );
  XOR2_X1 U429 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n496) );
  INV_X1 U430 ( .A(KEYINPUT38), .ZN(n380) );
  XNOR2_X1 U431 ( .A(n584), .B(KEYINPUT1), .ZN(n554) );
  OR2_X1 U432 ( .A1(n432), .A2(KEYINPUT0), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n362), .B(n361), .ZN(n493) );
  XNOR2_X1 U434 ( .A(G101), .B(KEYINPUT71), .ZN(n361) );
  XNOR2_X1 U435 ( .A(n481), .B(n363), .ZN(n362) );
  XNOR2_X1 U436 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n481) );
  XNOR2_X1 U437 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n490) );
  XOR2_X1 U438 ( .A(G134), .B(KEYINPUT103), .Z(n522) );
  NAND2_X1 U439 ( .A1(n403), .A2(n402), .ZN(n667) );
  XNOR2_X1 U440 ( .A(G101), .B(G107), .ZN(n459) );
  XNOR2_X1 U441 ( .A(G104), .B(KEYINPUT77), .ZN(n463) );
  NAND2_X1 U442 ( .A1(n390), .A2(KEYINPUT34), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n623), .B(n468), .ZN(n431) );
  NAND2_X1 U444 ( .A1(n381), .A2(n718), .ZN(n576) );
  NAND2_X1 U445 ( .A1(n735), .A2(n584), .ZN(n623) );
  XNOR2_X1 U446 ( .A(n669), .B(n668), .ZN(n670) );
  INV_X1 U447 ( .A(n656), .ZN(n396) );
  NAND2_X1 U448 ( .A1(n667), .A2(n715), .ZN(n694) );
  XOR2_X1 U449 ( .A(n686), .B(KEYINPUT59), .Z(n687) );
  NAND2_X1 U450 ( .A1(n664), .A2(G953), .ZN(n699) );
  INV_X1 U451 ( .A(KEYINPUT31), .ZN(n378) );
  NAND2_X1 U452 ( .A1(n741), .A2(n625), .ZN(n548) );
  NOR2_X1 U453 ( .A1(n414), .A2(n353), .ZN(n413) );
  INV_X1 U454 ( .A(KEYINPUT53), .ZN(n393) );
  NAND2_X1 U455 ( .A1(n607), .A2(n606), .ZN(n710) );
  AND2_X1 U456 ( .A1(n658), .A2(n358), .ZN(n346) );
  INV_X1 U457 ( .A(KEYINPUT64), .ZN(n408) );
  INV_X1 U458 ( .A(KEYINPUT105), .ZN(n417) );
  NOR2_X1 U459 ( .A1(n721), .A2(n729), .ZN(n347) );
  NOR2_X1 U460 ( .A1(n553), .A2(n552), .ZN(n348) );
  XOR2_X1 U461 ( .A(n448), .B(n447), .Z(n349) );
  XNOR2_X1 U462 ( .A(n505), .B(KEYINPUT79), .ZN(n350) );
  XNOR2_X1 U463 ( .A(n733), .B(KEYINPUT6), .ZN(n618) );
  AND2_X1 U464 ( .A1(n781), .A2(n592), .ZN(n351) );
  AND2_X1 U465 ( .A1(n658), .A2(n404), .ZN(n352) );
  INV_X1 U466 ( .A(n579), .ZN(n560) );
  BUF_X1 U467 ( .A(n554), .Z(n579) );
  NAND2_X1 U468 ( .A1(n635), .A2(n555), .ZN(n353) );
  AND2_X1 U469 ( .A1(n625), .A2(n620), .ZN(n354) );
  AND2_X1 U470 ( .A1(n387), .A2(n348), .ZN(n355) );
  XNOR2_X1 U471 ( .A(n619), .B(KEYINPUT33), .ZN(n356) );
  OR2_X1 U472 ( .A1(n641), .A2(KEYINPUT44), .ZN(n357) );
  INV_X1 U473 ( .A(n657), .ZN(n409) );
  XNOR2_X1 U474 ( .A(G902), .B(KEYINPUT15), .ZN(n657) );
  AND2_X1 U475 ( .A1(n409), .A2(KEYINPUT64), .ZN(n358) );
  INV_X1 U476 ( .A(KEYINPUT2), .ZN(n410) );
  NAND2_X1 U477 ( .A1(n410), .A2(n408), .ZN(n359) );
  XNOR2_X1 U478 ( .A(n483), .B(n484), .ZN(n669) );
  NAND2_X1 U479 ( .A1(n379), .A2(n626), .ZN(n377) );
  NOR2_X1 U480 ( .A1(n385), .A2(n376), .ZN(n386) );
  INV_X1 U481 ( .A(n766), .ZN(n384) );
  XNOR2_X1 U482 ( .A(n427), .B(n603), .ZN(n607) );
  XNOR2_X1 U483 ( .A(n514), .B(n489), .ZN(n492) );
  NAND2_X1 U484 ( .A1(n602), .A2(n601), .ZN(n429) );
  AND2_X1 U485 ( .A1(n488), .A2(n563), .ZN(n430) );
  NAND2_X1 U486 ( .A1(n364), .A2(n637), .ZN(n368) );
  INV_X1 U487 ( .A(n693), .ZN(n364) );
  NAND2_X1 U488 ( .A1(n640), .A2(n357), .ZN(n367) );
  NAND2_X1 U489 ( .A1(n547), .A2(n371), .ZN(n370) );
  AND2_X1 U490 ( .A1(n432), .A2(KEYINPUT0), .ZN(n371) );
  NAND2_X1 U491 ( .A1(n382), .A2(n377), .ZN(n376) );
  XNOR2_X2 U492 ( .A(n548), .B(n378), .ZN(n626) );
  INV_X1 U493 ( .A(n381), .ZN(n574) );
  XNOR2_X1 U494 ( .A(n574), .B(n380), .ZN(n717) );
  NAND2_X1 U495 ( .A1(n348), .A2(n381), .ZN(n535) );
  XNOR2_X2 U496 ( .A(G146), .B(G125), .ZN(n498) );
  NAND2_X1 U497 ( .A1(n727), .A2(n354), .ZN(n388) );
  XNOR2_X2 U498 ( .A(n420), .B(n356), .ZN(n727) );
  NAND2_X2 U499 ( .A1(n391), .A2(n389), .ZN(n621) );
  INV_X1 U500 ( .A(n727), .ZN(n390) );
  INV_X1 U501 ( .A(n625), .ZN(n392) );
  INV_X1 U502 ( .A(n646), .ZN(n661) );
  NAND2_X1 U503 ( .A1(n411), .A2(n346), .ZN(n402) );
  INV_X1 U504 ( .A(n694), .ZN(n685) );
  XNOR2_X2 U505 ( .A(n645), .B(n644), .ZN(n646) );
  NAND2_X1 U506 ( .A1(n401), .A2(n400), .ZN(n403) );
  XNOR2_X1 U507 ( .A(n663), .B(n396), .ZN(n395) );
  XNOR2_X1 U508 ( .A(n394), .B(n393), .ZN(G75) );
  NAND2_X1 U509 ( .A1(n762), .A2(n761), .ZN(n394) );
  NAND2_X1 U510 ( .A1(n395), .A2(n699), .ZN(n665) );
  XNOR2_X1 U511 ( .A(n398), .B(n397), .ZN(n593) );
  XNOR2_X1 U512 ( .A(n455), .B(KEYINPUT67), .ZN(n538) );
  NAND2_X1 U513 ( .A1(n399), .A2(n351), .ZN(n427) );
  XNOR2_X1 U514 ( .A(n429), .B(n428), .ZN(n399) );
  NAND2_X1 U515 ( .A1(n404), .A2(n359), .ZN(n400) );
  NAND2_X1 U516 ( .A1(n661), .A2(n352), .ZN(n401) );
  XNOR2_X2 U517 ( .A(n576), .B(KEYINPUT19), .ZN(n547) );
  NAND2_X1 U518 ( .A1(n419), .A2(n560), .ZN(n634) );
  NOR2_X1 U519 ( .A1(n418), .A2(n412), .ZN(n684) );
  NAND2_X1 U520 ( .A1(n415), .A2(n413), .ZN(n412) );
  NOR2_X1 U521 ( .A1(n560), .A2(KEYINPUT105), .ZN(n414) );
  NAND2_X1 U522 ( .A1(n419), .A2(n416), .ZN(n415) );
  AND2_X1 U523 ( .A1(n559), .A2(n417), .ZN(n418) );
  NAND2_X1 U524 ( .A1(n421), .A2(n567), .ZN(n420) );
  XNOR2_X1 U525 ( .A(n617), .B(n422), .ZN(n421) );
  INV_X1 U526 ( .A(KEYINPUT106), .ZN(n422) );
  XNOR2_X2 U527 ( .A(n540), .B(n539), .ZN(n617) );
  XNOR2_X2 U528 ( .A(n501), .B(n457), .ZN(n609) );
  XNOR2_X2 U529 ( .A(n523), .B(n423), .ZN(n501) );
  XNOR2_X2 U530 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n423) );
  XNOR2_X2 U531 ( .A(G143), .B(G128), .ZN(n523) );
  XNOR2_X2 U532 ( .A(n424), .B(n467), .ZN(n584) );
  XNOR2_X1 U533 ( .A(n425), .B(n345), .ZN(n434) );
  INV_X1 U534 ( .A(n454), .ZN(n555) );
  NAND2_X1 U535 ( .A1(n656), .A2(n533), .ZN(n426) );
  NAND2_X1 U536 ( .A1(n431), .A2(n430), .ZN(n537) );
  BUF_X1 U537 ( .A(n538), .Z(n735) );
  NOR2_X1 U538 ( .A1(n752), .A2(n546), .ZN(n432) );
  INV_X1 U539 ( .A(KEYINPUT100), .ZN(n627) );
  INV_X1 U540 ( .A(KEYINPUT98), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n434), .B(n433), .ZN(n438) );
  XNOR2_X1 U544 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U545 ( .A(n438), .B(n437), .ZN(n442) );
  NAND2_X1 U546 ( .A1(n757), .A2(G234), .ZN(n439) );
  XNOR2_X1 U547 ( .A(n439), .B(KEYINPUT8), .ZN(n528) );
  INV_X1 U548 ( .A(G221), .ZN(n440) );
  OR2_X1 U549 ( .A1(n528), .A2(n440), .ZN(n441) );
  XNOR2_X1 U550 ( .A(n443), .B(G137), .ZN(n460) );
  XNOR2_X1 U551 ( .A(n516), .B(n460), .ZN(n608) );
  NAND2_X1 U552 ( .A1(n657), .A2(G234), .ZN(n444) );
  XNOR2_X1 U553 ( .A(n444), .B(KEYINPUT20), .ZN(n449) );
  AND2_X1 U554 ( .A1(n449), .A2(G217), .ZN(n448) );
  XNOR2_X1 U555 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n446) );
  XNOR2_X1 U556 ( .A(KEYINPUT25), .B(KEYINPUT76), .ZN(n445) );
  XNOR2_X1 U557 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U558 ( .A1(n449), .A2(G221), .ZN(n452) );
  INV_X1 U559 ( .A(KEYINPUT97), .ZN(n450) );
  XNOR2_X1 U560 ( .A(n450), .B(KEYINPUT21), .ZN(n451) );
  XNOR2_X1 U561 ( .A(n452), .B(n451), .ZN(n729) );
  INV_X1 U562 ( .A(n729), .ZN(n453) );
  NAND2_X1 U563 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U564 ( .A(n456), .B(G131), .ZN(n457) );
  NAND2_X1 U565 ( .A1(n757), .A2(G227), .ZN(n458) );
  INV_X1 U566 ( .A(n460), .ZN(n461) );
  XNOR2_X1 U567 ( .A(n462), .B(n461), .ZN(n465) );
  XNOR2_X1 U568 ( .A(n489), .B(n463), .ZN(n464) );
  XNOR2_X1 U569 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U570 ( .A(KEYINPUT70), .B(G469), .ZN(n467) );
  NAND2_X1 U571 ( .A1(G234), .A2(G237), .ZN(n470) );
  INV_X1 U572 ( .A(KEYINPUT14), .ZN(n469) );
  XNOR2_X1 U573 ( .A(n470), .B(n469), .ZN(n752) );
  NOR2_X1 U574 ( .A1(n752), .A2(n542), .ZN(n471) );
  XNOR2_X1 U575 ( .A(n471), .B(KEYINPUT107), .ZN(n472) );
  NOR2_X1 U576 ( .A1(G900), .A2(n472), .ZN(n474) );
  NAND2_X1 U577 ( .A1(n757), .A2(G952), .ZN(n545) );
  NOR2_X1 U578 ( .A1(n752), .A2(n545), .ZN(n473) );
  OR2_X1 U579 ( .A1(n474), .A2(n473), .ZN(n563) );
  XOR2_X1 U580 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n476) );
  NAND2_X1 U581 ( .A1(G210), .A2(n507), .ZN(n475) );
  XNOR2_X1 U582 ( .A(n476), .B(n475), .ZN(n480) );
  XNOR2_X1 U583 ( .A(n482), .B(n493), .ZN(n484) );
  NAND2_X1 U584 ( .A1(n669), .A2(n533), .ZN(n485) );
  XNOR2_X2 U585 ( .A(n485), .B(G472), .ZN(n733) );
  INV_X1 U586 ( .A(G237), .ZN(n486) );
  NAND2_X1 U587 ( .A1(n533), .A2(n486), .ZN(n504) );
  AND2_X1 U588 ( .A1(n504), .A2(G214), .ZN(n597) );
  INV_X1 U589 ( .A(n597), .ZN(n718) );
  XNOR2_X1 U590 ( .A(n487), .B(KEYINPUT30), .ZN(n488) );
  XNOR2_X1 U591 ( .A(n524), .B(n490), .ZN(n491) );
  XNOR2_X1 U592 ( .A(n492), .B(n491), .ZN(n494) );
  XNOR2_X1 U593 ( .A(n494), .B(n493), .ZN(n651) );
  XNOR2_X1 U594 ( .A(n496), .B(n495), .ZN(n500) );
  NAND2_X1 U595 ( .A1(n757), .A2(G224), .ZN(n497) );
  XNOR2_X1 U596 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U597 ( .A(n500), .B(n499), .ZN(n502) );
  XNOR2_X1 U598 ( .A(n501), .B(n502), .ZN(n503) );
  XNOR2_X1 U599 ( .A(n651), .B(n503), .ZN(n677) );
  NAND2_X1 U600 ( .A1(n677), .A2(n657), .ZN(n506) );
  NAND2_X1 U601 ( .A1(n504), .A2(G210), .ZN(n505) );
  XOR2_X1 U602 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n509) );
  NAND2_X1 U603 ( .A1(n507), .A2(G214), .ZN(n508) );
  XNOR2_X1 U604 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U605 ( .A(n510), .B(KEYINPUT12), .Z(n518) );
  XNOR2_X1 U606 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U607 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U608 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U609 ( .A(n518), .B(n517), .ZN(n686) );
  NAND2_X1 U610 ( .A1(n686), .A2(n533), .ZN(n520) );
  XNOR2_X1 U611 ( .A(KEYINPUT13), .B(G475), .ZN(n519) );
  XNOR2_X1 U612 ( .A(n520), .B(n519), .ZN(n553) );
  XNOR2_X1 U613 ( .A(G122), .B(KEYINPUT102), .ZN(n521) );
  XNOR2_X1 U614 ( .A(n522), .B(n521), .ZN(n526) );
  XNOR2_X1 U615 ( .A(n523), .B(n524), .ZN(n525) );
  XNOR2_X1 U616 ( .A(n526), .B(n525), .ZN(n532) );
  INV_X1 U617 ( .A(G217), .ZN(n527) );
  OR2_X1 U618 ( .A1(n528), .A2(n527), .ZN(n530) );
  XOR2_X1 U619 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n529) );
  XNOR2_X1 U620 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U621 ( .A(n532), .B(n531), .ZN(n697) );
  NAND2_X1 U622 ( .A1(n697), .A2(n533), .ZN(n534) );
  INV_X1 U623 ( .A(G478), .ZN(n695) );
  XNOR2_X1 U624 ( .A(n534), .B(n695), .ZN(n552) );
  OR2_X1 U625 ( .A1(n537), .A2(n535), .ZN(n590) );
  XOR2_X1 U626 ( .A(G143), .B(KEYINPUT115), .Z(n536) );
  XNOR2_X1 U627 ( .A(n590), .B(n536), .ZN(G45) );
  INV_X1 U628 ( .A(n552), .ZN(n549) );
  NAND2_X1 U629 ( .A1(n549), .A2(n553), .ZN(n765) );
  INV_X1 U630 ( .A(n765), .ZN(n771) );
  NAND2_X1 U631 ( .A1(n593), .A2(n771), .ZN(n605) );
  XNOR2_X1 U632 ( .A(n605), .B(G134), .ZN(G36) );
  NAND2_X1 U633 ( .A1(n538), .A2(n554), .ZN(n540) );
  INV_X1 U634 ( .A(KEYINPUT75), .ZN(n539) );
  INV_X1 U635 ( .A(n617), .ZN(n541) );
  INV_X1 U636 ( .A(G898), .ZN(n652) );
  INV_X1 U637 ( .A(n542), .ZN(n543) );
  NAND2_X1 U638 ( .A1(n652), .A2(n543), .ZN(n544) );
  AND2_X1 U639 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U640 ( .A1(n549), .A2(n553), .ZN(n763) );
  NOR2_X1 U641 ( .A1(n626), .A2(n763), .ZN(n550) );
  XOR2_X1 U642 ( .A(G113), .B(n550), .Z(G15) );
  NOR2_X1 U643 ( .A1(n626), .A2(n765), .ZN(n551) );
  XOR2_X1 U644 ( .A(G116), .B(n551), .Z(G18) );
  NAND2_X1 U645 ( .A1(n553), .A2(n552), .ZN(n721) );
  INV_X1 U646 ( .A(n555), .ZN(n561) );
  NOR2_X1 U647 ( .A1(n560), .A2(n561), .ZN(n556) );
  NAND2_X1 U648 ( .A1(n556), .A2(n618), .ZN(n557) );
  NOR2_X1 U649 ( .A1(n559), .A2(n557), .ZN(n558) );
  XNOR2_X1 U650 ( .A(n558), .B(KEYINPUT32), .ZN(n636) );
  XOR2_X1 U651 ( .A(G119), .B(n636), .Z(G21) );
  NAND2_X1 U652 ( .A1(n618), .A2(n561), .ZN(n562) );
  NOR2_X1 U653 ( .A1(n634), .A2(n562), .ZN(n628) );
  XOR2_X1 U654 ( .A(G101), .B(n628), .Z(G3) );
  INV_X1 U655 ( .A(n563), .ZN(n564) );
  NOR2_X1 U656 ( .A1(n729), .A2(n564), .ZN(n565) );
  XOR2_X1 U657 ( .A(n565), .B(KEYINPUT69), .Z(n566) );
  AND2_X1 U658 ( .A1(n555), .A2(n566), .ZN(n581) );
  NAND2_X1 U659 ( .A1(n567), .A2(n581), .ZN(n568) );
  XNOR2_X1 U660 ( .A(KEYINPUT108), .B(n568), .ZN(n569) );
  NOR2_X1 U661 ( .A1(n763), .A2(n569), .ZN(n570) );
  XNOR2_X1 U662 ( .A(KEYINPUT109), .B(n570), .ZN(n577) );
  INV_X1 U663 ( .A(n577), .ZN(n571) );
  NAND2_X1 U664 ( .A1(n718), .A2(n571), .ZN(n572) );
  OR2_X1 U665 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U666 ( .A(n573), .B(KEYINPUT43), .ZN(n575) );
  NAND2_X1 U667 ( .A1(n575), .A2(n574), .ZN(n604) );
  XNOR2_X1 U668 ( .A(n604), .B(G140), .ZN(G42) );
  NOR2_X1 U669 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U670 ( .A(n578), .B(KEYINPUT36), .ZN(n580) );
  NAND2_X1 U671 ( .A1(n580), .A2(n579), .ZN(n781) );
  NAND2_X1 U672 ( .A1(n733), .A2(n581), .ZN(n583) );
  XNOR2_X1 U673 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n582) );
  XNOR2_X1 U674 ( .A(n583), .B(n582), .ZN(n585) );
  AND2_X1 U675 ( .A1(n584), .A2(n585), .ZN(n770) );
  AND2_X1 U676 ( .A1(n763), .A2(n765), .ZN(n723) );
  INV_X1 U677 ( .A(n723), .ZN(n586) );
  AND2_X1 U678 ( .A1(n547), .A2(n586), .ZN(n587) );
  NAND2_X1 U679 ( .A1(n770), .A2(n587), .ZN(n589) );
  INV_X1 U680 ( .A(KEYINPUT47), .ZN(n588) );
  XNOR2_X1 U681 ( .A(n589), .B(n588), .ZN(n591) );
  AND2_X1 U682 ( .A1(n591), .A2(n590), .ZN(n592) );
  INV_X1 U683 ( .A(n763), .ZN(n775) );
  NAND2_X1 U684 ( .A1(n593), .A2(n775), .ZN(n596) );
  INV_X1 U685 ( .A(KEYINPUT112), .ZN(n594) );
  XNOR2_X1 U686 ( .A(n594), .B(KEYINPUT40), .ZN(n595) );
  INV_X1 U687 ( .A(n683), .ZN(n602) );
  OR2_X1 U688 ( .A1(n717), .A2(n597), .ZN(n722) );
  OR2_X1 U689 ( .A1(n722), .A2(n721), .ZN(n598) );
  XNOR2_X1 U690 ( .A(n598), .B(KEYINPUT41), .ZN(n756) );
  NAND2_X1 U691 ( .A1(n756), .A2(n770), .ZN(n600) );
  INV_X1 U692 ( .A(KEYINPUT42), .ZN(n599) );
  XNOR2_X1 U693 ( .A(n600), .B(n599), .ZN(n783) );
  INV_X1 U694 ( .A(n783), .ZN(n601) );
  INV_X1 U695 ( .A(KEYINPUT48), .ZN(n603) );
  AND2_X1 U696 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U697 ( .A(n609), .B(n608), .ZN(n612) );
  XNOR2_X1 U698 ( .A(n612), .B(KEYINPUT125), .ZN(n610) );
  XNOR2_X1 U699 ( .A(n710), .B(n610), .ZN(n611) );
  NAND2_X1 U700 ( .A1(n611), .A2(n757), .ZN(n616) );
  XOR2_X1 U701 ( .A(G227), .B(n612), .Z(n613) );
  NAND2_X1 U702 ( .A1(n613), .A2(G900), .ZN(n614) );
  NAND2_X1 U703 ( .A1(n614), .A2(G953), .ZN(n615) );
  NAND2_X1 U704 ( .A1(n616), .A2(n615), .ZN(G72) );
  INV_X1 U705 ( .A(KEYINPUT89), .ZN(n619) );
  INV_X1 U706 ( .A(KEYINPUT34), .ZN(n620) );
  XNOR2_X2 U707 ( .A(n621), .B(KEYINPUT35), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n633), .A2(KEYINPUT44), .ZN(n622) );
  XNOR2_X1 U709 ( .A(n622), .B(KEYINPUT88), .ZN(n631) );
  NOR2_X1 U710 ( .A1(n623), .A2(n733), .ZN(n624) );
  NAND2_X1 U711 ( .A1(n625), .A2(n624), .ZN(n766) );
  XNOR2_X1 U712 ( .A(n629), .B(KEYINPUT104), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U714 ( .A(n632), .B(KEYINPUT87), .ZN(n643) );
  INV_X1 U715 ( .A(n733), .ZN(n635) );
  NOR2_X1 U716 ( .A1(n684), .A2(n636), .ZN(n639) );
  INV_X1 U717 ( .A(KEYINPUT65), .ZN(n641) );
  INV_X1 U718 ( .A(KEYINPUT44), .ZN(n637) );
  NOR2_X1 U719 ( .A1(n637), .A2(KEYINPUT65), .ZN(n638) );
  NOR2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n645) );
  INV_X1 U722 ( .A(KEYINPUT45), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n411), .A2(n757), .ZN(n650) );
  NAND2_X1 U724 ( .A1(G953), .A2(G224), .ZN(n647) );
  XNOR2_X1 U725 ( .A(KEYINPUT61), .B(n647), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n648), .A2(G898), .ZN(n649) );
  NAND2_X1 U727 ( .A1(n650), .A2(n649), .ZN(n655) );
  AND2_X1 U728 ( .A1(n652), .A2(G953), .ZN(n653) );
  NOR2_X1 U729 ( .A1(n651), .A2(n653), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n655), .B(n654), .ZN(G69) );
  INV_X1 U731 ( .A(KEYINPUT124), .ZN(n666) );
  INV_X1 U732 ( .A(n710), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n658), .A2(KEYINPUT2), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n659), .B(KEYINPUT85), .ZN(n660) );
  AND2_X1 U735 ( .A1(n715), .A2(G217), .ZN(n662) );
  AND2_X1 U736 ( .A1(n667), .A2(n662), .ZN(n663) );
  INV_X1 U737 ( .A(G952), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n666), .B(n665), .ZN(G66) );
  INV_X1 U739 ( .A(n694), .ZN(n701) );
  NAND2_X1 U740 ( .A1(n701), .A2(G472), .ZN(n671) );
  XOR2_X1 U741 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n668) );
  XNOR2_X1 U742 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U743 ( .A1(n672), .A2(n699), .ZN(n675) );
  XNOR2_X1 U744 ( .A(KEYINPUT114), .B(KEYINPUT63), .ZN(n673) );
  XNOR2_X1 U745 ( .A(n673), .B(KEYINPUT90), .ZN(n674) );
  XNOR2_X1 U746 ( .A(n675), .B(n674), .ZN(G57) );
  NAND2_X1 U747 ( .A1(n685), .A2(G210), .ZN(n679) );
  XOR2_X1 U748 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n676) );
  XNOR2_X1 U749 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U750 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U751 ( .A1(n680), .A2(n699), .ZN(n682) );
  XOR2_X1 U752 ( .A(KEYINPUT86), .B(KEYINPUT56), .Z(n681) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(G51) );
  XOR2_X1 U754 ( .A(n683), .B(G131), .Z(G33) );
  XOR2_X1 U755 ( .A(n684), .B(G110), .Z(G12) );
  NAND2_X1 U756 ( .A1(n701), .A2(G475), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n688), .B(n687), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n689), .A2(n699), .ZN(n691) );
  XOR2_X1 U759 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n690) );
  XNOR2_X1 U760 ( .A(n691), .B(n690), .ZN(G60) );
  XOR2_X1 U761 ( .A(G122), .B(KEYINPUT126), .Z(n692) );
  XNOR2_X1 U762 ( .A(n693), .B(n692), .ZN(G24) );
  BUF_X1 U763 ( .A(n694), .Z(n696) );
  NOR2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n698) );
  XNOR2_X1 U765 ( .A(n698), .B(n697), .ZN(n700) );
  INV_X1 U766 ( .A(n699), .ZN(n706) );
  NOR2_X1 U767 ( .A1(n700), .A2(n706), .ZN(G63) );
  NAND2_X1 U768 ( .A1(n685), .A2(G469), .ZN(n705) );
  XOR2_X1 U769 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n702) );
  XNOR2_X1 U770 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U771 ( .A(n705), .B(n704), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n707), .A2(n706), .ZN(G54) );
  XNOR2_X1 U773 ( .A(KEYINPUT2), .B(KEYINPUT81), .ZN(n709) );
  NAND2_X1 U774 ( .A1(n646), .A2(n709), .ZN(n708) );
  XNOR2_X1 U775 ( .A(n708), .B(KEYINPUT83), .ZN(n713) );
  NAND2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U777 ( .A(KEYINPUT84), .B(n711), .Z(n712) );
  XNOR2_X1 U778 ( .A(n714), .B(KEYINPUT80), .ZN(n716) );
  NAND2_X1 U779 ( .A1(n716), .A2(n715), .ZN(n762) );
  INV_X1 U780 ( .A(n717), .ZN(n719) );
  NOR2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n725) );
  NOR2_X1 U783 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U784 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U785 ( .A(n726), .B(KEYINPUT122), .ZN(n728) );
  NOR2_X1 U786 ( .A1(n728), .A2(n390), .ZN(n749) );
  NAND2_X1 U787 ( .A1(n555), .A2(n729), .ZN(n730) );
  XNOR2_X1 U788 ( .A(n730), .B(KEYINPUT49), .ZN(n731) );
  XNOR2_X1 U789 ( .A(n731), .B(KEYINPUT118), .ZN(n732) );
  NOR2_X1 U790 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U791 ( .A(KEYINPUT119), .B(n734), .Z(n740) );
  INV_X1 U792 ( .A(n735), .ZN(n736) );
  NAND2_X1 U793 ( .A1(n560), .A2(n736), .ZN(n737) );
  XNOR2_X1 U794 ( .A(n737), .B(KEYINPUT50), .ZN(n738) );
  XNOR2_X1 U795 ( .A(KEYINPUT120), .B(n738), .ZN(n739) );
  NAND2_X1 U796 ( .A1(n740), .A2(n739), .ZN(n743) );
  INV_X1 U797 ( .A(n741), .ZN(n742) );
  NAND2_X1 U798 ( .A1(n743), .A2(n742), .ZN(n745) );
  XOR2_X1 U799 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n744) );
  XNOR2_X1 U800 ( .A(n745), .B(n744), .ZN(n747) );
  INV_X1 U801 ( .A(n756), .ZN(n746) );
  NOR2_X1 U802 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U803 ( .A1(n749), .A2(n748), .ZN(n751) );
  XOR2_X1 U804 ( .A(KEYINPUT123), .B(KEYINPUT52), .Z(n750) );
  XNOR2_X1 U805 ( .A(n751), .B(n750), .ZN(n755) );
  INV_X1 U806 ( .A(n752), .ZN(n753) );
  NAND2_X1 U807 ( .A1(n753), .A2(G952), .ZN(n754) );
  NOR2_X1 U808 ( .A1(n755), .A2(n754), .ZN(n760) );
  NAND2_X1 U809 ( .A1(n727), .A2(n756), .ZN(n758) );
  NAND2_X1 U810 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U811 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U812 ( .A1(n766), .A2(n763), .ZN(n764) );
  XOR2_X1 U813 ( .A(G104), .B(n764), .Z(G6) );
  NOR2_X1 U814 ( .A1(n766), .A2(n765), .ZN(n768) );
  XNOR2_X1 U815 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n767) );
  XNOR2_X1 U816 ( .A(n768), .B(n767), .ZN(n769) );
  XNOR2_X1 U817 ( .A(G107), .B(n769), .ZN(G9) );
  INV_X1 U818 ( .A(n770), .ZN(n777) );
  NAND2_X1 U819 ( .A1(n547), .A2(n771), .ZN(n772) );
  NOR2_X1 U820 ( .A1(n777), .A2(n772), .ZN(n774) );
  XNOR2_X1 U821 ( .A(n345), .B(KEYINPUT29), .ZN(n773) );
  XNOR2_X1 U822 ( .A(n774), .B(n773), .ZN(G30) );
  NAND2_X1 U823 ( .A1(n547), .A2(n775), .ZN(n776) );
  NOR2_X1 U824 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U825 ( .A(KEYINPUT116), .B(n778), .Z(n779) );
  XNOR2_X1 U826 ( .A(G146), .B(n779), .ZN(G48) );
  XNOR2_X1 U827 ( .A(KEYINPUT37), .B(KEYINPUT117), .ZN(n780) );
  XNOR2_X1 U828 ( .A(n781), .B(n780), .ZN(n782) );
  XNOR2_X1 U829 ( .A(G125), .B(n782), .ZN(G27) );
  XOR2_X1 U830 ( .A(G137), .B(n783), .Z(G39) );
endmodule

