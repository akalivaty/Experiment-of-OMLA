//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1315, new_n1316, new_n1317, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1346, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1413,
    new_n1414, new_n1415;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND3_X1  g0010(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(new_n203), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n203), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n207), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n210), .B1(new_n211), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT64), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G58), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(G13), .ZN(new_n245));
  INV_X1    g0045(.A(G20), .ZN(new_n246));
  NOR3_X1   g0046(.A1(new_n245), .A2(new_n246), .A3(G1), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G1), .A2(G13), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n201), .B1(new_n252), .B2(G20), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n251), .A2(new_n253), .B1(new_n201), .B2(new_n247), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n246), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n246), .A2(new_n258), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n255), .A2(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n260), .B1(G20), .B2(new_n204), .ZN(new_n261));
  INV_X1    g0061(.A(new_n250), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n254), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT9), .ZN(new_n264));
  INV_X1    g0064(.A(G200), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  OAI211_X1 g0068(.A(G1), .B(G13), .C1(new_n258), .C2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(new_n269), .A3(G274), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT65), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n252), .B(KEYINPUT65), .C1(G41), .C2(G45), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G226), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT66), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT66), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G223), .A3(G1698), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G222), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n286), .B1(new_n220), .B2(new_n285), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n269), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n276), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n264), .B1(new_n265), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n294), .A2(G190), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n263), .B1(new_n294), .B2(G169), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n283), .B1(new_n281), .B2(new_n282), .ZN(new_n306));
  OAI211_X1 g0106(.A(G232), .B(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(G226), .B(new_n289), .C1(new_n305), .C2(new_n306), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G97), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n293), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n270), .B1(new_n274), .B2(new_n215), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT13), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n311), .A2(new_n316), .A3(new_n313), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G200), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n311), .B2(new_n313), .ZN(new_n320));
  AOI211_X1 g0120(.A(KEYINPUT13), .B(new_n312), .C1(new_n310), .C2(new_n293), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G190), .ZN(new_n323));
  INV_X1    g0123(.A(new_n259), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n220), .B2(new_n256), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n326), .A2(new_n250), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n328));
  INV_X1    g0128(.A(new_n247), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n262), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT68), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n252), .A2(G20), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(G68), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n247), .A2(new_n203), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT12), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n328), .A2(new_n336), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n319), .A2(new_n323), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n315), .A2(G179), .A3(new_n317), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT70), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT70), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n322), .A2(new_n346), .A3(G179), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(G169), .C1(new_n320), .C2(new_n321), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT69), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT14), .B1(new_n322), .B2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n318), .A2(KEYINPUT69), .A3(new_n349), .A4(G169), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n348), .A2(new_n352), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n343), .B1(new_n356), .B2(new_n340), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT76), .ZN(new_n358));
  INV_X1    g0158(.A(new_n255), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n335), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n360), .A2(new_n330), .B1(new_n329), .B2(new_n359), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT16), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT73), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n278), .A2(KEYINPUT73), .A3(G33), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n282), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT74), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n371), .A3(new_n368), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n280), .A2(new_n246), .A3(new_n284), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n367), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n203), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G58), .A2(G68), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n246), .B1(new_n212), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G159), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n259), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n362), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT71), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n278), .B2(G33), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n258), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(G20), .B1(new_n387), .B2(new_n281), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n203), .B1(new_n388), .B2(new_n367), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n277), .B1(new_n385), .B2(new_n386), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT7), .B1(new_n390), .B2(G20), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT72), .B1(new_n378), .B2(new_n380), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n381), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n389), .A2(new_n391), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n262), .B1(new_n395), .B2(KEYINPUT16), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n361), .B1(new_n383), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n272), .A2(G232), .A3(new_n269), .A4(new_n273), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n270), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(KEYINPUT75), .A3(new_n270), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  XNOR2_X1  g0205(.A(KEYINPUT67), .B(G1698), .ZN(new_n406));
  INV_X1    g0206(.A(G223), .ZN(new_n407));
  INV_X1    g0207(.A(G1698), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n406), .A2(new_n407), .B1(new_n275), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n405), .B1(new_n409), .B2(new_n390), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n300), .B1(new_n410), .B2(new_n269), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n403), .A2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n289), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n387), .A2(new_n281), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n404), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n293), .ZN(new_n416));
  INV_X1    g0216(.A(new_n399), .ZN(new_n417));
  AOI21_X1  g0217(.A(G169), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT18), .B1(new_n397), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n361), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n366), .A2(new_n371), .A3(new_n368), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n371), .B1(new_n366), .B2(new_n368), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n305), .A2(new_n306), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT7), .B1(new_n426), .B2(new_n246), .ZN(new_n427));
  OAI21_X1  g0227(.A(G68), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT16), .B1(new_n428), .B2(new_n381), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n388), .A2(new_n367), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(G68), .A3(new_n391), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n394), .A2(new_n392), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT16), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n250), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n422), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n419), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n358), .B1(new_n421), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  INV_X1    g0239(.A(G190), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n440), .A2(KEYINPUT77), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(KEYINPUT77), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n410), .B2(new_n269), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT78), .B1(new_n403), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n416), .A2(new_n417), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n265), .ZN(new_n447));
  INV_X1    g0247(.A(new_n443), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n415), .B2(new_n293), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT78), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(new_n401), .A4(new_n402), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n445), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n439), .B1(new_n435), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT76), .A2(KEYINPUT18), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n397), .B2(new_n420), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n445), .A2(new_n447), .A3(new_n451), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n438), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n285), .A2(G238), .A3(G1698), .ZN(new_n460));
  OAI221_X1 g0260(.A(new_n460), .B1(new_n222), .B2(new_n285), .C1(new_n290), .C2(new_n229), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n293), .ZN(new_n462));
  INV_X1    g0262(.A(new_n270), .ZN(new_n463));
  INV_X1    g0263(.A(new_n274), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(G244), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n300), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n334), .A2(G77), .A3(new_n335), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n255), .A2(new_n259), .B1(new_n246), .B2(new_n220), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT15), .B(G87), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n256), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n250), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n468), .B(new_n472), .C1(G77), .C2(new_n329), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n462), .A2(new_n465), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n353), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(G200), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n473), .B1(new_n466), .B2(G190), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n304), .A2(new_n357), .A3(new_n459), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT80), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n268), .A2(KEYINPUT5), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n252), .A2(G45), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G41), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(KEYINPUT80), .A3(new_n252), .A4(G45), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n268), .A2(KEYINPUT5), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G257), .A3(new_n269), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n252), .B(G45), .C1(new_n268), .C2(KEYINPUT5), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n492), .A2(new_n482), .B1(KEYINPUT5), .B2(new_n268), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(G274), .A3(new_n269), .A4(new_n488), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  OR2_X1    g0296(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n497));
  NAND2_X1  g0297(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n497), .A2(KEYINPUT4), .A3(G244), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G250), .A2(G1698), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n280), .A2(new_n284), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n287), .A2(new_n288), .A3(new_n221), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT4), .B1(new_n390), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n496), .B(G179), .C1(new_n506), .C2(new_n269), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n499), .A2(new_n500), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n285), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n503), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n269), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(G169), .B1(new_n511), .B2(new_n495), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n252), .A2(G33), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n251), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OR3_X1    g0316(.A1(new_n329), .A2(KEYINPUT79), .A3(G97), .ZN(new_n517));
  OAI21_X1  g0317(.A(KEYINPUT79), .B1(new_n329), .B2(G97), .ZN(new_n518));
  AOI22_X1  g0318(.A1(G97), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT6), .ZN(new_n520));
  INV_X1    g0320(.A(G97), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n521), .A2(new_n222), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G97), .A2(G107), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n222), .A2(KEYINPUT6), .A3(G97), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(G20), .B1(G77), .B2(new_n324), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n375), .B1(new_n423), .B2(new_n424), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(G107), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n519), .B1(new_n530), .B2(new_n262), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n513), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n496), .B(new_n440), .C1(new_n506), .C2(new_n269), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n265), .B1(new_n511), .B2(new_n495), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n519), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n370), .A2(new_n372), .B1(new_n374), .B2(new_n367), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n527), .B1(new_n537), .B2(new_n222), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n538), .B2(new_n250), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n532), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT81), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n490), .A2(KEYINPUT83), .A3(G270), .A4(new_n269), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n494), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n293), .B1(new_n493), .B2(new_n488), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT83), .B1(new_n546), .B2(G270), .ZN(new_n547));
  INV_X1    g0347(.A(G257), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n406), .A2(new_n548), .B1(new_n223), .B2(new_n408), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n390), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n280), .A2(G303), .A3(new_n284), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n269), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n545), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n514), .A2(G116), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n332), .A2(new_n333), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n245), .A2(G1), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G116), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G20), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n504), .B(new_n246), .C1(G33), .C2(new_n521), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(new_n250), .A3(new_n560), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT20), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n562), .A2(KEYINPUT20), .A3(new_n250), .A4(new_n560), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n561), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n556), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n553), .A2(G179), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n550), .A2(new_n551), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n293), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n490), .A2(G270), .A3(new_n269), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT83), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n571), .A2(new_n574), .A3(new_n494), .A4(new_n544), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT21), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n353), .B1(new_n556), .B2(new_n567), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n576), .B1(new_n575), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n569), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n568), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n575), .B2(new_n443), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n553), .A2(new_n265), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n532), .A2(new_n540), .A3(KEYINPUT81), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n484), .A2(G274), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n484), .A2(new_n217), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n269), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n258), .A2(new_n559), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n406), .A2(new_n215), .B1(new_n221), .B2(new_n408), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n390), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT82), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n293), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI211_X1 g0394(.A(KEYINPUT82), .B(new_n590), .C1(new_n591), .C2(new_n390), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n589), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n353), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n300), .B(new_n589), .C1(new_n594), .C2(new_n595), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n390), .A2(new_n246), .A3(G68), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT19), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n246), .B1(new_n309), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n523), .A2(new_n216), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n246), .A2(G33), .A3(G97), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n601), .A2(new_n602), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n605), .A2(new_n250), .B1(new_n247), .B2(new_n470), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n470), .B2(new_n515), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n597), .A2(new_n598), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n516), .A2(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(G190), .B(new_n589), .C1(new_n594), .C2(new_n595), .ZN(new_n612));
  INV_X1    g0412(.A(new_n589), .ZN(new_n613));
  INV_X1    g0413(.A(new_n590), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n289), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n414), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n269), .B1(new_n616), .B2(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n592), .A2(new_n593), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n613), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n611), .B(new_n612), .C1(new_n619), .C2(new_n265), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n608), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n543), .A2(new_n585), .A3(new_n586), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT24), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n390), .A2(new_n246), .A3(G87), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT22), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n216), .A2(KEYINPUT22), .A3(G20), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n285), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT23), .B1(new_n222), .B2(G20), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n222), .A2(KEYINPUT23), .A3(G20), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n630), .A2(new_n631), .B1(new_n590), .B2(new_n246), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n623), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n632), .ZN(new_n634));
  AOI211_X1 g0434(.A(KEYINPUT24), .B(new_n634), .C1(new_n625), .C2(new_n627), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n250), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n287), .A2(new_n288), .A3(new_n217), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n548), .A2(new_n408), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n390), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(G33), .A2(G294), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n293), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT85), .B1(new_n546), .B2(G264), .ZN(new_n643));
  AND4_X1   g0443(.A1(KEYINPUT85), .A2(new_n490), .A3(G264), .A4(new_n269), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n494), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G200), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n247), .A2(KEYINPUT25), .A3(new_n222), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT25), .B1(new_n247), .B2(new_n222), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n515), .A2(new_n222), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n269), .B1(new_n639), .B2(new_n640), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n490), .A2(G264), .A3(new_n269), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT85), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n546), .A2(KEYINPUT85), .A3(G264), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(G190), .A3(new_n494), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n636), .A2(new_n646), .A3(new_n651), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n645), .A2(G169), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT86), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n657), .A2(G179), .A3(new_n494), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n660), .B2(new_n662), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n628), .A2(new_n623), .A3(new_n632), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n624), .A2(KEYINPUT22), .B1(new_n285), .B2(new_n626), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT24), .B1(new_n667), .B2(new_n634), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n262), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT84), .B1(new_n669), .B2(new_n650), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT84), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n636), .A2(new_n671), .A3(new_n651), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  NOR4_X1   g0474(.A1(new_n481), .A2(new_n622), .A3(new_n659), .A4(new_n674), .ZN(G372));
  INV_X1    g0475(.A(new_n481), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT87), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n596), .A2(new_n677), .A3(new_n353), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n677), .B1(new_n596), .B2(new_n353), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n598), .B(new_n607), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n610), .A2(KEYINPUT88), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT88), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n606), .A2(new_n684), .A3(new_n609), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n596), .A2(G200), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(new_n687), .A3(new_n612), .ZN(new_n688));
  INV_X1    g0488(.A(new_n532), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n681), .A2(new_n682), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n608), .A2(new_n620), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT26), .B1(new_n691), .B2(new_n532), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n690), .A2(new_n681), .A3(new_n692), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n575), .A2(new_n581), .A3(new_n300), .ZN(new_n694));
  INV_X1    g0494(.A(new_n579), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n645), .A2(new_n300), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n353), .B1(new_n657), .B2(new_n494), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n698), .A2(new_n699), .B1(new_n669), .B2(new_n650), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(KEYINPUT89), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n688), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n598), .A2(new_n607), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n597), .A2(KEYINPUT87), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(new_n678), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n541), .A2(new_n659), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT89), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n636), .A2(new_n651), .B1(new_n660), .B2(new_n662), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n580), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n701), .A2(new_n706), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n693), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n676), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n303), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n421), .A2(new_n437), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n477), .B1(new_n356), .B2(new_n340), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n342), .A2(new_n453), .A3(new_n457), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n714), .B1(new_n718), .B2(new_n299), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n713), .A2(new_n719), .ZN(G369));
  INV_X1    g0520(.A(KEYINPUT93), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n557), .A2(new_n246), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n723));
  INV_X1    g0523(.A(G213), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT90), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT90), .B1(new_n722), .B2(KEYINPUT27), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT91), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n725), .B(KEYINPUT91), .C1(new_n728), .C2(new_n729), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(new_n733), .A3(G343), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n674), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n659), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n670), .A2(new_n672), .A3(new_n735), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n737), .B(new_n738), .C1(new_n665), .C2(new_n673), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n721), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n736), .A2(new_n721), .A3(new_n739), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT94), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n734), .A2(new_n581), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT92), .B1(new_n580), .B2(new_n745), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n569), .B1(new_n582), .B2(new_n583), .C1(new_n579), .C2(new_n578), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n746), .B1(new_n747), .B2(new_n745), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n580), .A2(KEYINPUT92), .A3(new_n745), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G330), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n743), .A2(new_n744), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n744), .B1(new_n743), .B2(new_n752), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n697), .A2(new_n735), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n736), .A2(new_n721), .A3(new_n739), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(new_n740), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n734), .B(KEYINPUT95), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n709), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n757), .A2(new_n765), .ZN(G399));
  INV_X1    g0566(.A(new_n208), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G41), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n602), .A2(G116), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(G1), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n213), .B2(new_n769), .ZN(new_n772));
  XOR2_X1   g0572(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n773));
  XNOR2_X1  g0573(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n586), .A2(new_n621), .ZN(new_n775));
  AOI21_X1  g0575(.A(KEYINPUT81), .B1(new_n532), .B2(new_n540), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n775), .A2(new_n747), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n670), .A2(new_n672), .ZN(new_n778));
  OAI21_X1  g0578(.A(KEYINPUT86), .B1(new_n698), .B2(new_n699), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n660), .A2(new_n662), .A3(new_n661), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n659), .B(new_n761), .C1(new_n778), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n777), .A2(new_n782), .A3(KEYINPUT98), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT98), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n737), .B(new_n762), .C1(new_n665), .C2(new_n673), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n622), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n511), .A2(new_n495), .A3(new_n300), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n788), .A2(new_n553), .A3(new_n619), .A4(new_n657), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT30), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n645), .A2(new_n575), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n300), .B1(new_n511), .B2(new_n495), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n619), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n789), .A2(new_n790), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  AND3_X1   g0594(.A1(new_n553), .A2(new_n619), .A3(new_n657), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT97), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n795), .A2(new_n796), .A3(KEYINPUT30), .A4(new_n788), .ZN(new_n797));
  OAI21_X1  g0597(.A(KEYINPUT97), .B1(new_n789), .B2(new_n790), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n794), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(KEYINPUT31), .B1(new_n799), .B2(new_n735), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT31), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n762), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n800), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n751), .B1(new_n787), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n706), .A2(new_n707), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n580), .B1(new_n778), .B2(new_n781), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n689), .A2(new_n682), .A3(new_n608), .A4(new_n620), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n681), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n681), .A2(new_n689), .A3(new_n688), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(KEYINPUT26), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n735), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT29), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n712), .A2(new_n762), .ZN(new_n814));
  XOR2_X1   g0614(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n804), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n774), .B1(new_n817), .B2(G1), .ZN(G364));
  NOR2_X1   g0618(.A1(new_n245), .A2(G20), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n252), .B1(new_n819), .B2(G45), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n768), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n752), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n750), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(G330), .ZN(new_n826));
  NOR2_X1   g0626(.A1(G13), .A2(G33), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(G20), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n750), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n822), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n426), .A2(new_n767), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G355), .B1(new_n559), .B2(new_n767), .ZN(new_n833));
  INV_X1    g0633(.A(G45), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n243), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n390), .A2(new_n767), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(G45), .B2(new_n213), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(G20), .B1(KEYINPUT100), .B2(G169), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(KEYINPUT100), .A2(G169), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n249), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n829), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n831), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n440), .A2(G179), .A3(G200), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n246), .ZN(new_n846));
  INV_X1    g0646(.A(G294), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n246), .A2(new_n300), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n265), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n443), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(G326), .ZN(new_n854));
  INV_X1    g0654(.A(G322), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n443), .A2(G200), .A3(new_n850), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n854), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n852), .A2(G190), .ZN(new_n859));
  XNOR2_X1  g0659(.A(KEYINPUT33), .B(G317), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n848), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n246), .A2(G179), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(new_n440), .A3(G200), .ZN(new_n863));
  INV_X1    g0663(.A(G283), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(G190), .A3(G200), .ZN(new_n865));
  INV_X1    g0665(.A(G303), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n863), .A2(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(G311), .ZN(new_n868));
  NOR2_X1   g0668(.A1(G190), .A2(G200), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n849), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n426), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n862), .A2(new_n869), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n872), .A2(KEYINPUT101), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(KEYINPUT101), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n867), .B(new_n871), .C1(G329), .C2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n853), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n878), .A2(new_n201), .B1(new_n216), .B2(new_n865), .ZN(new_n879));
  INV_X1    g0679(.A(new_n859), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n880), .A2(new_n203), .B1(new_n222), .B2(new_n863), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n285), .B1(new_n220), .B2(new_n870), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n857), .A2(new_n202), .B1(new_n521), .B2(new_n846), .ZN(new_n883));
  NOR4_X1   g0683(.A1(new_n879), .A2(new_n881), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n875), .A2(new_n379), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT32), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n861), .A2(new_n877), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n842), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n844), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n824), .A2(new_n826), .B1(new_n830), .B2(new_n889), .ZN(G396));
  INV_X1    g0690(.A(new_n804), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n761), .B1(new_n693), .B2(new_n711), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n467), .A2(new_n473), .A3(new_n475), .A4(new_n734), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n479), .A2(new_n478), .B1(new_n473), .B2(new_n735), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(new_n477), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n761), .B(new_n895), .C1(new_n693), .C2(new_n711), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n891), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n899), .A2(KEYINPUT104), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n891), .A2(new_n897), .A3(new_n898), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n900), .A2(new_n822), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(KEYINPUT104), .B2(new_n899), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n888), .A2(new_n828), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT102), .Z(new_n905));
  OAI21_X1  g0705(.A(new_n822), .B1(new_n905), .B2(G77), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT103), .Z(new_n907));
  AOI22_X1  g0707(.A1(new_n853), .A2(G137), .B1(G143), .B2(new_n856), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n908), .B1(new_n257), .B2(new_n880), .C1(new_n379), .C2(new_n870), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT34), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n390), .B1(new_n201), .B2(new_n865), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n846), .A2(new_n202), .B1(new_n863), .B2(new_n203), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(new_n876), .C2(G132), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n910), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n846), .A2(new_n521), .B1(new_n863), .B2(new_n216), .ZN(new_n917));
  INV_X1    g0717(.A(new_n870), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n285), .B(new_n917), .C1(G116), .C2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(G303), .A2(new_n853), .B1(new_n859), .B2(G283), .ZN(new_n920));
  INV_X1    g0720(.A(new_n865), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n856), .A2(G294), .B1(G107), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n876), .A2(G311), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n919), .A2(new_n920), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n907), .B1(new_n888), .B2(new_n925), .C1(new_n896), .C2(new_n828), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n903), .A2(new_n926), .ZN(G384));
  NOR2_X1   g0727(.A1(new_n819), .A2(new_n252), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n676), .A2(new_n813), .A3(new_n816), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n719), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT107), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n346), .B1(new_n322), .B2(G179), .ZN(new_n932));
  NOR4_X1   g0732(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT70), .A4(new_n300), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n355), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n352), .A2(new_n354), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n340), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n341), .A2(new_n734), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(new_n342), .A3(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n340), .B(new_n735), .C1(new_n356), .C2(new_n343), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n893), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n941), .B1(new_n898), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT16), .B1(new_n431), .B2(new_n432), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n422), .B1(new_n434), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n732), .A2(new_n733), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n438), .B2(new_n458), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n946), .B1(new_n412), .B2(new_n418), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n397), .A2(new_n456), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT37), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT106), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n383), .A2(new_n396), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n456), .A3(new_n422), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n945), .A2(new_n950), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT106), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT37), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n435), .A2(new_n419), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n435), .A2(new_n947), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n960), .A2(new_n961), .A3(new_n952), .A4(new_n955), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n953), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n949), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT38), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n949), .A2(new_n963), .A3(KEYINPUT38), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n943), .A2(new_n968), .B1(new_n715), .B2(new_n947), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n960), .A2(new_n961), .A3(new_n955), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(KEYINPUT37), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n453), .A2(new_n421), .A3(new_n437), .A4(new_n457), .ZN(new_n972));
  INV_X1    g0772(.A(new_n961), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n971), .A2(new_n962), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n967), .B1(KEYINPUT38), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT39), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n966), .A2(KEYINPUT39), .A3(new_n967), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n356), .A2(new_n340), .A3(new_n734), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n969), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n931), .B(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n799), .A2(KEYINPUT31), .A3(new_n735), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n800), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT98), .B1(new_n777), .B2(new_n782), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n622), .A2(new_n785), .A3(new_n784), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n895), .B1(new_n939), .B2(new_n940), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n949), .A2(new_n963), .A3(KEYINPUT38), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n971), .A2(new_n962), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n972), .A2(new_n973), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT38), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT40), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT109), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT40), .ZN(new_n998));
  INV_X1    g0798(.A(new_n995), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n998), .B1(new_n999), .B2(new_n967), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT109), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n1000), .A2(new_n1001), .A3(new_n990), .A4(new_n989), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n966), .A2(new_n967), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(new_n989), .A3(new_n990), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n997), .A2(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n799), .A2(new_n735), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n801), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n984), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n786), .B2(new_n783), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(new_n481), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n751), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n928), .B1(new_n983), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n983), .B2(new_n1013), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n211), .A2(new_n559), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n526), .B(KEYINPUT105), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT35), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n1019), .B2(new_n1018), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT36), .Z(new_n1022));
  NAND2_X1  g0822(.A1(new_n377), .A2(G77), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n213), .A2(new_n1023), .B1(G50), .B2(new_n203), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1024), .A2(G1), .A3(new_n245), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1015), .A2(new_n1022), .A3(new_n1025), .ZN(G367));
  OAI211_X1 g0826(.A(new_n532), .B(new_n540), .C1(new_n762), .C2(new_n539), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n689), .A2(new_n761), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n757), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n706), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n686), .A2(new_n734), .ZN(new_n1033));
  MUX2_X1   g0833(.A(new_n1032), .B(new_n681), .S(new_n1033), .Z(new_n1034));
  INV_X1    g0834(.A(KEYINPUT43), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n674), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n532), .B1(new_n1038), .B2(new_n1027), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n762), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n758), .B(new_n1029), .C1(new_n759), .C2(new_n740), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT110), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT42), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1040), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1041), .B(KEYINPUT110), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1046), .A2(KEYINPUT42), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1036), .B(new_n1037), .C1(new_n1045), .C2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1046), .A2(KEYINPUT42), .B1(new_n762), .B2(new_n1039), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1049), .A2(new_n1035), .A3(new_n1034), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1031), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1048), .A2(new_n1051), .A3(new_n1031), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT111), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT111), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1048), .A2(new_n1051), .A3(new_n1055), .A4(new_n1031), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1052), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n820), .B(KEYINPUT116), .Z(new_n1058));
  INV_X1    g0858(.A(new_n817), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT115), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n760), .A2(new_n763), .A3(new_n1029), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1061), .B(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(KEYINPUT44), .B1(new_n764), .B2(new_n1030), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT44), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1066), .B(new_n1029), .C1(new_n760), .C2(new_n763), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n757), .B(new_n1060), .C1(new_n1064), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1065), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1067), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1061), .B(new_n1062), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1060), .B1(new_n754), .B2(new_n755), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n755), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(KEYINPUT115), .A3(new_n753), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1069), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n741), .B(new_n742), .C1(new_n697), .C2(new_n735), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n760), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT114), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT113), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1081), .B1(new_n752), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1081), .B2(new_n752), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1083), .B1(new_n1079), .B2(new_n760), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n817), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1059), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n768), .B(KEYINPUT41), .Z(new_n1090));
  OAI21_X1  g0890(.A(new_n1058), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1057), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1034), .A2(new_n829), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n836), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n843), .B1(new_n208), .B2(new_n470), .C1(new_n235), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n831), .B1(new_n1095), .B2(KEYINPUT117), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(KEYINPUT117), .B2(new_n1095), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n880), .A2(new_n847), .B1(new_n222), .B2(new_n846), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G303), .B2(new_n856), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n876), .A2(G317), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n863), .A2(new_n521), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n414), .B1(new_n864), .B2(new_n870), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n853), .C2(G311), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n921), .A2(G116), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT46), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1099), .A2(new_n1100), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n876), .A2(G137), .B1(G58), .B2(new_n921), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(KEYINPUT118), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n857), .A2(new_n257), .B1(new_n220), .B2(new_n863), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n846), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1109), .B1(G68), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(KEYINPUT118), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n426), .B1(G50), .B2(new_n918), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G143), .A2(new_n853), .B1(new_n859), .B2(G159), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1106), .B1(new_n1108), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT47), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1097), .B1(new_n1117), .B2(new_n842), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1093), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1092), .A2(new_n1119), .ZN(G387));
  INV_X1    g0920(.A(new_n1086), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1059), .B(new_n1121), .C1(new_n1080), .C2(new_n1084), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n768), .A3(new_n1087), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n859), .A2(new_n359), .B1(G68), .B2(new_n918), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT120), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n856), .A2(G50), .B1(G77), .B2(new_n921), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n470), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n853), .A2(G159), .B1(new_n1127), .B2(new_n1110), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n414), .B(new_n1101), .C1(new_n876), .C2(G150), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n846), .A2(new_n864), .B1(new_n865), .B2(new_n847), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n853), .A2(G322), .B1(G317), .B2(new_n856), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n866), .B2(new_n870), .C1(new_n868), .C2(new_n880), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT48), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1134), .B2(new_n1133), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT49), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n414), .B1(new_n559), .B2(new_n863), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n876), .B2(G326), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1130), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n842), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n232), .A2(new_n834), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n770), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1144), .A2(new_n836), .B1(new_n1145), .B2(new_n832), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT119), .B(KEYINPUT50), .Z(new_n1147));
  AND3_X1   g0947(.A1(new_n359), .A2(new_n201), .A3(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n770), .B(new_n834), .C1(new_n203), .C2(new_n220), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1147), .B1(new_n359), .B2(new_n201), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1146), .A2(new_n1151), .B1(G107), .B2(new_n208), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n831), .B1(new_n1152), .B2(new_n843), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1143), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n759), .A2(new_n740), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n829), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1121), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1058), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1123), .A2(new_n1159), .ZN(G393));
  NAND2_X1  g0960(.A1(new_n1078), .A2(new_n1088), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1069), .A2(new_n1077), .A3(new_n1087), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n768), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1030), .A2(new_n829), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n843), .B1(new_n521), .B2(new_n208), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n240), .B2(new_n836), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n853), .A2(G150), .B1(G159), .B2(new_n856), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT51), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n859), .A2(G50), .B1(G68), .B2(new_n921), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n863), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1110), .A2(G77), .B1(new_n1170), .B2(G87), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n876), .A2(G143), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n414), .B1(new_n359), .B2(new_n918), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1169), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n853), .A2(G317), .B1(G311), .B2(new_n856), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT52), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n859), .A2(G303), .B1(G107), .B2(new_n1170), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1110), .A2(G116), .B1(new_n921), .B2(G283), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n876), .A2(G322), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n285), .B1(G294), .B2(new_n918), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1168), .A2(new_n1174), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n831), .B(new_n1166), .C1(new_n1182), .C2(new_n842), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1078), .A2(new_n1158), .B1(new_n1164), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1163), .A2(new_n1184), .ZN(G390));
  NAND2_X1  g0985(.A1(new_n941), .A2(new_n896), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1010), .A2(new_n1186), .A3(new_n751), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n943), .A2(new_n980), .B1(new_n977), .B2(new_n978), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n975), .A2(new_n980), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n810), .A2(KEYINPUT26), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n681), .A3(new_n808), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n805), .A2(new_n806), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n734), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n894), .A2(new_n477), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n893), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1189), .B1(new_n1195), .B2(new_n941), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1187), .B1(new_n1188), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n942), .B1(new_n892), .B2(new_n896), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n941), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n980), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n979), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1195), .A2(new_n941), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1189), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n804), .A2(new_n896), .A3(new_n941), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1201), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1197), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n979), .A2(new_n827), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n822), .B1(new_n905), .B2(new_n359), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n853), .A2(G283), .B1(G77), .B2(new_n1110), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n222), .B2(new_n880), .C1(new_n559), .C2(new_n857), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n285), .B1(G97), .B2(new_n918), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n921), .A2(G87), .B1(new_n1170), .B2(G68), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n847), .C2(new_n875), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n426), .B1(new_n856), .B2(G132), .ZN(new_n1215));
  INV_X1    g1015(.A(G125), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(KEYINPUT54), .B(G143), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT122), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1215), .B1(new_n1216), .B2(new_n875), .C1(new_n870), .C2(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G128), .A2(new_n853), .B1(new_n859), .B2(G137), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n865), .A2(new_n257), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1110), .A2(G159), .B1(new_n1170), .B2(G50), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1221), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1211), .A2(new_n1214), .B1(new_n1220), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1209), .B1(new_n1227), .B2(new_n842), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1207), .A2(new_n1158), .B1(new_n1208), .B2(new_n1228), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1010), .A2(new_n481), .A3(new_n751), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n930), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n893), .B1(new_n814), .B2(new_n1194), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n803), .B1(new_n987), .B2(new_n988), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(G330), .A3(new_n896), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(KEYINPUT121), .A3(new_n1199), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1010), .A2(new_n751), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n990), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT121), .B1(new_n1234), .B2(new_n1199), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1232), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1195), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1205), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n941), .B1(new_n1236), .B2(new_n896), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1231), .B1(new_n1240), .B2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n768), .B1(new_n1245), .B2(new_n1207), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT121), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n751), .B(new_n895), .C1(new_n787), .C2(new_n803), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(new_n941), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n1237), .A3(new_n1235), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1247), .B1(new_n1232), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1197), .A2(new_n1206), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1231), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1229), .B1(new_n1246), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT124), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT124), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1257), .B(new_n1229), .C1(new_n1246), .C2(new_n1254), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(G378));
  NAND2_X1  g1060(.A1(new_n997), .A2(new_n1002), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n751), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n299), .A2(new_n303), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n947), .A2(new_n263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT55), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1263), .B(new_n1265), .ZN(new_n1266));
  XOR2_X1   g1066(.A(KEYINPUT125), .B(KEYINPUT56), .Z(new_n1267));
  XNOR2_X1  g1067(.A(new_n1266), .B(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1261), .A2(new_n1262), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n982), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1010), .A2(new_n1186), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1001), .B1(new_n1272), .B2(new_n1000), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n991), .A2(KEYINPUT109), .A3(new_n996), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1262), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1268), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n969), .A2(new_n981), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1261), .A2(new_n1262), .A3(new_n1268), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1271), .A2(new_n1280), .A3(new_n1158), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n822), .B1(new_n904), .B2(G50), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n390), .A2(G41), .ZN(new_n1283));
  AOI211_X1 g1083(.A(G50), .B(new_n1283), .C1(new_n258), .C2(new_n268), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1110), .A2(G68), .B1(new_n918), .B2(new_n1127), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n1285), .B1(new_n220), .B2(new_n865), .C1(new_n880), .C2(new_n521), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n853), .A2(G116), .B1(G107), .B2(new_n856), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n202), .B2(new_n863), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1283), .B1(new_n875), .B2(new_n864), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1286), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1284), .B1(new_n1290), .B2(KEYINPUT58), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n856), .A2(G128), .B1(G137), .B2(new_n918), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n865), .B2(new_n1219), .ZN(new_n1293));
  INV_X1    g1093(.A(G132), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n880), .A2(new_n1294), .B1(new_n257), .B2(new_n846), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1293), .B(new_n1295), .C1(G125), .C2(new_n853), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(KEYINPUT59), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n876), .A2(G124), .ZN(new_n1299));
  AOI211_X1 g1099(.A(G33), .B(G41), .C1(new_n1170), .C2(G159), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT59), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1299), .B(new_n1300), .C1(new_n1296), .C2(new_n1301), .ZN(new_n1302));
  OAI221_X1 g1102(.A(new_n1291), .B1(KEYINPUT58), .B2(new_n1290), .C1(new_n1298), .C2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1282), .B1(new_n1303), .B2(new_n842), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1276), .B2(new_n828), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1281), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1269), .A2(new_n1270), .A3(new_n982), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1278), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n930), .A2(new_n1230), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT57), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1271), .A2(new_n1280), .A3(KEYINPUT57), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1240), .A2(new_n1244), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1231), .B1(new_n1207), .B2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n768), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1307), .B1(new_n1313), .B2(new_n1317), .ZN(G375));
  NAND2_X1  g1118(.A1(new_n1199), .A2(new_n827), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n822), .B1(new_n905), .B2(G68), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n853), .A2(G294), .B1(G283), .B2(new_n856), .ZN(new_n1321));
  OAI221_X1 g1121(.A(new_n1321), .B1(new_n521), .B2(new_n865), .C1(new_n559), .C2(new_n880), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n285), .B1(G107), .B2(new_n918), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1110), .A2(new_n1127), .B1(new_n1170), .B2(G77), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1323), .B(new_n1324), .C1(new_n866), .C2(new_n875), .ZN(new_n1325));
  AOI22_X1  g1125(.A1(new_n856), .A2(G137), .B1(G159), .B2(new_n921), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1326), .B1(new_n878), .B2(new_n1294), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n876), .A2(G128), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n859), .A2(new_n1218), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n414), .B1(G150), .B2(new_n918), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1110), .A2(G50), .B1(new_n1170), .B2(G58), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1328), .A2(new_n1329), .A3(new_n1330), .A4(new_n1331), .ZN(new_n1332));
  OAI22_X1  g1132(.A1(new_n1322), .A2(new_n1325), .B1(new_n1327), .B2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1320), .B1(new_n1333), .B2(new_n842), .ZN(new_n1334));
  AOI22_X1  g1134(.A1(new_n1315), .A2(new_n1158), .B1(new_n1319), .B2(new_n1334), .ZN(new_n1335));
  OR2_X1    g1135(.A1(new_n1245), .A2(new_n1090), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1315), .A2(new_n1311), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1335), .B1(new_n1336), .B2(new_n1337), .ZN(G381));
  INV_X1    g1138(.A(G387), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1255), .ZN(new_n1340));
  INV_X1    g1140(.A(G396), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1123), .A2(new_n1159), .A3(new_n1341), .ZN(new_n1342));
  NOR4_X1   g1142(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(G375), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1339), .A2(new_n1340), .A3(new_n1343), .A4(new_n1344), .ZN(G407));
  OR3_X1    g1145(.A1(G375), .A2(G343), .A3(new_n1255), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(G407), .A2(G213), .A3(new_n1346), .ZN(G409));
  INV_X1    g1147(.A(new_n1342), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1341), .B1(new_n1123), .B2(new_n1159), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1069), .A2(new_n1077), .A3(new_n1087), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1087), .B1(new_n1069), .B2(new_n1077), .ZN(new_n1352));
  NOR3_X1   g1152(.A1(new_n1351), .A2(new_n1352), .A3(new_n769), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1078), .A2(new_n1158), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1164), .A2(new_n1183), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1350), .B1(new_n1353), .B2(new_n1356), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1163), .B(new_n1184), .C1(new_n1348), .C2(new_n1349), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(G387), .A2(new_n1359), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1092), .A2(new_n1357), .A3(new_n1358), .A4(new_n1119), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1271), .A2(new_n1280), .ZN(new_n1363));
  NOR3_X1   g1163(.A1(new_n1363), .A2(new_n1316), .A3(new_n1090), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1340), .B1(new_n1364), .B2(new_n1306), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1365), .B1(new_n1259), .B2(G375), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT62), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n724), .A2(G343), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n941), .B1(new_n804), .B2(new_n896), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1187), .B1(new_n1370), .B2(KEYINPUT121), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1198), .B1(new_n1371), .B2(new_n1250), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1311), .B1(new_n1372), .B2(new_n1247), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1240), .A2(new_n1231), .A3(new_n1244), .A4(KEYINPUT60), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1373), .A2(new_n1374), .A3(new_n768), .ZN(new_n1375));
  AOI21_X1  g1175(.A(KEYINPUT60), .B1(new_n1252), .B2(new_n1231), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1335), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1377));
  INV_X1    g1177(.A(G384), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  OAI211_X1 g1179(.A(G384), .B(new_n1335), .C1(new_n1375), .C2(new_n1376), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1381), .ZN(new_n1382));
  NAND4_X1  g1182(.A1(new_n1366), .A2(new_n1367), .A3(new_n1369), .A4(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(KEYINPUT61), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1368), .A2(KEYINPUT126), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1379), .A2(new_n1380), .A3(new_n1385), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1368), .A2(G2897), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1386), .A2(new_n1387), .ZN(new_n1388));
  INV_X1    g1188(.A(new_n1387), .ZN(new_n1389));
  NAND4_X1  g1189(.A1(new_n1379), .A2(new_n1380), .A3(new_n1389), .A4(new_n1385), .ZN(new_n1390));
  AND2_X1   g1190(.A1(new_n1388), .A2(new_n1390), .ZN(new_n1391));
  INV_X1    g1191(.A(KEYINPUT57), .ZN(new_n1392));
  OAI21_X1  g1192(.A(new_n1392), .B1(new_n1363), .B2(new_n1316), .ZN(new_n1393));
  NAND4_X1  g1193(.A1(new_n1312), .A2(KEYINPUT57), .A3(new_n1280), .A4(new_n1271), .ZN(new_n1394));
  NAND3_X1  g1194(.A1(new_n1393), .A2(new_n768), .A3(new_n1394), .ZN(new_n1395));
  NAND4_X1  g1195(.A1(new_n1395), .A2(new_n1256), .A3(new_n1258), .A4(new_n1307), .ZN(new_n1396));
  AOI21_X1  g1196(.A(new_n1368), .B1(new_n1396), .B2(new_n1365), .ZN(new_n1397));
  OAI211_X1 g1197(.A(new_n1383), .B(new_n1384), .C1(new_n1391), .C2(new_n1397), .ZN(new_n1398));
  AOI211_X1 g1198(.A(new_n1368), .B(new_n1381), .C1(new_n1396), .C2(new_n1365), .ZN(new_n1399));
  NOR2_X1   g1199(.A1(new_n1399), .A2(new_n1367), .ZN(new_n1400));
  OAI21_X1  g1200(.A(new_n1362), .B1(new_n1398), .B2(new_n1400), .ZN(new_n1401));
  NAND3_X1  g1201(.A1(new_n1360), .A2(new_n1384), .A3(new_n1361), .ZN(new_n1402));
  AOI21_X1  g1202(.A(new_n1402), .B1(new_n1399), .B2(KEYINPUT63), .ZN(new_n1403));
  INV_X1    g1203(.A(KEYINPUT127), .ZN(new_n1404));
  OAI21_X1  g1204(.A(new_n1404), .B1(new_n1391), .B2(new_n1397), .ZN(new_n1405));
  NAND2_X1  g1205(.A1(new_n1366), .A2(new_n1369), .ZN(new_n1406));
  NAND2_X1  g1206(.A1(new_n1388), .A2(new_n1390), .ZN(new_n1407));
  NAND3_X1  g1207(.A1(new_n1406), .A2(KEYINPUT127), .A3(new_n1407), .ZN(new_n1408));
  INV_X1    g1208(.A(KEYINPUT63), .ZN(new_n1409));
  OAI21_X1  g1209(.A(new_n1409), .B1(new_n1406), .B2(new_n1381), .ZN(new_n1410));
  NAND4_X1  g1210(.A1(new_n1403), .A2(new_n1405), .A3(new_n1408), .A4(new_n1410), .ZN(new_n1411));
  NAND2_X1  g1211(.A1(new_n1401), .A2(new_n1411), .ZN(G405));
  NAND2_X1  g1212(.A1(G375), .A2(new_n1340), .ZN(new_n1413));
  NAND2_X1  g1213(.A1(new_n1413), .A2(new_n1396), .ZN(new_n1414));
  XNOR2_X1  g1214(.A(new_n1414), .B(new_n1382), .ZN(new_n1415));
  XNOR2_X1  g1215(.A(new_n1415), .B(new_n1362), .ZN(G402));
endmodule


