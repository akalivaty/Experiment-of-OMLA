

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580;

  OR2_X2 U324 ( .A1(n381), .A2(n563), .ZN(n383) );
  XNOR2_X1 U325 ( .A(n426), .B(n425), .ZN(n567) );
  INV_X1 U326 ( .A(KEYINPUT65), .ZN(n425) );
  XNOR2_X1 U327 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U328 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U329 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n317) );
  XNOR2_X1 U330 ( .A(n429), .B(n317), .ZN(n318) );
  XNOR2_X1 U331 ( .A(n357), .B(n356), .ZN(n358) );
  INV_X1 U332 ( .A(n567), .ZN(n445) );
  XNOR2_X1 U333 ( .A(n360), .B(n326), .ZN(n327) );
  XNOR2_X1 U334 ( .A(n328), .B(n327), .ZN(n384) );
  XNOR2_X1 U335 ( .A(n365), .B(n364), .ZN(n558) );
  XNOR2_X1 U336 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U337 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n293) );
  XNOR2_X1 U339 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U341 ( .A(KEYINPUT19), .B(n294), .Z(n399) );
  XOR2_X1 U342 ( .A(KEYINPUT20), .B(G183GAT), .Z(n296) );
  XNOR2_X1 U343 ( .A(G15GAT), .B(G71GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U345 ( .A(KEYINPUT66), .B(KEYINPUT80), .Z(n298) );
  XNOR2_X1 U346 ( .A(KEYINPUT81), .B(KEYINPUT83), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U348 ( .A(n300), .B(n299), .Z(n313) );
  XOR2_X1 U349 ( .A(KEYINPUT0), .B(KEYINPUT78), .Z(n302) );
  XNOR2_X1 U350 ( .A(G134GAT), .B(G120GAT), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U352 ( .A(n303), .B(G127GAT), .Z(n305) );
  XNOR2_X1 U353 ( .A(G113GAT), .B(KEYINPUT79), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n411) );
  XOR2_X1 U355 ( .A(G176GAT), .B(G190GAT), .Z(n307) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G99GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U358 ( .A(KEYINPUT84), .B(n308), .Z(n310) );
  NAND2_X1 U359 ( .A1(G227GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n411), .B(n311), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n399), .B(n314), .ZN(n533) );
  XOR2_X1 U364 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n316) );
  XNOR2_X1 U365 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n315) );
  XOR2_X1 U366 ( .A(n316), .B(n315), .Z(n319) );
  XOR2_X1 U367 ( .A(G148GAT), .B(G106GAT), .Z(n429) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n325) );
  XOR2_X1 U369 ( .A(G64GAT), .B(G204GAT), .Z(n321) );
  XNOR2_X1 U370 ( .A(G176GAT), .B(G92GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n396) );
  XOR2_X1 U372 ( .A(G78GAT), .B(KEYINPUT13), .Z(n323) );
  XNOR2_X1 U373 ( .A(G71GAT), .B(G57GAT), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n373) );
  XOR2_X1 U375 ( .A(n396), .B(n373), .Z(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n328) );
  XOR2_X1 U377 ( .A(G99GAT), .B(G85GAT), .Z(n360) );
  NAND2_X1 U378 ( .A1(G230GAT), .A2(G233GAT), .ZN(n326) );
  XOR2_X1 U379 ( .A(n384), .B(KEYINPUT64), .Z(n329) );
  XNOR2_X1 U380 ( .A(KEYINPUT41), .B(n329), .ZN(n550) );
  XNOR2_X1 U381 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n330), .B(G15GAT), .ZN(n369) );
  XOR2_X1 U383 ( .A(G36GAT), .B(n369), .Z(n332) );
  NAND2_X1 U384 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U386 ( .A(n333), .B(G50GAT), .Z(n341) );
  XOR2_X1 U387 ( .A(G141GAT), .B(G197GAT), .Z(n335) );
  XNOR2_X1 U388 ( .A(G169GAT), .B(G22GAT), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U390 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n337) );
  XNOR2_X1 U391 ( .A(G113GAT), .B(KEYINPUT29), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U395 ( .A(n342), .B(G8GAT), .Z(n346) );
  XOR2_X1 U396 ( .A(G29GAT), .B(G43GAT), .Z(n344) );
  XNOR2_X1 U397 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n355) );
  XNOR2_X1 U399 ( .A(n355), .B(KEYINPUT68), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n568) );
  NAND2_X1 U401 ( .A1(n550), .A2(n568), .ZN(n349) );
  XOR2_X1 U402 ( .A(KEYINPUT46), .B(KEYINPUT110), .Z(n347) );
  XNOR2_X1 U403 ( .A(KEYINPUT109), .B(n347), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n366) );
  XOR2_X1 U405 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n351) );
  XNOR2_X1 U406 ( .A(G134GAT), .B(KEYINPUT74), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n365) );
  XNOR2_X1 U408 ( .A(G36GAT), .B(G190GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n352), .B(G218GAT), .ZN(n398) );
  XOR2_X1 U410 ( .A(G50GAT), .B(G162GAT), .Z(n440) );
  XNOR2_X1 U411 ( .A(n398), .B(n440), .ZN(n354) );
  AND2_X1 U412 ( .A1(G232GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n355), .B(G106GAT), .ZN(n357) );
  INV_X1 U415 ( .A(G92GAT), .ZN(n356) );
  XOR2_X1 U416 ( .A(n361), .B(n360), .Z(n363) );
  XNOR2_X1 U417 ( .A(KEYINPUT73), .B(KEYINPUT10), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n364) );
  INV_X1 U419 ( .A(n558), .ZN(n457) );
  NAND2_X1 U420 ( .A1(n366), .A2(n457), .ZN(n381) );
  XOR2_X1 U421 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n368) );
  XNOR2_X1 U422 ( .A(G127GAT), .B(KEYINPUT15), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n380) );
  XOR2_X1 U424 ( .A(G8GAT), .B(G183GAT), .Z(n393) );
  XOR2_X1 U425 ( .A(n369), .B(n393), .Z(n371) );
  NAND2_X1 U426 ( .A1(G231GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U428 ( .A(n372), .B(KEYINPUT12), .Z(n375) );
  XNOR2_X1 U429 ( .A(n373), .B(KEYINPUT14), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U431 ( .A(G22GAT), .B(G155GAT), .Z(n430) );
  XOR2_X1 U432 ( .A(n376), .B(n430), .Z(n378) );
  XNOR2_X1 U433 ( .A(G64GAT), .B(G211GAT), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n489) );
  XNOR2_X1 U436 ( .A(KEYINPUT108), .B(n489), .ZN(n563) );
  XOR2_X1 U437 ( .A(KEYINPUT47), .B(KEYINPUT111), .Z(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n390) );
  XNOR2_X1 U439 ( .A(KEYINPUT36), .B(n558), .ZN(n577) );
  NAND2_X1 U440 ( .A1(n577), .A2(n489), .ZN(n386) );
  XOR2_X1 U441 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n385) );
  INV_X1 U442 ( .A(n568), .ZN(n507) );
  NAND2_X1 U443 ( .A1(n387), .A2(n507), .ZN(n388) );
  NOR2_X1 U444 ( .A1(n384), .A2(n388), .ZN(n389) );
  NOR2_X1 U445 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U446 ( .A(KEYINPUT48), .B(n391), .ZN(n530) );
  XNOR2_X1 U447 ( .A(G197GAT), .B(G211GAT), .ZN(n392) );
  XOR2_X1 U448 ( .A(n392), .B(KEYINPUT21), .Z(n427) );
  XNOR2_X1 U449 ( .A(n427), .B(n393), .ZN(n395) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n397) );
  XOR2_X1 U452 ( .A(n397), .B(n396), .Z(n401) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U454 ( .A(n401), .B(n400), .Z(n522) );
  XOR2_X1 U455 ( .A(n522), .B(KEYINPUT121), .Z(n402) );
  NOR2_X1 U456 ( .A1(n530), .A2(n402), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n403), .B(KEYINPUT54), .ZN(n424) );
  NAND2_X1 U458 ( .A1(G225GAT), .A2(G233GAT), .ZN(n409) );
  XOR2_X1 U459 ( .A(G57GAT), .B(G148GAT), .Z(n405) );
  XNOR2_X1 U460 ( .A(G29GAT), .B(G1GAT), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U462 ( .A(G162GAT), .B(G85GAT), .Z(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n423) );
  XOR2_X1 U466 ( .A(KEYINPUT89), .B(KEYINPUT87), .Z(n413) );
  XNOR2_X1 U467 ( .A(KEYINPUT5), .B(KEYINPUT91), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U469 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n415) );
  XNOR2_X1 U470 ( .A(G155GAT), .B(KEYINPUT1), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n421) );
  XNOR2_X1 U473 ( .A(KEYINPUT88), .B(KEYINPUT90), .ZN(n419) );
  XOR2_X1 U474 ( .A(G141GAT), .B(KEYINPUT3), .Z(n418) );
  XOR2_X1 U475 ( .A(KEYINPUT2), .B(n418), .Z(n428) );
  XOR2_X1 U476 ( .A(n419), .B(n428), .Z(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n520) );
  NAND2_X1 U479 ( .A1(n424), .A2(n520), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n444) );
  XOR2_X1 U481 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U483 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U484 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n434) );
  XNOR2_X1 U485 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U487 ( .A(n436), .B(n435), .Z(n442) );
  XOR2_X1 U488 ( .A(KEYINPUT24), .B(G78GAT), .Z(n438) );
  XNOR2_X1 U489 ( .A(G218GAT), .B(G204GAT), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U492 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U493 ( .A(n444), .B(n443), .ZN(n470) );
  NAND2_X1 U494 ( .A1(n445), .A2(n470), .ZN(n447) );
  INV_X1 U495 ( .A(KEYINPUT55), .ZN(n446) );
  XNOR2_X1 U496 ( .A(n447), .B(n446), .ZN(n448) );
  NOR2_X1 U497 ( .A1(n533), .A2(n448), .ZN(n564) );
  NAND2_X1 U498 ( .A1(n564), .A2(n558), .ZN(n452) );
  XOR2_X1 U499 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n450) );
  XNOR2_X1 U500 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n449) );
  NAND2_X1 U501 ( .A1(n564), .A2(n550), .ZN(n456) );
  XOR2_X1 U502 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n454) );
  XOR2_X1 U503 ( .A(G176GAT), .B(KEYINPUT56), .Z(n453) );
  XNOR2_X1 U504 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U505 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  NOR2_X1 U506 ( .A1(n384), .A2(n507), .ZN(n494) );
  NAND2_X1 U507 ( .A1(n489), .A2(n457), .ZN(n458) );
  XNOR2_X1 U508 ( .A(n458), .B(KEYINPUT16), .ZN(n459) );
  XNOR2_X1 U509 ( .A(n459), .B(KEYINPUT77), .ZN(n477) );
  XNOR2_X1 U510 ( .A(n522), .B(KEYINPUT92), .ZN(n460) );
  XNOR2_X1 U511 ( .A(KEYINPUT27), .B(n460), .ZN(n472) );
  INV_X1 U512 ( .A(n533), .ZN(n461) );
  NOR2_X1 U513 ( .A1(n461), .A2(n470), .ZN(n463) );
  XNOR2_X1 U514 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n462) );
  XOR2_X1 U515 ( .A(n463), .B(n462), .Z(n566) );
  NOR2_X1 U516 ( .A1(n472), .A2(n566), .ZN(n464) );
  XNOR2_X1 U517 ( .A(KEYINPUT95), .B(n464), .ZN(n468) );
  OR2_X1 U518 ( .A1(n533), .A2(n522), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n470), .A2(n465), .ZN(n466) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n466), .Z(n467) );
  NAND2_X1 U521 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U522 ( .A1(n520), .A2(n469), .ZN(n476) );
  XNOR2_X1 U523 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n471) );
  XNOR2_X1 U524 ( .A(n471), .B(n470), .ZN(n536) );
  NOR2_X1 U525 ( .A1(n472), .A2(n520), .ZN(n473) );
  XNOR2_X1 U526 ( .A(n473), .B(KEYINPUT93), .ZN(n531) );
  NOR2_X1 U527 ( .A1(n536), .A2(n531), .ZN(n474) );
  NAND2_X1 U528 ( .A1(n474), .A2(n533), .ZN(n475) );
  NAND2_X1 U529 ( .A1(n476), .A2(n475), .ZN(n490) );
  NAND2_X1 U530 ( .A1(n477), .A2(n490), .ZN(n478) );
  XOR2_X1 U531 ( .A(KEYINPUT96), .B(n478), .Z(n508) );
  NAND2_X1 U532 ( .A1(n494), .A2(n508), .ZN(n486) );
  NOR2_X1 U533 ( .A1(n520), .A2(n486), .ZN(n480) );
  XNOR2_X1 U534 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NOR2_X1 U537 ( .A1(n522), .A2(n486), .ZN(n482) );
  XOR2_X1 U538 ( .A(G8GAT), .B(n482), .Z(G1325GAT) );
  NOR2_X1 U539 ( .A1(n533), .A2(n486), .ZN(n484) );
  XNOR2_X1 U540 ( .A(KEYINPUT35), .B(KEYINPUT98), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  INV_X1 U543 ( .A(n536), .ZN(n526) );
  NOR2_X1 U544 ( .A1(n526), .A2(n486), .ZN(n488) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(G1327GAT) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n497) );
  NAND2_X1 U548 ( .A1(n577), .A2(n490), .ZN(n491) );
  NOR2_X1 U549 ( .A1(n489), .A2(n491), .ZN(n493) );
  XOR2_X1 U550 ( .A(KEYINPUT37), .B(KEYINPUT100), .Z(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n518) );
  NAND2_X1 U552 ( .A1(n518), .A2(n494), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(KEYINPUT38), .ZN(n502) );
  NOR2_X1 U554 ( .A1(n520), .A2(n502), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n502), .A2(n522), .ZN(n498) );
  XOR2_X1 U557 ( .A(G36GAT), .B(n498), .Z(G1329GAT) );
  NOR2_X1 U558 ( .A1(n502), .A2(n533), .ZN(n500) );
  XNOR2_X1 U559 ( .A(KEYINPUT40), .B(KEYINPUT101), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NOR2_X1 U562 ( .A1(n526), .A2(n502), .ZN(n503) );
  XOR2_X1 U563 ( .A(G50GAT), .B(n503), .Z(n504) );
  XNOR2_X1 U564 ( .A(KEYINPUT102), .B(n504), .ZN(G1331GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT104), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(n510) );
  AND2_X1 U568 ( .A1(n507), .A2(n550), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n517), .A2(n508), .ZN(n514) );
  NOR2_X1 U570 ( .A1(n520), .A2(n514), .ZN(n509) );
  XOR2_X1 U571 ( .A(n510), .B(n509), .Z(G1332GAT) );
  NOR2_X1 U572 ( .A1(n522), .A2(n514), .ZN(n511) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n533), .A2(n514), .ZN(n513) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(G1334GAT) );
  NOR2_X1 U577 ( .A1(n526), .A2(n514), .ZN(n516) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n519), .B(KEYINPUT106), .ZN(n525) );
  NOR2_X1 U582 ( .A1(n520), .A2(n525), .ZN(n521) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n521), .Z(G1336GAT) );
  NOR2_X1 U584 ( .A1(n525), .A2(n522), .ZN(n523) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n525), .A2(n533), .ZN(n524) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  XNOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT107), .ZN(n528) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NOR2_X1 U592 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U593 ( .A(n532), .B(KEYINPUT113), .ZN(n548) );
  NOR2_X1 U594 ( .A1(n533), .A2(n548), .ZN(n534) );
  XOR2_X1 U595 ( .A(KEYINPUT114), .B(n534), .Z(n535) );
  NOR2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n568), .A2(n545), .ZN(n537) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n539) );
  NAND2_X1 U600 ( .A1(n545), .A2(n550), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT115), .Z(n540) );
  XNOR2_X1 U603 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n543) );
  NAND2_X1 U605 ( .A1(n545), .A2(n563), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U609 ( .A1(n545), .A2(n558), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U611 ( .A1(n548), .A2(n566), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n568), .A2(n557), .ZN(n549) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U615 ( .A1(n557), .A2(n550), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n555) );
  NAND2_X1 U619 ( .A1(n557), .A2(n489), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n556), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n559), .B(KEYINPUT120), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n568), .A2(n564), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n578) );
  AND2_X1 U631 ( .A1(n568), .A2(n578), .ZN(n570) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U633 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U636 ( .A1(n578), .A2(n384), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n575) );
  NAND2_X1 U639 ( .A1(n578), .A2(n489), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

