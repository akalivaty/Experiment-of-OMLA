

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U554 ( .A1(n523), .A2(G2104), .ZN(n892) );
  INV_X1 U555 ( .A(n764), .ZN(n748) );
  AND2_X1 U556 ( .A1(n747), .A2(n921), .ZN(n520) );
  OR2_X1 U557 ( .A1(n711), .A2(n926), .ZN(n521) );
  XNOR2_X1 U558 ( .A(KEYINPUT87), .B(n795), .ZN(n522) );
  INV_X2 U559 ( .A(n717), .ZN(n711) );
  INV_X1 U560 ( .A(KEYINPUT88), .ZN(n718) );
  XNOR2_X1 U561 ( .A(n737), .B(KEYINPUT32), .ZN(n744) );
  NAND2_X1 U562 ( .A1(n744), .A2(n743), .ZN(n760) );
  XNOR2_X1 U563 ( .A(KEYINPUT12), .B(KEYINPUT70), .ZN(n564) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n770) );
  XNOR2_X1 U565 ( .A(n565), .B(n564), .ZN(n567) );
  NAND2_X1 U566 ( .A1(n522), .A2(n796), .ZN(n797) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n654) );
  OR2_X1 U568 ( .A1(n798), .A2(n797), .ZN(n813) );
  NAND2_X1 U569 ( .A1(n894), .A2(G137), .ZN(n531) );
  NOR2_X1 U570 ( .A1(n570), .A2(n569), .ZN(n935) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n887) );
  NAND2_X1 U572 ( .A1(n887), .A2(G113), .ZN(n526) );
  INV_X1 U573 ( .A(G2105), .ZN(n523) );
  NAND2_X1 U574 ( .A1(G101), .A2(n892), .ZN(n524) );
  XOR2_X1 U575 ( .A(KEYINPUT23), .B(n524), .Z(n525) );
  NAND2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n533) );
  XNOR2_X1 U577 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n528) );
  NOR2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XNOR2_X2 U579 ( .A(n528), .B(n527), .ZN(n894) );
  NOR2_X1 U580 ( .A1(n523), .A2(G2104), .ZN(n529) );
  XNOR2_X2 U581 ( .A(n529), .B(KEYINPUT64), .ZN(n888) );
  NAND2_X1 U582 ( .A1(G125), .A2(n888), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U584 ( .A1(n533), .A2(n532), .ZN(G160) );
  NAND2_X1 U585 ( .A1(G102), .A2(n892), .ZN(n535) );
  NAND2_X1 U586 ( .A1(G138), .A2(n894), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U588 ( .A1(G114), .A2(n887), .ZN(n537) );
  NAND2_X1 U589 ( .A1(G126), .A2(n888), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U591 ( .A1(n539), .A2(n538), .ZN(G164) );
  INV_X1 U592 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U593 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U594 ( .A(G82), .ZN(G220) );
  INV_X1 U595 ( .A(G132), .ZN(G219) );
  NAND2_X1 U596 ( .A1(G69), .A2(G120), .ZN(n540) );
  NOR2_X1 U597 ( .A1(G237), .A2(n540), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G108), .A2(n541), .ZN(n833) );
  NAND2_X1 U599 ( .A1(n833), .A2(G567), .ZN(n546) );
  NOR2_X1 U600 ( .A1(G220), .A2(G219), .ZN(n542) );
  XOR2_X1 U601 ( .A(KEYINPUT22), .B(n542), .Z(n543) );
  NOR2_X1 U602 ( .A1(G218), .A2(n543), .ZN(n544) );
  NAND2_X1 U603 ( .A1(G96), .A2(n544), .ZN(n834) );
  NAND2_X1 U604 ( .A1(n834), .A2(G2106), .ZN(n545) );
  AND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(G319) );
  INV_X1 U606 ( .A(G651), .ZN(n549) );
  NOR2_X1 U607 ( .A1(G543), .A2(n549), .ZN(n547) );
  XOR2_X1 U608 ( .A(KEYINPUT1), .B(n547), .Z(n650) );
  NAND2_X1 U609 ( .A1(G64), .A2(n650), .ZN(n548) );
  XNOR2_X1 U610 ( .A(n548), .B(KEYINPUT67), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G90), .A2(n654), .ZN(n551) );
  XOR2_X1 U612 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  NOR2_X1 U613 ( .A1(n623), .A2(n549), .ZN(n655) );
  NAND2_X1 U614 ( .A1(G77), .A2(n655), .ZN(n550) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n552), .B(KEYINPUT9), .ZN(n554) );
  NOR2_X2 U617 ( .A1(G651), .A2(n623), .ZN(n651) );
  NAND2_X1 U618 ( .A1(G52), .A2(n651), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U620 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U621 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U622 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n558) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G223) );
  INV_X1 U625 ( .A(G223), .ZN(n826) );
  NAND2_X1 U626 ( .A1(n826), .A2(G567), .ZN(n559) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n559), .Z(G234) );
  NAND2_X1 U628 ( .A1(G56), .A2(n650), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n560), .B(KEYINPUT14), .ZN(n563) );
  NAND2_X1 U630 ( .A1(G43), .A2(n651), .ZN(n561) );
  XOR2_X1 U631 ( .A(KEYINPUT71), .B(n561), .Z(n562) );
  NAND2_X1 U632 ( .A1(n563), .A2(n562), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G81), .A2(n654), .ZN(n565) );
  NAND2_X1 U634 ( .A1(G68), .A2(n655), .ZN(n566) );
  NAND2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U636 ( .A(KEYINPUT13), .B(n568), .Z(n569) );
  NAND2_X1 U637 ( .A1(n935), .A2(G860), .ZN(G153) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G92), .A2(n654), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n571), .B(KEYINPUT72), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G66), .A2(n650), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G79), .A2(n655), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G54), .A2(n651), .ZN(n574) );
  XNOR2_X1 U646 ( .A(KEYINPUT73), .B(n574), .ZN(n575) );
  NOR2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U649 ( .A(KEYINPUT15), .B(n579), .ZN(n927) );
  OR2_X1 U650 ( .A1(n927), .A2(G868), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U652 ( .A1(n654), .A2(G89), .ZN(n582) );
  XNOR2_X1 U653 ( .A(n582), .B(KEYINPUT4), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G76), .A2(n655), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U656 ( .A(n585), .B(KEYINPUT5), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G63), .A2(n650), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G51), .A2(n651), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U660 ( .A(KEYINPUT6), .B(n588), .Z(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U662 ( .A(n591), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U663 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U664 ( .A1(G65), .A2(n650), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G53), .A2(n651), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n654), .A2(G91), .ZN(n594) );
  XOR2_X1 U668 ( .A(KEYINPUT68), .B(n594), .Z(n595) );
  NOR2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n655), .A2(G78), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(G299) );
  INV_X1 U672 ( .A(G868), .ZN(n666) );
  NOR2_X1 U673 ( .A1(G286), .A2(n666), .ZN(n600) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n600), .A2(n599), .ZN(G297) );
  INV_X1 U676 ( .A(G860), .ZN(n836) );
  NAND2_X1 U677 ( .A1(n836), .A2(G559), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n601), .A2(n927), .ZN(n602) );
  XNOR2_X1 U679 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G559), .A2(n666), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n927), .A2(n603), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n935), .A2(n666), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U684 ( .A(KEYINPUT74), .B(n606), .Z(G282) );
  NAND2_X1 U685 ( .A1(G99), .A2(n892), .ZN(n608) );
  NAND2_X1 U686 ( .A1(G111), .A2(n887), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n888), .A2(G123), .ZN(n609) );
  XNOR2_X1 U689 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n894), .A2(G135), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n995) );
  XNOR2_X1 U693 ( .A(G2096), .B(n995), .ZN(n615) );
  INV_X1 U694 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G88), .A2(n654), .ZN(n617) );
  NAND2_X1 U697 ( .A1(G75), .A2(n655), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G62), .A2(n650), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G50), .A2(n651), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U702 ( .A1(n621), .A2(n620), .ZN(G166) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n622) );
  XNOR2_X1 U704 ( .A(n622), .B(KEYINPUT78), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G49), .A2(n651), .ZN(n625) );
  NAND2_X1 U706 ( .A1(G87), .A2(n623), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U708 ( .A1(n650), .A2(n626), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G60), .A2(n650), .ZN(n630) );
  NAND2_X1 U711 ( .A1(G47), .A2(n651), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U713 ( .A(KEYINPUT66), .B(n631), .Z(n635) );
  NAND2_X1 U714 ( .A1(G85), .A2(n654), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G72), .A2(n655), .ZN(n632) );
  AND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(G290) );
  XOR2_X1 U718 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n637) );
  NAND2_X1 U719 ( .A1(G73), .A2(n655), .ZN(n636) );
  XNOR2_X1 U720 ( .A(n637), .B(n636), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G61), .A2(n650), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G86), .A2(n654), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U724 ( .A(KEYINPUT79), .B(n640), .Z(n641) );
  NOR2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n651), .A2(G48), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(G305) );
  XOR2_X1 U728 ( .A(n935), .B(KEYINPUT75), .Z(n646) );
  NAND2_X1 U729 ( .A1(G559), .A2(n927), .ZN(n645) );
  XNOR2_X1 U730 ( .A(n646), .B(n645), .ZN(n835) );
  XOR2_X1 U731 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n648) );
  INV_X1 U732 ( .A(G299), .ZN(n918) );
  XNOR2_X1 U733 ( .A(n918), .B(G166), .ZN(n647) );
  XNOR2_X1 U734 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U735 ( .A(n649), .B(G288), .ZN(n662) );
  NAND2_X1 U736 ( .A1(G67), .A2(n650), .ZN(n653) );
  NAND2_X1 U737 ( .A1(G55), .A2(n651), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n653), .A2(n652), .ZN(n660) );
  NAND2_X1 U739 ( .A1(G93), .A2(n654), .ZN(n657) );
  NAND2_X1 U740 ( .A1(G80), .A2(n655), .ZN(n656) );
  NAND2_X1 U741 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U742 ( .A(KEYINPUT76), .B(n658), .ZN(n659) );
  NOR2_X1 U743 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n661), .B(KEYINPUT77), .ZN(n837) );
  XNOR2_X1 U745 ( .A(n662), .B(n837), .ZN(n663) );
  XNOR2_X1 U746 ( .A(n663), .B(G290), .ZN(n664) );
  XNOR2_X1 U747 ( .A(n664), .B(G305), .ZN(n906) );
  XNOR2_X1 U748 ( .A(n835), .B(n906), .ZN(n665) );
  NAND2_X1 U749 ( .A1(n665), .A2(G868), .ZN(n668) );
  NAND2_X1 U750 ( .A1(n837), .A2(n666), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U754 ( .A1(n670), .A2(G2090), .ZN(n671) );
  XNOR2_X1 U755 ( .A(n671), .B(KEYINPUT21), .ZN(n672) );
  XNOR2_X1 U756 ( .A(KEYINPUT82), .B(n672), .ZN(n673) );
  NAND2_X1 U757 ( .A1(G2072), .A2(n673), .ZN(G158) );
  NAND2_X1 U758 ( .A1(G661), .A2(G483), .ZN(n674) );
  XNOR2_X1 U759 ( .A(KEYINPUT83), .B(n674), .ZN(n675) );
  NAND2_X1 U760 ( .A1(n675), .A2(G319), .ZN(n676) );
  XOR2_X1 U761 ( .A(KEYINPUT84), .B(n676), .Z(n832) );
  NAND2_X1 U762 ( .A1(G36), .A2(n832), .ZN(G176) );
  XNOR2_X1 U763 ( .A(KEYINPUT85), .B(G166), .ZN(G303) );
  NAND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n769) );
  INV_X1 U765 ( .A(n769), .ZN(n677) );
  NAND2_X2 U766 ( .A1(n677), .A2(n770), .ZN(n717) );
  NAND2_X1 U767 ( .A1(G1996), .A2(n711), .ZN(n678) );
  XNOR2_X1 U768 ( .A(n678), .B(KEYINPUT26), .ZN(n679) );
  NAND2_X1 U769 ( .A1(n717), .A2(G1341), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n679), .A2(n682), .ZN(n680) );
  NAND2_X1 U771 ( .A1(n680), .A2(KEYINPUT92), .ZN(n681) );
  NAND2_X1 U772 ( .A1(n935), .A2(n681), .ZN(n686) );
  INV_X1 U773 ( .A(KEYINPUT26), .ZN(n683) );
  NOR2_X1 U774 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U775 ( .A1(KEYINPUT92), .A2(n684), .ZN(n685) );
  NOR2_X2 U776 ( .A1(n686), .A2(n685), .ZN(n688) );
  NOR2_X1 U777 ( .A1(n688), .A2(n927), .ZN(n687) );
  XNOR2_X1 U778 ( .A(n687), .B(KEYINPUT95), .ZN(n698) );
  NAND2_X1 U779 ( .A1(n688), .A2(n927), .ZN(n696) );
  NAND2_X1 U780 ( .A1(G2067), .A2(n711), .ZN(n689) );
  XNOR2_X1 U781 ( .A(KEYINPUT94), .B(n689), .ZN(n690) );
  INV_X1 U782 ( .A(G1348), .ZN(n926) );
  NAND2_X1 U783 ( .A1(n690), .A2(n521), .ZN(n691) );
  NOR2_X1 U784 ( .A1(KEYINPUT93), .A2(n691), .ZN(n694) );
  NAND2_X1 U785 ( .A1(KEYINPUT94), .A2(KEYINPUT93), .ZN(n692) );
  NOR2_X1 U786 ( .A1(n692), .A2(n521), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n704) );
  NAND2_X1 U790 ( .A1(n717), .A2(G1956), .ZN(n701) );
  NAND2_X1 U791 ( .A1(n711), .A2(G2072), .ZN(n699) );
  XOR2_X1 U792 ( .A(KEYINPUT27), .B(n699), .Z(n700) );
  NAND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U794 ( .A(n702), .B(KEYINPUT91), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n918), .A2(n705), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U797 ( .A1(n918), .A2(n705), .ZN(n706) );
  XOR2_X1 U798 ( .A(n706), .B(KEYINPUT28), .Z(n707) );
  NAND2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U800 ( .A(n709), .B(KEYINPUT29), .ZN(n716) );
  XNOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .ZN(n971) );
  NAND2_X1 U802 ( .A1(n711), .A2(n971), .ZN(n710) );
  XNOR2_X1 U803 ( .A(n710), .B(KEYINPUT89), .ZN(n713) );
  NOR2_X1 U804 ( .A1(n711), .A2(G1961), .ZN(n712) );
  NOR2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U806 ( .A(KEYINPUT90), .B(n714), .Z(n724) );
  AND2_X1 U807 ( .A1(G171), .A2(n724), .ZN(n715) );
  NOR2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n729) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n717), .ZN(n738) );
  NAND2_X1 U810 ( .A1(G8), .A2(n717), .ZN(n764) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n764), .ZN(n719) );
  XNOR2_X1 U812 ( .A(n719), .B(n718), .ZN(n739) );
  NAND2_X1 U813 ( .A1(n739), .A2(G8), .ZN(n720) );
  NOR2_X1 U814 ( .A1(n738), .A2(n720), .ZN(n722) );
  XOR2_X1 U815 ( .A(KEYINPUT96), .B(KEYINPUT30), .Z(n721) );
  XNOR2_X1 U816 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U817 ( .A1(G168), .A2(n723), .ZN(n726) );
  NOR2_X1 U818 ( .A1(G171), .A2(n724), .ZN(n725) );
  NOR2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U820 ( .A(n727), .B(KEYINPUT31), .ZN(n728) );
  NOR2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U822 ( .A(n730), .B(KEYINPUT97), .ZN(n740) );
  NAND2_X1 U823 ( .A1(n740), .A2(G286), .ZN(n735) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n764), .ZN(n732) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n717), .ZN(n731) );
  NOR2_X1 U826 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U827 ( .A1(n733), .A2(G303), .ZN(n734) );
  NAND2_X1 U828 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n736), .A2(G8), .ZN(n737) );
  NAND2_X1 U830 ( .A1(G8), .A2(n738), .ZN(n742) );
  AND2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n745) );
  NOR2_X1 U835 ( .A1(n751), .A2(n745), .ZN(n924) );
  XNOR2_X1 U836 ( .A(KEYINPUT98), .B(n924), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n760), .A2(n746), .ZN(n747) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n921) );
  NAND2_X1 U839 ( .A1(n520), .A2(n748), .ZN(n750) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n749) );
  NAND2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U843 ( .A1(n752), .A2(n764), .ZN(n754) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n938) );
  INV_X1 U845 ( .A(n938), .ZN(n753) );
  NOR2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U848 ( .A(KEYINPUT99), .B(n757), .ZN(n768) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U850 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n764), .A2(n761), .ZN(n766) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U854 ( .A(n762), .B(KEYINPUT24), .Z(n763) );
  OR2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n798) );
  NOR2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n810) );
  NAND2_X1 U859 ( .A1(G104), .A2(n892), .ZN(n772) );
  NAND2_X1 U860 ( .A1(G140), .A2(n894), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U862 ( .A(KEYINPUT34), .B(n773), .ZN(n778) );
  NAND2_X1 U863 ( .A1(G116), .A2(n887), .ZN(n775) );
  NAND2_X1 U864 ( .A1(G128), .A2(n888), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U866 ( .A(KEYINPUT35), .B(n776), .Z(n777) );
  NOR2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U868 ( .A(KEYINPUT36), .B(n779), .ZN(n903) );
  XNOR2_X1 U869 ( .A(KEYINPUT37), .B(G2067), .ZN(n808) );
  NOR2_X1 U870 ( .A1(n903), .A2(n808), .ZN(n1015) );
  NAND2_X1 U871 ( .A1(n810), .A2(n1015), .ZN(n806) );
  NAND2_X1 U872 ( .A1(n888), .A2(G129), .ZN(n780) );
  XNOR2_X1 U873 ( .A(n780), .B(KEYINPUT86), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G141), .A2(n894), .ZN(n782) );
  NAND2_X1 U875 ( .A1(G117), .A2(n887), .ZN(n781) );
  NAND2_X1 U876 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n892), .A2(G105), .ZN(n783) );
  XOR2_X1 U878 ( .A(KEYINPUT38), .B(n783), .Z(n784) );
  NOR2_X1 U879 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n872) );
  AND2_X1 U881 ( .A1(n872), .A2(G1996), .ZN(n998) );
  NAND2_X1 U882 ( .A1(G95), .A2(n892), .ZN(n789) );
  NAND2_X1 U883 ( .A1(G107), .A2(n887), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U885 ( .A1(G131), .A2(n894), .ZN(n791) );
  NAND2_X1 U886 ( .A1(G119), .A2(n888), .ZN(n790) );
  NAND2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n868) );
  INV_X1 U889 ( .A(G1991), .ZN(n800) );
  NOR2_X1 U890 ( .A1(n868), .A2(n800), .ZN(n996) );
  OR2_X1 U891 ( .A1(n998), .A2(n996), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n810), .A2(n794), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n806), .A2(n799), .ZN(n795) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n933) );
  NAND2_X1 U895 ( .A1(n933), .A2(n810), .ZN(n796) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n872), .ZN(n992) );
  INV_X1 U897 ( .A(n799), .ZN(n803) );
  AND2_X1 U898 ( .A1(n800), .A2(n868), .ZN(n997) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U900 ( .A1(n997), .A2(n801), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U902 ( .A1(n992), .A2(n804), .ZN(n805) );
  XNOR2_X1 U903 ( .A(n805), .B(KEYINPUT39), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n903), .A2(n808), .ZN(n1004) );
  NAND2_X1 U906 ( .A1(n809), .A2(n1004), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n815) );
  XNOR2_X1 U909 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n814) );
  XNOR2_X1 U910 ( .A(n815), .B(n814), .ZN(G329) );
  XOR2_X1 U911 ( .A(G2430), .B(G2451), .Z(n817) );
  XNOR2_X1 U912 ( .A(G2446), .B(G2427), .ZN(n816) );
  XNOR2_X1 U913 ( .A(n817), .B(n816), .ZN(n824) );
  XOR2_X1 U914 ( .A(G2438), .B(KEYINPUT101), .Z(n819) );
  XNOR2_X1 U915 ( .A(G2443), .B(G2454), .ZN(n818) );
  XNOR2_X1 U916 ( .A(n819), .B(n818), .ZN(n820) );
  XOR2_X1 U917 ( .A(n820), .B(G2435), .Z(n822) );
  XNOR2_X1 U918 ( .A(G1348), .B(G1341), .ZN(n821) );
  XNOR2_X1 U919 ( .A(n822), .B(n821), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n824), .B(n823), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n825), .A2(G14), .ZN(n912) );
  XOR2_X1 U922 ( .A(KEYINPUT102), .B(n912), .Z(G401) );
  NAND2_X1 U923 ( .A1(n826), .A2(G2106), .ZN(n827) );
  XOR2_X1 U924 ( .A(KEYINPUT103), .B(n827), .Z(G217) );
  INV_X1 U925 ( .A(G661), .ZN(n829) );
  NAND2_X1 U926 ( .A1(G2), .A2(G15), .ZN(n828) );
  NOR2_X1 U927 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U928 ( .A(KEYINPUT104), .B(n830), .Z(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U930 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  NAND2_X1 U937 ( .A1(n836), .A2(n835), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(G145) );
  XNOR2_X1 U939 ( .A(G1981), .B(KEYINPUT106), .ZN(n848) );
  XOR2_X1 U940 ( .A(G1976), .B(G1971), .Z(n840) );
  XNOR2_X1 U941 ( .A(G1966), .B(G1956), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U943 ( .A(G1961), .B(G1986), .Z(n842) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U946 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2474), .B(KEYINPUT41), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(G229) );
  XOR2_X1 U950 ( .A(KEYINPUT105), .B(G2090), .Z(n850) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2072), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U953 ( .A(n851), .B(G2096), .Z(n853) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2084), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U956 ( .A(G2678), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U957 ( .A(KEYINPUT42), .B(G2100), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U959 ( .A(n857), .B(n856), .Z(G227) );
  NAND2_X1 U960 ( .A1(G100), .A2(n892), .ZN(n859) );
  NAND2_X1 U961 ( .A1(G112), .A2(n887), .ZN(n858) );
  NAND2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n888), .A2(G124), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n894), .A2(G136), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U967 ( .A1(n864), .A2(n863), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT110), .B(KEYINPUT48), .Z(n866) );
  XNOR2_X1 U969 ( .A(KEYINPUT115), .B(KEYINPUT114), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U971 ( .A(n867), .B(KEYINPUT113), .Z(n870) );
  XNOR2_X1 U972 ( .A(n868), .B(KEYINPUT46), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U974 ( .A(n871), .B(G162), .Z(n874) );
  XOR2_X1 U975 ( .A(G160), .B(n872), .Z(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(n875), .B(n995), .Z(n886) );
  NAND2_X1 U978 ( .A1(n894), .A2(G139), .ZN(n876) );
  XOR2_X1 U979 ( .A(KEYINPUT111), .B(n876), .Z(n878) );
  NAND2_X1 U980 ( .A1(n892), .A2(G103), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U982 ( .A(KEYINPUT112), .B(n879), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G115), .A2(n887), .ZN(n881) );
  NAND2_X1 U984 ( .A1(G127), .A2(n888), .ZN(n880) );
  NAND2_X1 U985 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U986 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n1006) );
  XNOR2_X1 U988 ( .A(G164), .B(n1006), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n902) );
  NAND2_X1 U990 ( .A1(G118), .A2(n887), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G130), .A2(n888), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U993 ( .A(KEYINPUT107), .B(n891), .Z(n900) );
  NAND2_X1 U994 ( .A1(n892), .A2(G106), .ZN(n893) );
  XNOR2_X1 U995 ( .A(KEYINPUT108), .B(n893), .ZN(n897) );
  NAND2_X1 U996 ( .A1(n894), .A2(G142), .ZN(n895) );
  XOR2_X1 U997 ( .A(KEYINPUT109), .B(n895), .Z(n896) );
  NAND2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U999 ( .A(n898), .B(KEYINPUT45), .Z(n899) );
  NOR2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1001 ( .A(n902), .B(n901), .Z(n904) );
  XOR2_X1 U1002 ( .A(n904), .B(n903), .Z(n905) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n905), .ZN(G395) );
  XOR2_X1 U1004 ( .A(n906), .B(G286), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G171), .B(n935), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n909), .B(n927), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n910), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(KEYINPUT116), .B(n911), .ZN(G397) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n912), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1018 ( .A(KEYINPUT56), .B(G16), .ZN(n944) );
  XNOR2_X1 U1019 ( .A(n918), .B(G1956), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(n919), .B(KEYINPUT123), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(G1971), .A2(G303), .ZN(n920) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n931) );
  XNOR2_X1 U1024 ( .A(G171), .B(G1961), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n927), .B(n926), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1030 ( .A(KEYINPUT124), .B(n934), .Z(n937) );
  XOR2_X1 U1031 ( .A(n935), .B(G1341), .Z(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(G1966), .B(G168), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(n940), .B(KEYINPUT57), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n1024) );
  XNOR2_X1 U1038 ( .A(G1986), .B(G24), .ZN(n949) );
  XNOR2_X1 U1039 ( .A(G1971), .B(G22), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G1976), .B(G23), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(KEYINPUT127), .B(n947), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT58), .B(n950), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G21), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G5), .B(G1961), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n965) );
  XOR2_X1 U1049 ( .A(G19), .B(G1341), .Z(n958) );
  XNOR2_X1 U1050 ( .A(G1956), .B(G20), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(G1981), .B(G6), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1054 ( .A(KEYINPUT59), .B(G1348), .Z(n959) );
  XNOR2_X1 U1055 ( .A(G4), .B(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1057 ( .A(KEYINPUT60), .B(n962), .Z(n963) );
  XNOR2_X1 U1058 ( .A(KEYINPUT126), .B(n963), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n966), .B(KEYINPUT61), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT125), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n969), .ZN(n1022) );
  XNOR2_X1 U1064 ( .A(G2072), .B(KEYINPUT121), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n970), .B(G33), .ZN(n975) );
  XOR2_X1 U1066 ( .A(n971), .B(G27), .Z(n973) );
  XNOR2_X1 U1067 ( .A(G1996), .B(G32), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(KEYINPUT120), .B(G2067), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(G26), .B(n976), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1073 ( .A(KEYINPUT122), .B(n979), .Z(n981) );
  XNOR2_X1 U1074 ( .A(G1991), .B(G25), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(G28), .A2(n982), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(n983), .B(KEYINPUT53), .ZN(n986) );
  XOR2_X1 U1078 ( .A(G2084), .B(G34), .Z(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT54), .B(n984), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(G35), .B(G2090), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(G29), .A2(n989), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(n990), .B(KEYINPUT55), .ZN(n1020) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1087 ( .A(KEYINPUT51), .B(n993), .Z(n994) );
  XNOR2_X1 U1088 ( .A(KEYINPUT118), .B(n994), .ZN(n1013) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G2084), .B(G160), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(KEYINPUT117), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1011) );
  XOR2_X1 U1096 ( .A(G2072), .B(n1006), .Z(n1008) );
  XOR2_X1 U1097 ( .A(G164), .B(G2078), .Z(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1099 ( .A(KEYINPUT50), .B(n1009), .Z(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(n1017), .B(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(G29), .A2(n1018), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

