//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n469), .B(KEYINPUT65), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n463), .A2(new_n464), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G125), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n458), .B1(new_n477), .B2(new_n470), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT66), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n468), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n480), .B(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n466), .A2(G136), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT69), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n465), .A2(new_n458), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G124), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n484), .A2(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(new_n476), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n458), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI22_X1  g069(.A1(new_n491), .A2(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n466), .A2(G138), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n466), .A2(new_n498), .A3(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  AND3_X1   g086(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(G543), .B1(KEYINPUT70), .B2(KEYINPUT5), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n505), .A2(KEYINPUT71), .A3(new_n510), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI221_X1 g096(.A(new_n508), .B1(new_n509), .B2(new_n511), .C1(new_n520), .C2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n511), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT74), .B(G51), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n516), .A2(new_n517), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT71), .B1(new_n505), .B2(new_n510), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(G76), .A2(G543), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n507), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n527), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n505), .B(KEYINPUT72), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G63), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n532), .A2(new_n533), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n507), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n535), .A2(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n505), .B(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n525), .A2(G52), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n530), .A2(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n536), .A2(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n507), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n511), .B(KEYINPUT73), .ZN(new_n554));
  INV_X1    g129(.A(G43), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n520), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  AND2_X1   g138(.A1(new_n510), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(new_n565), .A3(G53), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n511), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n566), .A2(new_n571), .A3(new_n568), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT77), .B1(new_n528), .B2(new_n529), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n518), .A2(new_n575), .A3(new_n519), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(G91), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n505), .A2(G65), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT78), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n573), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  INV_X1    g159(.A(G74), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n507), .B1(new_n543), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(G49), .B2(new_n564), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n574), .A2(new_n576), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G87), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(new_n588), .A2(G86), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n505), .A2(G61), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n597), .A3(G651), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n596), .A2(new_n598), .B1(G48), .B2(new_n564), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n591), .A2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n530), .A2(G85), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT80), .B(G47), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n525), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n601), .B(new_n603), .C1(new_n604), .C2(new_n507), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n505), .A2(G66), .ZN(new_n607));
  INV_X1    g182(.A(G79), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n502), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n525), .A2(G54), .B1(G651), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n574), .A2(G92), .A3(new_n576), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(KEYINPUT81), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n574), .A2(new_n614), .A3(G92), .A4(new_n576), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n613), .B1(new_n612), .B2(new_n615), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n606), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n606), .B1(new_n619), .B2(G868), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n582), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(G868), .B2(new_n582), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n619), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n619), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n460), .A2(new_n476), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT13), .Z(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n466), .A2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n488), .A2(G123), .ZN(new_n638));
  OR2_X1    g213(.A1(G99), .A2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n639), .B(G2104), .C1(G111), .C2(new_n458), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n637), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2096), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n635), .A2(new_n636), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT84), .ZN(G401));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n666), .B1(new_n662), .B2(new_n665), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n664), .B2(new_n665), .ZN(new_n669));
  INV_X1    g244(.A(new_n665), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n670), .A2(new_n666), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n662), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  OR3_X1    g248(.A1(new_n667), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  MUX2_X1   g265(.A(new_n690), .B(new_n689), .S(new_n682), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n694), .A2(new_n695), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(new_n695), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n700), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT26), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G129), .B2(new_n488), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n460), .A2(G105), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n466), .A2(G141), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(KEYINPUT95), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(KEYINPUT95), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G32), .B(new_n713), .S(G29), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G27), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G164), .B2(new_n717), .ZN(new_n719));
  INV_X1    g294(.A(G2078), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G29), .A2(G33), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT93), .Z(new_n723));
  NAND3_X1  g298(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT25), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n476), .A2(G127), .ZN(new_n726));
  NAND2_X1  g301(.A1(G115), .A2(G2104), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n458), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI211_X1 g303(.A(new_n725), .B(new_n728), .C1(G139), .C2(new_n466), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n723), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G2072), .Z(new_n731));
  NAND3_X1  g306(.A1(new_n716), .A2(new_n721), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G29), .A2(G35), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G162), .B2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT29), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2090), .ZN(new_n736));
  NOR2_X1   g311(.A1(G16), .A2(G19), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n558), .B2(G16), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(G1341), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n717), .A2(G26), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT28), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n466), .A2(G140), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n488), .A2(G128), .ZN(new_n743));
  OR2_X1    g318(.A1(G104), .A2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT92), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n742), .A2(new_n743), .A3(KEYINPUT92), .A4(new_n745), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n741), .B1(new_n750), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2067), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n738), .A2(G1341), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n739), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n732), .A2(new_n736), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G16), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G20), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT23), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n582), .B2(new_n756), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1956), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT24), .B(G34), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(new_n717), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT94), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n480), .B(KEYINPUT68), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n717), .ZN(new_n766));
  INV_X1    g341(.A(G2084), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G1961), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n756), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n756), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT97), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n768), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  AND3_X1   g348(.A1(new_n755), .A2(new_n761), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n619), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G4), .B2(G16), .ZN(new_n776));
  INV_X1    g351(.A(G1348), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n756), .A2(G21), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G168), .B2(new_n756), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G1966), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT96), .Z(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT30), .B(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n784), .A2(new_n717), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n641), .B2(new_n717), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n781), .B2(G1966), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n783), .B(new_n789), .C1(new_n769), .C2(new_n772), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT98), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n779), .B(new_n791), .C1(new_n777), .C2(new_n776), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n756), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n756), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1971), .ZN(new_n795));
  NOR2_X1   g370(.A1(G6), .A2(G16), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n591), .A2(new_n599), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G23), .B(G288), .S(G16), .Z(new_n801));
  XOR2_X1   g376(.A(KEYINPUT33), .B(G1976), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT90), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n801), .B(new_n803), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n800), .B(new_n804), .C1(new_n798), .C2(new_n799), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n756), .A2(G24), .ZN(new_n808));
  INV_X1    g383(.A(G290), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n756), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1986), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n717), .A2(G25), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT88), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n466), .A2(G131), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n488), .A2(G119), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n458), .A2(G107), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n814), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT89), .Z(new_n819));
  AOI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(G29), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  AOI211_X1 g397(.A(new_n811), .B(new_n822), .C1(KEYINPUT91), .C2(KEYINPUT36), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n806), .A2(new_n807), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n792), .A2(new_n826), .A3(new_n827), .ZN(G311));
  INV_X1    g403(.A(G311), .ZN(G150));
  NAND2_X1  g404(.A1(new_n619), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n536), .A2(G67), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n507), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G55), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n554), .A2(new_n835), .B1(new_n836), .B2(new_n520), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n558), .A2(new_n838), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n557), .A2(new_n553), .B1(new_n834), .B2(new_n837), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n831), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n842), .ZN(new_n845));
  INV_X1    g420(.A(new_n838), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n845), .A2(new_n849), .ZN(G145));
  INV_X1    g425(.A(new_n641), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n765), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(G160), .A2(new_n641), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n852), .A2(new_n853), .A3(G162), .ZN(new_n854));
  AOI21_X1  g429(.A(G162), .B1(new_n852), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n497), .A2(new_n499), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n495), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n493), .A2(new_n494), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n488), .B2(G126), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT100), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n857), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n711), .B2(new_n712), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n711), .A2(new_n712), .A3(new_n863), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT101), .B1(new_n748), .B2(new_n749), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n748), .A2(KEYINPUT101), .A3(new_n749), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n865), .B(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n867), .ZN(new_n870));
  INV_X1    g445(.A(new_n866), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(new_n864), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n729), .B(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n869), .A2(new_n876), .A3(new_n729), .A4(new_n872), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n488), .A2(G130), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n458), .A2(G118), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(G142), .B2(new_n466), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n818), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n633), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT103), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n856), .B1(new_n878), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n875), .A2(KEYINPUT103), .A3(new_n886), .A4(new_n877), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n875), .A2(new_n886), .A3(new_n877), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n886), .B1(new_n875), .B2(new_n877), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n856), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g471(.A(new_n627), .B(new_n841), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n618), .A2(G299), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n582), .B(new_n610), .C1(new_n616), .C2(new_n617), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n612), .A2(new_n615), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT10), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n582), .B1(new_n909), .B2(new_n610), .ZN(new_n910));
  INV_X1    g485(.A(new_n900), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n898), .A2(KEYINPUT104), .A3(new_n900), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n904), .B1(new_n897), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(G288), .A2(G166), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n587), .A2(new_n589), .A3(G303), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(G305), .A2(new_n809), .ZN(new_n919));
  NAND3_X1  g494(.A1(G290), .A2(new_n591), .A3(new_n599), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n916), .A2(new_n919), .A3(new_n917), .A4(new_n920), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT42), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n922), .A2(KEYINPUT105), .A3(new_n923), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT105), .B1(new_n922), .B2(new_n923), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n924), .B2(KEYINPUT106), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n926), .B1(new_n930), .B2(KEYINPUT42), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n915), .B(new_n931), .Z(new_n932));
  MUX2_X1   g507(.A(new_n846), .B(new_n932), .S(G868), .Z(G295));
  MUX2_X1   g508(.A(new_n846), .B(new_n932), .S(G868), .Z(G331));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  NAND2_X1  g510(.A1(G168), .A2(G301), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n547), .A2(new_n548), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n937), .B(new_n546), .C1(new_n535), .C2(new_n539), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n841), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n936), .A2(new_n938), .A3(new_n839), .A4(new_n840), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n901), .B2(new_n902), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n924), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n922), .A2(KEYINPUT105), .A3(new_n923), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n942), .A2(new_n898), .A3(new_n900), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  XNOR2_X1  g526(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT41), .B1(new_n910), .B2(new_n911), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n942), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n949), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n929), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n954), .B2(new_n955), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n943), .B1(new_n902), .B2(KEYINPUT108), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n912), .A2(new_n913), .A3(new_n942), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n929), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n950), .A2(new_n951), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n935), .B1(new_n959), .B2(new_n968), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n963), .A2(new_n965), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n958), .A2(new_n950), .A3(new_n951), .ZN(new_n971));
  INV_X1    g546(.A(new_n952), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n953), .A2(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n969), .B1(new_n935), .B2(new_n973), .ZN(G397));
  XOR2_X1   g549(.A(new_n750), .B(G2067), .Z(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT109), .ZN(new_n976));
  INV_X1    g551(.A(G1996), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n713), .B(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n818), .B(new_n821), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n863), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(KEYINPUT45), .ZN(new_n986));
  INV_X1    g561(.A(G40), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n987), .B(new_n468), .C1(new_n479), .C2(new_n475), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n983), .A2(new_n990), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n989), .A2(G1986), .A3(G290), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT124), .B(KEYINPUT48), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n821), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n819), .A2(new_n995), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n980), .A2(new_n996), .B1(G2067), .B2(new_n750), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n991), .A2(new_n994), .B1(new_n990), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n990), .B1(new_n976), .B2(new_n713), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT123), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n990), .A2(new_n977), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT46), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n998), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n863), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(G164), .B2(G1384), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n988), .A3(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(G2078), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G164), .A2(G1384), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n857), .A2(new_n861), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n984), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n480), .A2(G40), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n985), .B2(new_n1015), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1011), .A2(new_n1012), .B1(new_n1023), .B2(new_n769), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n988), .B1(new_n1018), .B2(new_n1008), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n720), .A2(KEYINPUT53), .ZN(new_n1026));
  OR3_X1    g601(.A1(new_n986), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G301), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT113), .B(G1981), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n797), .A2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n530), .A2(G86), .ZN(new_n1031));
  INV_X1    g606(.A(G48), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n595), .B1(new_n1032), .B2(new_n511), .ZN(new_n1033));
  OAI21_X1  g608(.A(G1981), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n863), .A2(new_n984), .ZN(new_n1038));
  OAI21_X1  g613(.A(G8), .B1(new_n1021), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1042));
  AOI211_X1 g617(.A(KEYINPUT114), .B(KEYINPUT49), .C1(new_n1030), .C2(new_n1034), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G288), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(new_n1039), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1044), .A2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT110), .B(G1971), .Z(new_n1053));
  NAND2_X1  g628(.A1(new_n1010), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1023), .B2(G2090), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1058), .B2(KEYINPUT55), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(KEYINPUT112), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(KEYINPUT55), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1055), .A2(G8), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1017), .A2(new_n1015), .A3(new_n984), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n988), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1015), .B1(new_n863), .B2(new_n984), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1054), .B1(new_n1068), .B2(G2090), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1063), .B1(new_n1069), .B2(G8), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1052), .A2(new_n1064), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1020), .A2(new_n1022), .A3(new_n767), .ZN(new_n1072));
  INV_X1    g647(.A(G1966), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n986), .B2(new_n1025), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1074), .A3(G168), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT51), .B1(new_n1075), .B2(G8), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(KEYINPUT122), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G8), .ZN(new_n1080));
  AOI211_X1 g655(.A(new_n1080), .B(G168), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1076), .B2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1079), .A2(KEYINPUT62), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1028), .B(new_n1071), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1070), .A2(KEYINPUT63), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1080), .B(G286), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1064), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G288), .A2(G1976), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1044), .A2(new_n1090), .B1(new_n797), .B2(new_n1029), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1089), .A2(new_n1052), .B1(new_n1091), .B2(new_n1039), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1044), .A2(new_n1088), .A3(new_n1051), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1055), .A2(G8), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1063), .B1(new_n1095), .B2(KEYINPUT115), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(KEYINPUT115), .B2(new_n1095), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1093), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1086), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n566), .A2(new_n1101), .A3(new_n568), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n569), .A2(KEYINPUT117), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(new_n577), .A3(new_n581), .A4(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(KEYINPUT118), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(KEYINPUT118), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1007), .A2(new_n988), .A3(new_n1009), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n582), .A2(KEYINPUT57), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1110), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1021), .A2(new_n1038), .A3(G2067), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(new_n1023), .B2(new_n777), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1119), .B2(new_n618), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1109), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1116), .B1(new_n1121), .B2(new_n1107), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1119), .A2(KEYINPUT60), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(new_n619), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(KEYINPUT60), .B2(new_n1119), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1117), .A3(KEYINPUT61), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1007), .A2(new_n988), .A3(new_n977), .A4(new_n1009), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT58), .B(G1341), .Z(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1021), .B2(new_n1038), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1130), .B1(new_n1134), .B2(new_n558), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n558), .ZN(new_n1137));
  AOI211_X1 g712(.A(KEYINPUT119), .B(new_n1137), .C1(new_n1131), .C2(new_n1133), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1129), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1135), .A2(new_n1138), .A3(KEYINPUT59), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1128), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1117), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1115), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT120), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1142), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1127), .B1(new_n1150), .B2(KEYINPUT121), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n1152), .B(new_n1142), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1124), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n1155));
  INV_X1    g730(.A(new_n986), .ZN(new_n1156));
  NOR4_X1   g731(.A1(new_n468), .A2(new_n478), .A3(new_n987), .A4(new_n1026), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1007), .A3(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1024), .A2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1159), .A2(G301), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1155), .B1(new_n1160), .B2(new_n1028), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1024), .A2(G301), .A3(new_n1027), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1162), .B(KEYINPUT54), .C1(new_n1159), .C2(G301), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1071), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1100), .B1(new_n1154), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n983), .ZN(new_n1167));
  XOR2_X1   g742(.A(G290), .B(G1986), .Z(new_n1168));
  AOI21_X1  g743(.A(new_n989), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1006), .B1(new_n1166), .B2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n677), .A2(G319), .A3(new_n678), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n1173), .A2(KEYINPUT125), .ZN(new_n1174));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n1175));
  NAND4_X1  g749(.A1(new_n677), .A2(new_n1175), .A3(G319), .A4(new_n678), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n703), .A2(new_n659), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g752(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n895), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g754(.A(new_n1172), .B1(new_n973), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n890), .B2(new_n894), .ZN(new_n1182));
  AND2_X1   g756(.A1(new_n971), .A2(new_n972), .ZN(new_n1183));
  NAND3_X1  g757(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n1184));
  NOR2_X1   g758(.A1(new_n1184), .A2(new_n966), .ZN(new_n1185));
  OAI211_X1 g759(.A(new_n1182), .B(KEYINPUT126), .C1(new_n1183), .C2(new_n1185), .ZN(new_n1186));
  AND3_X1   g760(.A1(new_n1181), .A2(KEYINPUT127), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g761(.A(KEYINPUT127), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1188));
  NOR2_X1   g762(.A1(new_n1187), .A2(new_n1188), .ZN(G308));
  NAND2_X1  g763(.A1(new_n1181), .A2(new_n1186), .ZN(G225));
endmodule


