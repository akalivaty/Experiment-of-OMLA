

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U320 ( .A(G113GAT), .B(G197GAT), .Z(n288) );
  NOR2_X1 U321 ( .A1(n553), .A2(n372), .ZN(n374) );
  XOR2_X1 U322 ( .A(G169GAT), .B(G8GAT), .Z(n331) );
  NOR2_X1 U323 ( .A1(n568), .A2(n462), .ZN(n426) );
  XNOR2_X1 U324 ( .A(n355), .B(n288), .ZN(n336) );
  XNOR2_X1 U325 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U326 ( .A(n573), .B(KEYINPUT41), .Z(n547) );
  XNOR2_X1 U327 ( .A(n377), .B(KEYINPUT69), .ZN(n556) );
  INV_X1 U328 ( .A(n556), .ZN(n532) );
  XOR2_X1 U329 ( .A(n448), .B(n447), .Z(n557) );
  XOR2_X1 U330 ( .A(n462), .B(KEYINPUT28), .Z(n525) );
  XNOR2_X1 U331 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U332 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(G43GAT), .B(G29GAT), .Z(n290) );
  XNOR2_X1 U334 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n289) );
  XNOR2_X1 U335 ( .A(n290), .B(n289), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n291), .B(KEYINPUT67), .ZN(n293) );
  XOR2_X1 U337 ( .A(G36GAT), .B(KEYINPUT8), .Z(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n339) );
  XOR2_X1 U339 ( .A(G190GAT), .B(KEYINPUT77), .Z(n316) );
  XOR2_X1 U340 ( .A(n316), .B(G106GAT), .Z(n295) );
  XNOR2_X1 U341 ( .A(G134GAT), .B(G218GAT), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n339), .B(n296), .ZN(n298) );
  AND2_X1 U344 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U346 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n300) );
  XNOR2_X1 U347 ( .A(G162GAT), .B(KEYINPUT76), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n310) );
  XOR2_X1 U350 ( .A(KEYINPUT72), .B(G85GAT), .Z(n304) );
  XNOR2_X1 U351 ( .A(G99GAT), .B(KEYINPUT71), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U353 ( .A(G92GAT), .B(n305), .Z(n351) );
  XOR2_X1 U354 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n307) );
  XNOR2_X1 U355 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n351), .B(n308), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n449) );
  XOR2_X1 U359 ( .A(KEYINPUT18), .B(KEYINPUT81), .Z(n312) );
  XNOR2_X1 U360 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U362 ( .A(KEYINPUT19), .B(n313), .Z(n446) );
  XOR2_X1 U363 ( .A(G176GAT), .B(G64GAT), .Z(n346) );
  XOR2_X1 U364 ( .A(n346), .B(KEYINPUT92), .Z(n315) );
  NAND2_X1 U365 ( .A1(G226GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n317) );
  XOR2_X1 U367 ( .A(n317), .B(n316), .Z(n326) );
  XOR2_X1 U368 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n319) );
  XNOR2_X1 U369 ( .A(G218GAT), .B(KEYINPUT84), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U371 ( .A(n320), .B(G211GAT), .Z(n322) );
  XNOR2_X1 U372 ( .A(G197GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n421) );
  XNOR2_X1 U374 ( .A(G36GAT), .B(n331), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n323), .B(G92GAT), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n421), .B(n324), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U378 ( .A(n446), .B(n327), .Z(n519) );
  INV_X1 U379 ( .A(n519), .ZN(n385) );
  INV_X1 U380 ( .A(n449), .ZN(n553) );
  XOR2_X1 U381 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n329) );
  XNOR2_X1 U382 ( .A(KEYINPUT66), .B(KEYINPUT29), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U384 ( .A(G141GAT), .B(G22GAT), .Z(n413) );
  XNOR2_X1 U385 ( .A(n330), .B(n413), .ZN(n335) );
  XOR2_X1 U386 ( .A(n331), .B(KEYINPUT65), .Z(n333) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n337) );
  XOR2_X1 U390 ( .A(G15GAT), .B(G1GAT), .Z(n355) );
  XOR2_X1 U391 ( .A(n339), .B(n338), .Z(n377) );
  XNOR2_X1 U392 ( .A(G106GAT), .B(G78GAT), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n340), .B(G148GAT), .ZN(n416) );
  XOR2_X1 U394 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n341) );
  XNOR2_X1 U395 ( .A(n416), .B(n341), .ZN(n345) );
  XOR2_X1 U396 ( .A(KEYINPUT70), .B(KEYINPUT31), .Z(n343) );
  XNOR2_X1 U397 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n350) );
  XOR2_X1 U400 ( .A(KEYINPUT13), .B(G57GAT), .Z(n366) );
  XOR2_X1 U401 ( .A(n366), .B(n346), .Z(n348) );
  NAND2_X1 U402 ( .A1(G230GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n353) );
  XOR2_X1 U405 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XNOR2_X1 U406 ( .A(n435), .B(n351), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n573) );
  NAND2_X1 U408 ( .A1(n377), .A2(n547), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n354), .B(KEYINPUT46), .ZN(n371) );
  XNOR2_X1 U410 ( .A(n355), .B(G127GAT), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n356), .B(G71GAT), .ZN(n370) );
  XOR2_X1 U412 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n358) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U415 ( .A(KEYINPUT14), .B(G64GAT), .Z(n360) );
  XNOR2_X1 U416 ( .A(G8GAT), .B(G78GAT), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U418 ( .A(n362), .B(n361), .Z(n368) );
  XOR2_X1 U419 ( .A(G211GAT), .B(G155GAT), .Z(n364) );
  XNOR2_X1 U420 ( .A(G22GAT), .B(G183GAT), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U424 ( .A(n370), .B(n369), .Z(n577) );
  INV_X1 U425 ( .A(n577), .ZN(n489) );
  NAND2_X1 U426 ( .A1(n371), .A2(n489), .ZN(n372) );
  XNOR2_X1 U427 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n375), .B(KEYINPUT47), .ZN(n382) );
  XOR2_X1 U430 ( .A(KEYINPUT36), .B(n553), .Z(n581) );
  NOR2_X1 U431 ( .A1(n581), .A2(n489), .ZN(n376) );
  XNOR2_X1 U432 ( .A(KEYINPUT45), .B(n376), .ZN(n380) );
  INV_X1 U433 ( .A(n573), .ZN(n378) );
  AND2_X1 U434 ( .A1(n378), .A2(n556), .ZN(n379) );
  AND2_X1 U435 ( .A1(n380), .A2(n379), .ZN(n381) );
  NOR2_X1 U436 ( .A1(n382), .A2(n381), .ZN(n384) );
  INV_X1 U437 ( .A(KEYINPUT48), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n526) );
  NAND2_X1 U439 ( .A1(n385), .A2(n526), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n386), .B(KEYINPUT54), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n387), .B(KEYINPUT117), .ZN(n409) );
  XOR2_X1 U442 ( .A(G127GAT), .B(KEYINPUT0), .Z(n389) );
  XNOR2_X1 U443 ( .A(G113GAT), .B(G134GAT), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n438) );
  XOR2_X1 U445 ( .A(G85GAT), .B(n438), .Z(n391) );
  NAND2_X1 U446 ( .A1(G225GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U448 ( .A(G29GAT), .B(n392), .ZN(n408) );
  XOR2_X1 U449 ( .A(G57GAT), .B(G148GAT), .Z(n394) );
  XNOR2_X1 U450 ( .A(G141GAT), .B(G120GAT), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U452 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n396) );
  XNOR2_X1 U453 ( .A(G1GAT), .B(KEYINPUT90), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U455 ( .A(n398), .B(n397), .Z(n406) );
  XOR2_X1 U456 ( .A(KEYINPUT85), .B(G162GAT), .Z(n400) );
  XNOR2_X1 U457 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U459 ( .A(KEYINPUT2), .B(n401), .Z(n422) );
  XOR2_X1 U460 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n403) );
  XNOR2_X1 U461 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n422), .B(n404), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U465 ( .A(n408), .B(n407), .Z(n467) );
  INV_X1 U466 ( .A(n467), .ZN(n516) );
  NAND2_X1 U467 ( .A1(n409), .A2(n516), .ZN(n568) );
  XOR2_X1 U468 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n411) );
  XNOR2_X1 U469 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U471 ( .A(n412), .B(KEYINPUT24), .Z(n415) );
  XNOR2_X1 U472 ( .A(G50GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n420) );
  XOR2_X1 U474 ( .A(n416), .B(KEYINPUT23), .Z(n418) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U477 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n462) );
  XNOR2_X1 U480 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  NAND2_X1 U482 ( .A1(KEYINPUT118), .A2(n427), .ZN(n431) );
  INV_X1 U483 ( .A(KEYINPUT118), .ZN(n429) );
  INV_X1 U484 ( .A(n427), .ZN(n428) );
  NAND2_X1 U485 ( .A1(n429), .A2(n428), .ZN(n430) );
  NAND2_X1 U486 ( .A1(n431), .A2(n430), .ZN(n559) );
  XOR2_X1 U487 ( .A(KEYINPUT80), .B(G190GAT), .Z(n433) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(G15GAT), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U490 ( .A(n434), .B(G99GAT), .Z(n437) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n442) );
  XOR2_X1 U493 ( .A(n438), .B(KEYINPUT82), .Z(n440) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n442), .B(n441), .Z(n448) );
  XOR2_X1 U497 ( .A(KEYINPUT20), .B(G176GAT), .Z(n444) );
  XNOR2_X1 U498 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  INV_X1 U501 ( .A(n557), .ZN(n459) );
  NAND2_X1 U502 ( .A1(n559), .A2(n459), .ZN(n453) );
  NOR2_X1 U503 ( .A1(n449), .A2(n453), .ZN(n452) );
  XNOR2_X1 U504 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n450) );
  NOR2_X1 U505 ( .A1(n489), .A2(n453), .ZN(n456) );
  XNOR2_X1 U506 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(G183GAT), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n456), .B(n455), .ZN(G1350GAT) );
  NOR2_X1 U509 ( .A1(n556), .A2(n573), .ZN(n492) );
  XNOR2_X1 U510 ( .A(KEYINPUT27), .B(n519), .ZN(n464) );
  NOR2_X1 U511 ( .A1(n516), .A2(n464), .ZN(n527) );
  NAND2_X1 U512 ( .A1(n525), .A2(n527), .ZN(n457) );
  XOR2_X1 U513 ( .A(KEYINPUT93), .B(n457), .Z(n458) );
  NOR2_X1 U514 ( .A1(n459), .A2(n458), .ZN(n471) );
  NOR2_X1 U515 ( .A1(n519), .A2(n557), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n462), .A2(n460), .ZN(n461) );
  XOR2_X1 U517 ( .A(KEYINPUT25), .B(n461), .Z(n466) );
  NAND2_X1 U518 ( .A1(n557), .A2(n462), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT26), .ZN(n569) );
  NOR2_X1 U520 ( .A1(n569), .A2(n464), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n466), .A2(n465), .ZN(n468) );
  NOR2_X1 U522 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U523 ( .A(n469), .B(KEYINPUT94), .ZN(n470) );
  NOR2_X1 U524 ( .A1(n471), .A2(n470), .ZN(n488) );
  NOR2_X1 U525 ( .A1(n553), .A2(n489), .ZN(n472) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(n472), .Z(n473) );
  NOR2_X1 U527 ( .A1(n488), .A2(n473), .ZN(n503) );
  NAND2_X1 U528 ( .A1(n492), .A2(n503), .ZN(n483) );
  NOR2_X1 U529 ( .A1(n516), .A2(n483), .ZN(n478) );
  XOR2_X1 U530 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n475) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(KEYINPUT96), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT95), .B(n476), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U535 ( .A1(n519), .A2(n483), .ZN(n479) );
  XOR2_X1 U536 ( .A(G8GAT), .B(n479), .Z(G1325GAT) );
  NOR2_X1 U537 ( .A1(n557), .A2(n483), .ZN(n481) );
  XNOR2_X1 U538 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U541 ( .A1(n525), .A2(n483), .ZN(n485) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1327GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n487) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT100), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n496) );
  XOR2_X1 U547 ( .A(KEYINPUT38), .B(KEYINPUT101), .Z(n494) );
  NOR2_X1 U548 ( .A1(n581), .A2(n488), .ZN(n490) );
  NAND2_X1 U549 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT37), .B(n491), .ZN(n515) );
  NAND2_X1 U551 ( .A1(n492), .A2(n515), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(n501) );
  NOR2_X1 U553 ( .A1(n516), .A2(n501), .ZN(n495) );
  XOR2_X1 U554 ( .A(n496), .B(n495), .Z(G1328GAT) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n498) );
  NOR2_X1 U556 ( .A1(n519), .A2(n501), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1329GAT) );
  NOR2_X1 U558 ( .A1(n501), .A2(n557), .ZN(n499) );
  XOR2_X1 U559 ( .A(KEYINPUT40), .B(n499), .Z(n500) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NOR2_X1 U561 ( .A1(n525), .A2(n501), .ZN(n502) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n502), .Z(G1331GAT) );
  INV_X1 U563 ( .A(n547), .ZN(n562) );
  NOR2_X1 U564 ( .A1(n377), .A2(n562), .ZN(n514) );
  NAND2_X1 U565 ( .A1(n514), .A2(n503), .ZN(n510) );
  NOR2_X1 U566 ( .A1(n516), .A2(n510), .ZN(n504) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n504), .Z(n505) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n519), .A2(n510), .ZN(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n557), .A2(n510), .ZN(n509) );
  XOR2_X1 U574 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U575 ( .A1(n525), .A2(n510), .ZN(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n522) );
  NOR2_X1 U580 ( .A1(n516), .A2(n522), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n522), .ZN(n520) );
  XOR2_X1 U584 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U585 ( .A1(n557), .A2(n522), .ZN(n521) );
  XOR2_X1 U586 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U587 ( .A1(n525), .A2(n522), .ZN(n523) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(n523), .Z(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT112), .ZN(n534) );
  INV_X1 U591 ( .A(n525), .ZN(n531) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(KEYINPUT110), .B(n528), .ZN(n545) );
  OR2_X1 U594 ( .A1(n557), .A2(n545), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT111), .B(n529), .Z(n530) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n532), .A2(n542), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U600 ( .A1(n542), .A2(n547), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  NAND2_X1 U603 ( .A1(n542), .A2(n577), .ZN(n541) );
  XOR2_X1 U604 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n539) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U609 ( .A1(n542), .A2(n553), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NOR2_X1 U611 ( .A1(n545), .A2(n569), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n377), .A2(n554), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U615 ( .A1(n554), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n554), .A2(n577), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(KEYINPUT116), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(n552), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  AND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT120), .B(n560), .Z(n561) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n561), .ZN(G1348GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n453), .ZN(n567) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n564) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT56), .B(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NOR2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n579), .A2(n377), .ZN(n572) );
  XOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT60), .Z(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT59), .B(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n579), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n579), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U644 ( .A(n579), .ZN(n580) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

