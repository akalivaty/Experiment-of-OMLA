//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n572, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OR2_X1    g045(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n476), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n464), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n479), .A2(G137), .A3(new_n473), .A4(new_n467), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(G101), .A3(G2104), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT68), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n480), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n480), .B2(new_n483), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n475), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  OAI221_X1 g063(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n473), .C2(G112), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n464), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT67), .B1(new_n464), .B2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n467), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n464), .A2(G2104), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n477), .B2(new_n478), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n494), .A2(new_n474), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G124), .ZN(new_n499));
  INV_X1    g074(.A(G136), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n494), .A2(new_n481), .A3(new_n497), .ZN(new_n501));
  OAI221_X1 g076(.A(new_n489), .B1(new_n498), .B2(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G162));
  NAND3_X1  g078(.A1(new_n481), .A2(G102), .A3(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(G114), .A2(G2104), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(new_n496), .B2(G126), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n504), .B1(new_n507), .B2(new_n481), .ZN(new_n508));
  INV_X1    g083(.A(G138), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n471), .B2(new_n472), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n510), .A2(new_n479), .A3(KEYINPUT4), .A4(new_n467), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n514));
  OAI21_X1  g089(.A(G138), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n515), .B2(new_n468), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n508), .A2(new_n517), .ZN(G164));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT72), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT5), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n520), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n522), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n527), .A2(G651), .B1(new_n531), .B2(G50), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n523), .A2(new_n525), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n528), .A2(new_n529), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(KEYINPUT71), .B1(new_n526), .B2(new_n530), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n532), .B1(new_n533), .B2(new_n539), .ZN(G303));
  INV_X1    g115(.A(G303), .ZN(G166));
  XOR2_X1   g116(.A(KEYINPUT73), .B(G51), .Z(new_n542));
  NAND2_X1  g117(.A1(new_n531), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n537), .A2(new_n538), .A3(G89), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n545), .A2(KEYINPUT74), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(KEYINPUT74), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n543), .B(new_n544), .C1(new_n548), .C2(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  AND2_X1   g126(.A1(new_n537), .A2(new_n538), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G90), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G651), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n531), .A2(G52), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n553), .A2(new_n556), .A3(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  XNOR2_X1  g134(.A(KEYINPUT76), .B(G81), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n537), .A2(new_n538), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G43), .ZN(new_n562));
  INV_X1    g137(.A(new_n531), .ZN(new_n563));
  NAND2_X1  g138(.A1(G68), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G56), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n526), .B2(new_n565), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n566), .A2(KEYINPUT75), .A3(G651), .ZN(new_n567));
  AOI21_X1  g142(.A(KEYINPUT75), .B1(new_n566), .B2(G651), .ZN(new_n568));
  OAI221_X1 g143(.A(new_n561), .B1(new_n562), .B2(new_n563), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  AND3_X1   g146(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G36), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(G188));
  OAI211_X1 g151(.A(G53), .B(G543), .C1(new_n528), .C2(new_n529), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n526), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  INV_X1    g157(.A(G91), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n578), .B(new_n582), .C1(new_n539), .C2(new_n583), .ZN(G299));
  NAND3_X1  g159(.A1(new_n537), .A2(new_n538), .A3(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n531), .A2(G49), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT77), .ZN(G288));
  NAND2_X1  g164(.A1(new_n531), .A2(G48), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n552), .A2(G86), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n534), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n555), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n526), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n531), .A2(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n600), .B(new_n601), .C1(new_n539), .C2(new_n602), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT79), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n539), .A2(KEYINPUT10), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n526), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(new_n531), .B2(G54), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT10), .B1(new_n539), .B2(new_n606), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n607), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n605), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n605), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(G299), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G168), .B2(new_n617), .ZN(G297));
  XOR2_X1   g194(.A(G297), .B(KEYINPUT80), .Z(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n569), .A2(new_n617), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n613), .A2(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g201(.A(new_n498), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G123), .ZN(new_n628));
  INV_X1    g203(.A(new_n501), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G135), .ZN(new_n630));
  OAI221_X1 g205(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n473), .C2(G111), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G2096), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n481), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2435), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2438), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2451), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2454), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n646), .A2(new_n649), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n650), .B2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n641), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n640), .A3(new_n653), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n658), .A3(G14), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g236(.A1(new_n656), .A2(new_n658), .A3(KEYINPUT82), .A4(G14), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  INV_X1    g239(.A(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n666), .B(KEYINPUT17), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n667), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT83), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n669), .A2(new_n666), .A3(new_n667), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT18), .Z(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(new_n669), .A3(new_n673), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(KEYINPUT84), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n681));
  NAND4_X1  g256(.A1(new_n675), .A2(new_n681), .A3(new_n677), .A4(new_n678), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n680), .A2(new_n633), .A3(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n633), .B1(new_n680), .B2(new_n682), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n665), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n687), .A2(G2100), .A3(new_n683), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G227));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n691), .A2(new_n692), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n697), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n694), .A2(new_n696), .A3(new_n698), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n701), .B(new_n702), .C1(new_n700), .C2(new_n699), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT85), .B(G1981), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n703), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1991), .B(G1996), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1986), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(G229));
  OR2_X1    g285(.A1(G16), .A2(G21), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(G286), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G1966), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT30), .B(G28), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n713), .A2(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G5), .A2(G16), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G171), .B2(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G1961), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT31), .B(G11), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n715), .A2(new_n718), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n632), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(G29), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT93), .Z(new_n726));
  AND2_X1   g301(.A1(new_n716), .A2(G32), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n629), .A2(G141), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT91), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n481), .A2(G105), .A3(G2104), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n627), .A2(G129), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT26), .Z(new_n733));
  AND2_X1   g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n729), .A2(new_n730), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n727), .B1(new_n735), .B2(G29), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT27), .B(G1996), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n716), .B1(new_n743), .B2(G34), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(KEYINPUT89), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(G34), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(KEYINPUT89), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI22_X1  g323(.A1(new_n487), .A2(new_n716), .B1(KEYINPUT90), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(KEYINPUT90), .B2(new_n748), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2084), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  NOR2_X1   g327(.A1(G164), .A2(new_n716), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G27), .B2(new_n716), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n716), .A2(G26), .ZN(new_n756));
  OAI221_X1 g331(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n473), .C2(G116), .ZN(new_n757));
  INV_X1    g332(.A(G128), .ZN(new_n758));
  INV_X1    g333(.A(G140), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n757), .B1(new_n498), .B2(new_n758), .C1(new_n759), .C2(new_n501), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n756), .B1(new_n760), .B2(G29), .ZN(new_n761));
  MUX2_X1   g336(.A(new_n756), .B(new_n761), .S(KEYINPUT28), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2067), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n737), .A2(new_n740), .A3(new_n738), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n742), .A2(new_n755), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n716), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n716), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT94), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT29), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AOI21_X1  g346(.A(G2090), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n770), .A2(new_n771), .A3(G2090), .ZN(new_n773));
  NAND2_X1  g348(.A1(G299), .A2(G16), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n712), .A2(KEYINPUT23), .A3(G20), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT23), .ZN(new_n776));
  INV_X1    g351(.A(G20), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G16), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n774), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1956), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n754), .A2(new_n752), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n720), .A2(G1961), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n773), .A2(new_n783), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n726), .A2(new_n765), .A3(new_n772), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT87), .ZN(new_n786));
  INV_X1    g361(.A(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G16), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(G16), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G303), .B2(G16), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n788), .B1(new_n790), .B2(new_n786), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1971), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(new_n588), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G16), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT33), .B(G1976), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n712), .A2(G6), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n712), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT86), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT32), .B(G1981), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n803), .B2(new_n804), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n798), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT34), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n798), .A2(new_n807), .A3(new_n811), .A4(new_n808), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n810), .A2(KEYINPUT88), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n814));
  INV_X1    g389(.A(G290), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G16), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G16), .B2(G24), .ZN(new_n817));
  INV_X1    g392(.A(G1986), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI221_X1 g395(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n473), .C2(G107), .ZN(new_n821));
  INV_X1    g396(.A(G119), .ZN(new_n822));
  INV_X1    g397(.A(G131), .ZN(new_n823));
  OAI221_X1 g398(.A(new_n821), .B1(new_n498), .B2(new_n822), .C1(new_n823), .C2(new_n501), .ZN(new_n824));
  MUX2_X1   g399(.A(G25), .B(new_n824), .S(G29), .Z(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT35), .B(G1991), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n825), .B(new_n826), .Z(new_n827));
  NAND4_X1  g402(.A1(new_n813), .A2(new_n814), .A3(new_n820), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n810), .A2(KEYINPUT88), .A3(new_n827), .A4(new_n812), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT36), .B1(new_n829), .B2(new_n819), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT25), .Z(new_n833));
  INV_X1    g408(.A(G139), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n465), .A2(new_n467), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n835), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n836));
  OAI221_X1 g411(.A(new_n833), .B1(new_n834), .B2(new_n501), .C1(new_n473), .C2(new_n836), .ZN(new_n837));
  MUX2_X1   g412(.A(G33), .B(new_n837), .S(G29), .Z(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(G2072), .Z(new_n839));
  AND3_X1   g414(.A1(new_n785), .A2(new_n831), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT95), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n614), .A2(G16), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(G4), .B2(G16), .ZN(new_n843));
  INV_X1    g418(.A(G1348), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n712), .A2(G19), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n570), .B2(new_n712), .ZN(new_n848));
  INV_X1    g423(.A(G1341), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n840), .A2(new_n841), .A3(new_n846), .A4(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n785), .A2(new_n831), .A3(new_n850), .A4(new_n839), .ZN(new_n852));
  OAI21_X1  g427(.A(KEYINPUT95), .B1(new_n852), .B2(new_n845), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(G311));
  NAND3_X1  g429(.A1(new_n840), .A2(new_n846), .A3(new_n850), .ZN(G150));
  NAND2_X1  g430(.A1(new_n531), .A2(G55), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n534), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT97), .B(G93), .ZN(new_n858));
  OAI221_X1 g433(.A(new_n856), .B1(new_n555), .B2(new_n857), .C1(new_n539), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NOR2_X1   g436(.A1(new_n613), .A2(new_n621), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT39), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n569), .B(new_n859), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n861), .B1(new_n867), .B2(G860), .ZN(G145));
  INV_X1    g443(.A(new_n504), .ZN(new_n869));
  OAI211_X1 g444(.A(G126), .B(new_n467), .C1(new_n490), .C2(new_n491), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n505), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n871), .B2(G2105), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n511), .A2(KEYINPUT98), .A3(new_n516), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT98), .B1(new_n511), .B2(new_n516), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n636), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT91), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n728), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n734), .A2(new_n730), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI221_X1 g456(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n473), .C2(G118), .ZN(new_n882));
  INV_X1    g457(.A(G130), .ZN(new_n883));
  INV_X1    g458(.A(G142), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n882), .B1(new_n498), .B2(new_n883), .C1(new_n884), .C2(new_n501), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n824), .B(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n881), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n837), .B(new_n760), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n632), .A2(G160), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n632), .A2(G160), .ZN(new_n891));
  AOI21_X1  g466(.A(G162), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n893), .A2(new_n889), .A3(new_n502), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n888), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n888), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n502), .B1(new_n893), .B2(new_n889), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n890), .A2(G162), .A3(new_n891), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n887), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n887), .B1(new_n899), .B2(new_n895), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n877), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n895), .A2(new_n899), .ZN(new_n904));
  INV_X1    g479(.A(new_n887), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n887), .A2(new_n895), .A3(new_n899), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n876), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n903), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n902), .A2(KEYINPUT99), .A3(new_n908), .A4(new_n903), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT100), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(KEYINPUT40), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(G395));
  NOR2_X1   g496(.A1(new_n859), .A2(G868), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n924));
  NAND2_X1  g499(.A1(G166), .A2(new_n588), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n794), .A2(G303), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n815), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(G290), .A2(new_n925), .A3(new_n926), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n800), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n800), .B1(new_n928), .B2(new_n929), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n924), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n929), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G305), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(KEYINPUT102), .A3(new_n930), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT42), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n930), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(KEYINPUT42), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n866), .B(KEYINPUT101), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(new_n624), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n613), .B(G299), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT41), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n943), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n947), .B2(new_n942), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n923), .B1(new_n940), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n940), .A2(new_n948), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n949), .B(new_n950), .Z(new_n951));
  AOI21_X1  g526(.A(new_n922), .B1(new_n951), .B2(G868), .ZN(G295));
  AOI21_X1  g527(.A(new_n922), .B1(new_n951), .B2(G868), .ZN(G331));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n954));
  XNOR2_X1  g529(.A(G286), .B(G171), .ZN(new_n955));
  INV_X1    g530(.A(new_n866), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(G286), .B(G301), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT105), .B1(new_n958), .B2(new_n866), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n955), .A2(new_n960), .A3(new_n956), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(KEYINPUT104), .A3(new_n866), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n957), .A2(new_n959), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n958), .B(new_n956), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n963), .A2(new_n944), .B1(new_n964), .B2(new_n947), .ZN(new_n965));
  AOI21_X1  g540(.A(G37), .B1(new_n965), .B2(new_n937), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  OAI22_X1  g542(.A1(new_n963), .A2(new_n943), .B1(new_n945), .B2(new_n964), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n933), .A2(new_n936), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT106), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n965), .A2(new_n937), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n903), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n965), .A2(new_n937), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT43), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n966), .A2(new_n977), .A3(new_n967), .A4(new_n970), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n967), .B1(new_n974), .B2(new_n975), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n966), .A2(KEYINPUT43), .A3(new_n970), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  MUX2_X1   g557(.A(new_n979), .B(new_n982), .S(KEYINPUT44), .Z(G397));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT45), .B1(new_n875), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(G40), .B(new_n475), .C1(new_n485), .C2(new_n486), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1996), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n881), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n735), .A2(G1996), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n760), .B(G2067), .Z(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n824), .A2(new_n826), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n826), .B2(new_n824), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n818), .B2(new_n815), .ZN(new_n999));
  NOR2_X1   g574(.A1(G290), .A2(G1986), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n989), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT121), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n985), .B2(new_n986), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT98), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT4), .B(G138), .C1(new_n513), .C2(new_n514), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n492), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT4), .B1(new_n510), .B2(new_n835), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n511), .A2(KEYINPUT98), .A3(new_n516), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n1011), .B2(new_n872), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT112), .B(new_n987), .C1(new_n1012), .C2(KEYINPUT45), .ZN(new_n1013));
  INV_X1    g588(.A(new_n517), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1384), .B1(new_n872), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT45), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G2078), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1004), .A2(new_n1013), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n984), .B1(new_n508), .B2(new_n517), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT50), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n875), .A2(new_n984), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n1024));
  OAI211_X1 g599(.A(new_n987), .B(new_n1022), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1961), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1019), .A2(new_n1020), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1020), .B1(new_n1019), .B2(new_n1027), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n875), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1021), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1030), .A2(new_n1032), .A3(new_n752), .A4(new_n987), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1033), .A2(KEYINPUT120), .A3(new_n1017), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT120), .B1(new_n1033), .B2(new_n1017), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1028), .A2(new_n1029), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1002), .B1(new_n1037), .B2(G301), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1019), .A2(new_n1027), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT119), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1035), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1033), .A2(KEYINPUT120), .A3(new_n1017), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1019), .A2(new_n1020), .A3(new_n1027), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1046));
  INV_X1    g621(.A(new_n985), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1047), .A2(new_n987), .A3(new_n1030), .A4(new_n1018), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1027), .B(new_n1048), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1049), .A2(G171), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1038), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(G171), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT122), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1040), .A2(G301), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1049), .A2(new_n1057), .A3(G171), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1055), .A2(KEYINPUT54), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1012), .A2(new_n987), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n794), .A2(G1976), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(G8), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(KEYINPUT109), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT110), .B(G1976), .ZN(new_n1067));
  NAND3_X1  g642(.A1(G288), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1060), .A2(G8), .A3(new_n1061), .A4(new_n1064), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G305), .A2(G1981), .ZN(new_n1071));
  INV_X1    g646(.A(G1981), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n592), .A2(new_n1072), .A3(new_n593), .A4(new_n595), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT49), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1071), .A2(KEYINPUT49), .A3(new_n1073), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1076), .A2(G8), .A3(new_n1060), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1070), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G8), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n1081));
  NAND4_X1  g656(.A1(G303), .A2(KEYINPUT108), .A3(new_n1081), .A4(G8), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G166), .A2(new_n1080), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT108), .B(KEYINPUT55), .Z(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1024), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n986), .B1(new_n1012), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G2090), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n1022), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1030), .A2(new_n987), .A3(new_n1032), .ZN(new_n1090));
  INV_X1    g665(.A(G1971), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1080), .B(new_n1085), .C1(new_n1089), .C2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1079), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n986), .B1(new_n1096), .B2(new_n1015), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1097), .A3(new_n1088), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT111), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1092), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G8), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1099), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1085), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1094), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1025), .A2(G2084), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1004), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n714), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1080), .B1(new_n1108), .B2(G168), .ZN(new_n1109));
  NAND2_X1  g684(.A1(G286), .A2(G8), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT51), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1108), .A2(new_n1080), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G286), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1113), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1110), .B(new_n1117), .C1(new_n1108), .C2(new_n1080), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1059), .A2(new_n1105), .A3(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1053), .A2(new_n1120), .A3(KEYINPUT123), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT123), .B1(new_n1053), .B2(new_n1120), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1123));
  INV_X1    g698(.A(G1956), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1030), .A2(new_n1032), .A3(new_n987), .A4(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1125), .A2(KEYINPUT115), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT115), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n552), .A2(G91), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT114), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(new_n582), .A4(new_n578), .ZN(new_n1132));
  NAND2_X1  g707(.A1(G299), .A2(KEYINPUT114), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1132), .A2(new_n1133), .A3(KEYINPUT57), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT57), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1128), .A2(new_n1129), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1025), .A2(new_n844), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(G2067), .B2(new_n1060), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n614), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1136), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  OR2_X1    g719(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1145));
  NAND2_X1  g720(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1060), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(G1996), .B2(new_n1090), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n570), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1125), .A2(KEYINPUT117), .A3(new_n1136), .A4(new_n1127), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT61), .B1(new_n1137), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1136), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1158));
  OR3_X1    g733(.A1(new_n1143), .A2(new_n1158), .A3(KEYINPUT61), .ZN(new_n1159));
  AOI211_X1 g734(.A(new_n1151), .B(new_n1152), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n613), .B1(new_n1139), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1139), .A2(new_n1161), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1144), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1121), .A2(new_n1122), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1114), .A2(new_n1116), .A3(new_n1168), .A4(new_n1118), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1167), .A2(new_n1105), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1119), .A2(KEYINPUT62), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1167), .A2(KEYINPUT124), .A3(new_n1105), .A4(new_n1169), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(G8), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1079), .A2(new_n1177), .A3(new_n1085), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1060), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1180));
  OR3_X1    g755(.A1(new_n1180), .A2(G1976), .A3(G288), .ZN(new_n1181));
  AOI211_X1 g756(.A(new_n1080), .B(new_n1179), .C1(new_n1181), .C2(new_n1073), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT113), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1108), .A2(new_n1080), .A3(G286), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1104), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1094), .A2(new_n1103), .A3(KEYINPUT113), .A4(new_n1184), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1177), .B2(new_n1085), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1094), .A2(new_n1190), .A3(new_n1184), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1178), .B(new_n1182), .C1(new_n1189), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1175), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1001), .B1(new_n1166), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n989), .A2(new_n1000), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT48), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n998), .B2(new_n988), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n989), .B1(new_n994), .B2(new_n735), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT46), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1199), .B1(new_n988), .B2(G1996), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n989), .A2(KEYINPUT46), .A3(new_n990), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT47), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n996), .B(KEYINPUT125), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n995), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1205), .B1(G2067), .B2(new_n760), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n989), .ZN(new_n1207));
  AND3_X1   g782(.A1(new_n1197), .A2(new_n1203), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1194), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g784(.A1(G229), .A2(new_n461), .ZN(new_n1211));
  NAND3_X1  g785(.A1(new_n689), .A2(new_n663), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n1214), .B1(new_n911), .B2(new_n912), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1216));
  NAND3_X1  g790(.A1(new_n979), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n1218));
  XNOR2_X1  g792(.A(new_n1217), .B(new_n1218), .ZN(G308));
  XNOR2_X1  g793(.A(new_n1217), .B(KEYINPUT127), .ZN(G225));
endmodule


