//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n205), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT14), .B(G29gat), .Z(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G36gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n202), .A2(new_n203), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n204), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n211), .B2(KEYINPUT93), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(KEYINPUT93), .B2(new_n211), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(G1gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT95), .ZN(new_n220));
  INV_X1    g019(.A(G8gat), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n216), .A2(G1gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(KEYINPUT95), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT94), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n225), .A3(new_n218), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n226), .B(G8gat), .C1(new_n225), .C2(new_n218), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n215), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n214), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n230), .A2(new_n231), .B1(new_n228), .B2(new_n213), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(KEYINPUT18), .A3(new_n233), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n213), .B(new_n228), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT96), .B(KEYINPUT13), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(new_n233), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT97), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G197gat), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT11), .B(G169gat), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT12), .Z(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT92), .Z(new_n249));
  NAND3_X1  g048(.A1(new_n242), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n248), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n236), .A2(new_n237), .A3(new_n241), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n243), .B1(new_n242), .B2(new_n249), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G225gat), .A2(G233gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(G155gat), .A2(G162gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT2), .ZN(new_n258));
  INV_X1    g057(.A(G141gat), .ZN(new_n259));
  INV_X1    g058(.A(G148gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G141gat), .A2(G148gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT80), .ZN(new_n264));
  AND2_X1   g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G155gat), .ZN(new_n268));
  INV_X1    g067(.A(G162gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT80), .A3(new_n257), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n263), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n257), .B1(new_n270), .B2(KEYINPUT2), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n274));
  AND2_X1   g073(.A1(G141gat), .A2(G148gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n261), .A2(KEYINPUT81), .A3(new_n262), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n281));
  INV_X1    g080(.A(G127gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G134gat), .ZN(new_n283));
  INV_X1    g082(.A(G134gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(G127gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT68), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(G127gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n282), .A2(G134gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G113gat), .ZN(new_n291));
  INV_X1    g090(.A(G120gat), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G113gat), .A2(G120gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n286), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n287), .A2(new_n288), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n297), .A2(KEYINPUT68), .A3(new_n294), .A4(new_n293), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n272), .A2(new_n279), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n272), .A2(new_n279), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n296), .A2(new_n298), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n303), .B2(new_n305), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n256), .B(new_n302), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n308), .A2(KEYINPUT5), .ZN(new_n309));
  XNOR2_X1  g108(.A(G1gat), .B(G29gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT0), .ZN(new_n311));
  XNOR2_X1  g110(.A(G57gat), .B(G85gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(KEYINPUT82), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT4), .B1(new_n299), .B2(new_n280), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT82), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n256), .A4(new_n302), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n305), .B(new_n280), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT5), .B1(new_n321), .B2(new_n256), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT83), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT83), .ZN(new_n325));
  AOI211_X1 g124(.A(new_n325), .B(new_n322), .C1(new_n314), .C2(new_n319), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n309), .B(new_n313), .C1(new_n324), .C2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n309), .B1(new_n324), .B2(new_n326), .ZN(new_n330));
  INV_X1    g129(.A(new_n313), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT6), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n327), .B2(new_n328), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n332), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n338));
  INV_X1    g137(.A(G226gat), .ZN(new_n339));
  INV_X1    g138(.A(G233gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343));
  AND2_X1   g142(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(G190gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n346), .A2(KEYINPUT64), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT64), .B1(new_n346), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT65), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n345), .B(KEYINPUT65), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT23), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(G169gat), .B2(G176gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(new_n353), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n355), .A2(new_n358), .A3(new_n357), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT27), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G183gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT66), .ZN(new_n371));
  INV_X1    g170(.A(G190gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G183gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT27), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT66), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n368), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT27), .B(G183gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n368), .A2(G190gat), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT67), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT26), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n354), .B2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n358), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n388), .B1(new_n384), .B2(new_n354), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n387), .A2(new_n389), .B1(G183gat), .B2(G190gat), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n361), .A2(new_n367), .B1(new_n382), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n342), .B1(new_n391), .B2(KEYINPUT29), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT75), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n391), .B2(new_n342), .ZN(new_n394));
  NAND3_X1  g193(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(G183gat), .B2(G190gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT64), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n363), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n346), .A2(KEYINPUT64), .A3(new_n347), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n360), .B1(new_n400), .B2(KEYINPUT65), .ZN(new_n401));
  INV_X1    g200(.A(new_n353), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n367), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n382), .A2(new_n390), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT75), .A3(new_n341), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n392), .A2(new_n394), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G211gat), .A2(G218gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT22), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT74), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(KEYINPUT74), .A3(new_n409), .ZN(new_n413));
  XNOR2_X1  g212(.A(G197gat), .B(G204gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G211gat), .ZN(new_n416));
  INV_X1    g215(.A(G218gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n408), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n408), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n412), .A2(new_n420), .A3(new_n414), .A4(new_n413), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT76), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n392), .A2(KEYINPUT77), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT77), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(new_n342), .C1(new_n391), .C2(KEYINPUT29), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n405), .A2(new_n341), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n427), .A2(new_n422), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n407), .A2(KEYINPUT76), .A3(new_n423), .ZN(new_n432));
  XOR2_X1   g231(.A(G8gat), .B(G36gat), .Z(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT78), .ZN(new_n434));
  XNOR2_X1  g233(.A(G64gat), .B(G92gat), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n434), .B(new_n435), .Z(new_n436));
  NAND4_X1  g235(.A1(new_n426), .A2(new_n431), .A3(new_n432), .A4(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n338), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n431), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT76), .B1(new_n407), .B2(new_n423), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n442), .A2(KEYINPUT79), .A3(KEYINPUT30), .A4(new_n436), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n437), .A2(new_n438), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n431), .A3(new_n432), .ZN(new_n446));
  INV_X1    g245(.A(new_n436), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n335), .A2(new_n337), .A3(new_n444), .A4(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT29), .B1(new_n419), .B2(new_n421), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n280), .B1(new_n451), .B2(KEYINPUT3), .ZN(new_n452));
  INV_X1    g251(.A(G228gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(new_n340), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT29), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n301), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n423), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n452), .A2(new_n457), .A3(KEYINPUT87), .A4(new_n454), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n452), .A2(new_n457), .ZN(new_n465));
  INV_X1    g264(.A(new_n454), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT86), .B(new_n454), .C1(new_n452), .C2(new_n457), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(G22gat), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G78gat), .B(G106gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n471), .B(KEYINPUT85), .Z(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n465), .A2(new_n466), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT86), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n465), .A2(new_n464), .A3(new_n466), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G22gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n462), .A3(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n470), .A2(new_n473), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n473), .B1(new_n470), .B2(new_n479), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT31), .B(G50gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n463), .A2(new_n469), .A3(G22gat), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n478), .B1(new_n477), .B2(new_n462), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n472), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n473), .A3(new_n479), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n482), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n450), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n359), .B1(new_n350), .B2(new_n351), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n492), .A2(new_n353), .B1(new_n366), .B2(new_n365), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n372), .B(new_n371), .C1(new_n378), .C2(KEYINPUT66), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n380), .B1(new_n494), .B2(new_n368), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n387), .A2(new_n389), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n346), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT69), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n493), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT69), .B1(new_n403), .B2(new_n404), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n299), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G227gat), .A2(G233gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n499), .B1(new_n493), .B2(new_n498), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n305), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT34), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n502), .A2(new_n503), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n403), .A2(KEYINPUT69), .A3(new_n404), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n305), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n501), .A2(new_n299), .ZN(new_n511));
  INV_X1    g310(.A(new_n503), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n503), .B1(new_n502), .B2(new_n505), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT32), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT70), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n512), .B1(new_n510), .B2(new_n511), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT70), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT32), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G43gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(G71gat), .B(G99gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n518), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n524), .A2(new_n525), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n519), .A2(KEYINPUT32), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n519), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n515), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n526), .A3(new_n521), .ZN(new_n535));
  INV_X1    g334(.A(new_n515), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n535), .A2(new_n536), .A3(new_n531), .A4(new_n532), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(KEYINPUT73), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT36), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n540), .B(new_n515), .C1(new_n527), .C2(new_n533), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n534), .A2(KEYINPUT36), .A3(new_n537), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n444), .A2(new_n449), .A3(KEYINPUT88), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT88), .B1(new_n444), .B2(new_n449), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n305), .B1(KEYINPUT3), .B2(new_n280), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n315), .A2(new_n316), .B1(new_n547), .B2(new_n301), .ZN(new_n548));
  OR3_X1    g347(.A1(new_n548), .A2(KEYINPUT39), .A3(new_n256), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n256), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n321), .A2(new_n256), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT39), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n549), .B(new_n313), .C1(new_n550), .C2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(KEYINPUT89), .A2(KEYINPUT40), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n332), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n545), .A2(new_n546), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n483), .B1(new_n480), .B2(new_n481), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n487), .A2(new_n482), .A3(new_n488), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n318), .B1(new_n548), .B2(new_n256), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n308), .A2(KEYINPUT82), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n323), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n325), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n320), .A2(KEYINPUT83), .A3(new_n323), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n566), .A2(KEYINPUT84), .A3(new_n309), .A4(new_n313), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n567), .A2(new_n334), .B1(new_n330), .B2(new_n331), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT6), .B1(new_n329), .B2(new_n332), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n437), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT90), .B(KEYINPUT38), .Z(new_n571));
  OAI21_X1  g370(.A(new_n447), .B1(new_n446), .B2(KEYINPUT37), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n442), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n571), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n436), .B1(new_n442), .B2(new_n573), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n573), .B1(new_n407), .B2(new_n422), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n427), .A2(new_n423), .A3(new_n429), .A4(new_n430), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n571), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(KEYINPUT91), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n447), .B(new_n579), .C1(new_n446), .C2(KEYINPUT37), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT91), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n575), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n560), .B1(new_n570), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n491), .B(new_n544), .C1(new_n557), .C2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n560), .A2(new_n534), .A3(new_n537), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT35), .B1(new_n587), .B2(new_n450), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n545), .A2(new_n546), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n538), .A2(new_n541), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n568), .A2(new_n569), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT35), .B1(new_n558), .B2(new_n559), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n588), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n255), .B1(new_n586), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n591), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT102), .B(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT7), .ZN(new_n602));
  INV_X1    g401(.A(G99gat), .ZN(new_n603));
  INV_X1    g402(.A(G106gat), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT8), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G99gat), .B(G106gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n215), .A2(new_n231), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n213), .A2(new_n608), .B1(KEYINPUT41), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G190gat), .B(G218gat), .Z(new_n614));
  NOR2_X1   g413(.A1(new_n611), .A2(KEYINPUT41), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G134gat), .B(G162gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n613), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G57gat), .B(G64gat), .Z(new_n623));
  INV_X1    g422(.A(KEYINPUT9), .ZN(new_n624));
  INV_X1    g423(.A(G71gat), .ZN(new_n625));
  INV_X1    g424(.A(G78gat), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G71gat), .B(G78gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n623), .A2(new_n629), .A3(new_n627), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT101), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n228), .B1(new_n635), .B2(KEYINPUT21), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT98), .B(KEYINPUT21), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G127gat), .B(G155gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n636), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT99), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT100), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G183gat), .B(G211gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n641), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n622), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n634), .A2(new_n609), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n608), .B(new_n633), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(G230gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n340), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n655), .A2(new_n657), .A3(new_n340), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  OR2_X1    g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n664), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n597), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g469(.A1(new_n595), .A2(new_n668), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n221), .B1(new_n672), .B2(new_n589), .ZN(new_n673));
  INV_X1    g472(.A(new_n589), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT16), .B(G8gat), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT42), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(KEYINPUT42), .B2(new_n676), .ZN(G1325gat));
  NAND2_X1  g477(.A1(new_n595), .A2(new_n590), .ZN(new_n679));
  OR4_X1    g478(.A1(G15gat), .A2(new_n679), .A3(new_n652), .A4(new_n667), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n544), .A2(KEYINPUT105), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n542), .A2(new_n682), .A3(new_n543), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G15gat), .B1(new_n671), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(new_n685), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n560), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT106), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n667), .A2(new_n651), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n621), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n597), .A2(new_n205), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT45), .Z(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n586), .A2(new_n594), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(new_n621), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n593), .A2(new_n589), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT35), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n444), .A2(new_n449), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(new_n569), .A3(new_n568), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n534), .A2(new_n537), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n490), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n701), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n699), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n588), .B(KEYINPUT108), .C1(new_n589), .C2(new_n593), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n542), .A2(new_n682), .A3(new_n543), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n682), .B1(new_n542), .B2(new_n543), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n491), .B1(new_n557), .B2(new_n585), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n546), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n444), .A2(new_n449), .A3(KEYINPUT88), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n716), .A2(new_n332), .A3(new_n717), .A4(new_n555), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n335), .A2(new_n337), .B1(new_n442), .B2(new_n436), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n575), .A2(new_n580), .A3(new_n583), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n490), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n684), .A2(new_n722), .A3(KEYINPUT107), .A4(new_n491), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n709), .A2(new_n715), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n622), .A2(KEYINPUT44), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n698), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n255), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n691), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n205), .B1(new_n729), .B2(new_n596), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n695), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT109), .Z(G1328gat));
  INV_X1    g531(.A(new_n729), .ZN(new_n733));
  OAI21_X1  g532(.A(G36gat), .B1(new_n733), .B2(new_n674), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735));
  AOI21_X1  g534(.A(G36gat), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n595), .A2(new_n589), .A3(new_n693), .A4(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n737), .B(new_n739), .Z(new_n740));
  NAND2_X1  g539(.A1(new_n734), .A2(new_n740), .ZN(G1329gat));
  NOR2_X1   g540(.A1(new_n733), .A2(new_n684), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743));
  OAI21_X1  g542(.A(G43gat), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n743), .B2(new_n742), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n679), .A2(G43gat), .A3(new_n692), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT47), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n713), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n746), .B1(new_n749), .B2(G43gat), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n745), .A2(new_n748), .B1(KEYINPUT47), .B2(new_n750), .ZN(G1330gat));
  INV_X1    g550(.A(G50gat), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n729), .B2(new_n490), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n490), .A2(new_n752), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n693), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n754), .B2(new_n755), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n753), .B1(new_n595), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g558(.A(new_n667), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n727), .A2(new_n652), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n724), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n596), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g564(.A1(new_n762), .A2(new_n674), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  AND2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n766), .B2(new_n767), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n762), .B2(new_n684), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n590), .A2(new_n625), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n762), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g573(.A1(new_n762), .A2(new_n560), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(new_n626), .ZN(G1335gat));
  NOR3_X1   g575(.A1(new_n727), .A2(new_n651), .A3(new_n760), .ZN(new_n777));
  INV_X1    g576(.A(new_n725), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n713), .A2(new_n714), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n779), .A2(KEYINPUT107), .B1(new_n707), .B2(new_n708), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(new_n780), .B2(new_n715), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n777), .B1(new_n781), .B2(new_n698), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n591), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n727), .A2(new_n651), .A3(new_n622), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n724), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n724), .A2(KEYINPUT51), .A3(new_n784), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n596), .A2(new_n598), .A3(new_n667), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n783), .A2(new_n598), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n791), .B(KEYINPUT113), .Z(G1336gat));
  OAI21_X1  g591(.A(G92gat), .B1(new_n782), .B2(new_n674), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n787), .A2(KEYINPUT114), .A3(new_n788), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n785), .A2(new_n795), .A3(new_n786), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n589), .A2(new_n599), .A3(new_n667), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT52), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n793), .B(new_n801), .C1(new_n789), .C2(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n782), .B2(new_n684), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n590), .A2(new_n603), .A3(new_n667), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n789), .B2(new_n805), .ZN(G1338gat));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n807));
  INV_X1    g606(.A(new_n777), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n726), .A2(new_n560), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n809), .B2(new_n604), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n560), .A2(new_n760), .A3(G106gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n796), .A3(new_n811), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n490), .B(new_n777), .C1(new_n781), .C2(new_n698), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n810), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT53), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  INV_X1    g616(.A(new_n811), .ZN(new_n818));
  OAI221_X1 g617(.A(new_n817), .B1(new_n809), .B2(new_n604), .C1(new_n789), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n816), .A2(KEYINPUT116), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1339gat));
  NOR2_X1   g623(.A1(new_n232), .A2(new_n233), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n238), .A2(new_n240), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n247), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n252), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n621), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n659), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n656), .A2(new_n658), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n664), .B1(new_n659), .B2(new_n831), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n666), .A4(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n666), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n830), .A2(new_n841), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n841), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT118), .B1(new_n846), .B2(new_n829), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n828), .A2(new_n667), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n255), .B2(new_n846), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n622), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n651), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n668), .A2(new_n255), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n589), .A2(new_n591), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n855), .A2(new_n587), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n727), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n590), .A2(new_n560), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n856), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n255), .A2(new_n291), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(G1340gat));
  AOI21_X1  g664(.A(G120gat), .B1(new_n858), .B2(new_n667), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n760), .A2(new_n292), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n863), .B2(new_n867), .ZN(G1341gat));
  INV_X1    g667(.A(new_n651), .ZN(new_n869));
  OAI21_X1  g668(.A(G127gat), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n858), .A2(new_n282), .A3(new_n651), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  OAI21_X1  g671(.A(G134gat), .B1(new_n862), .B2(new_n622), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n284), .A3(new_n621), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT119), .B1(new_n874), .B2(KEYINPUT56), .ZN(new_n876));
  OAI221_X1 g675(.A(new_n873), .B1(KEYINPUT56), .B2(new_n874), .C1(new_n875), .C2(new_n876), .ZN(G1343gat));
  OAI21_X1  g676(.A(new_n849), .B1(new_n255), .B2(new_n843), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n622), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n651), .B1(new_n848), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n490), .B1(new_n880), .B2(new_n854), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n713), .A2(new_n857), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n884), .B(new_n490), .C1(new_n852), .C2(new_n854), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886), .B2(new_n255), .ZN(new_n887));
  NOR4_X1   g686(.A1(new_n855), .A2(new_n560), .A3(new_n713), .A4(new_n857), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n255), .A2(G141gat), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n888), .A2(new_n889), .B1(new_n890), .B2(KEYINPUT58), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n890), .A2(KEYINPUT58), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n892), .B(new_n893), .Z(G1344gat));
  NOR3_X1   g693(.A1(new_n855), .A2(new_n560), .A3(new_n857), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n760), .A2(G148gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n684), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n897), .B(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n879), .B1(new_n829), .B2(new_n843), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n869), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n853), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n560), .A2(KEYINPUT57), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n490), .B1(new_n852), .B2(new_n854), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n903), .A2(new_n904), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n883), .A2(KEYINPUT122), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n883), .A2(KEYINPUT122), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n906), .A2(new_n667), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n900), .B1(new_n909), .B2(G148gat), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n886), .A2(new_n760), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n900), .A2(G148gat), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n899), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n899), .B(KEYINPUT123), .C1(new_n910), .C2(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1345gat));
  OAI21_X1  g717(.A(G155gat), .B1(new_n886), .B2(new_n869), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n888), .A2(new_n268), .A3(new_n651), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  OR2_X1    g720(.A1(new_n886), .A2(new_n622), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n269), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n888), .A2(new_n269), .A3(new_n621), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n674), .A2(new_n596), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n861), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(G169gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n929), .A2(new_n930), .A3(new_n255), .ZN(new_n931));
  NOR4_X1   g730(.A1(new_n855), .A2(new_n596), .A3(new_n674), .A4(new_n587), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n727), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n931), .A2(new_n933), .ZN(G1348gat));
  OAI21_X1  g733(.A(G176gat), .B1(new_n929), .B2(new_n760), .ZN(new_n935));
  INV_X1    g734(.A(G176gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n932), .A2(new_n936), .A3(new_n667), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n929), .B2(new_n869), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n932), .A2(new_n651), .A3(new_n378), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g740(.A(KEYINPUT125), .B(KEYINPUT60), .Z(new_n942));
  XNOR2_X1  g741(.A(new_n941), .B(new_n942), .ZN(G1350gat));
  NAND3_X1  g742(.A1(new_n932), .A2(new_n372), .A3(new_n621), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n861), .A2(new_n621), .A3(new_n928), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n945), .A2(new_n946), .A3(G190gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n945), .B2(G190gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT126), .ZN(G1351gat));
  NAND2_X1  g749(.A1(new_n684), .A2(new_n928), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n905), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G197gat), .B1(new_n952), .B2(new_n727), .ZN(new_n953));
  INV_X1    g752(.A(new_n951), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n906), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n727), .A2(G197gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1352gat));
  INV_X1    g756(.A(G204gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n952), .A2(new_n958), .A3(new_n667), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n906), .A2(new_n667), .A3(new_n954), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n960), .B(new_n961), .C1(new_n958), .C2(new_n962), .ZN(G1353gat));
  NAND3_X1  g762(.A1(new_n952), .A2(new_n416), .A3(new_n651), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n955), .A2(new_n651), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  AOI21_X1  g767(.A(G218gat), .B1(new_n952), .B2(new_n621), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n622), .A2(new_n417), .ZN(new_n973));
  AOI22_X1  g772(.A1(new_n971), .A2(new_n972), .B1(new_n955), .B2(new_n973), .ZN(G1355gat));
endmodule


