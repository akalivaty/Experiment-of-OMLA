//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0002(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT65), .ZN(new_n205));
  INV_X1    g0005(.A(G13), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G116), .A2(G270), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT66), .B(G77), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT67), .B(G244), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n213), .B(new_n226), .C1(G68), .C2(G238), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT69), .ZN(new_n228));
  OAI22_X1  g0028(.A1(new_n227), .A2(new_n205), .B1(new_n228), .B2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n210), .B(new_n231), .C1(new_n234), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT70), .B(G250), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n242), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  INV_X1    g0048(.A(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G68), .B(G77), .Z(new_n253));
  XNOR2_X1  g0053(.A(G50), .B(G58), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n253), .B(new_n254), .Z(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G223), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n212), .A2(G1698), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n262), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G87), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n259), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n259), .A2(G232), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G179), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NOR4_X1   g0074(.A1(new_n268), .A2(new_n271), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n266), .A2(new_n267), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n271), .ZN(new_n279));
  INV_X1    g0079(.A(new_n274), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n275), .B1(new_n281), .B2(G169), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT16), .ZN(new_n283));
  INV_X1    g0083(.A(G68), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n257), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n233), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT7), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n233), .A4(new_n287), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n284), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G58), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n284), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G58), .A2(G68), .ZN(new_n295));
  OAI21_X1  g0095(.A(G20), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G159), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n283), .B1(new_n292), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT80), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n232), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n290), .A2(new_n291), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n299), .B1(new_n306), .B2(G68), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n305), .B1(new_n307), .B2(KEYINPUT16), .ZN(new_n308));
  OAI211_X1 g0108(.A(KEYINPUT80), .B(new_n283), .C1(new_n292), .C2(new_n299), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n302), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT8), .B(G58), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT72), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT8), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(G58), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT72), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n304), .B1(new_n269), .B2(G20), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n317), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n282), .B1(new_n310), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(KEYINPUT18), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT18), .ZN(new_n324));
  AOI211_X1 g0124(.A(new_n324), .B(new_n282), .C1(new_n310), .C2(new_n321), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n281), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(G190), .B2(new_n281), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n310), .A2(new_n321), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT17), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n310), .A2(KEYINPUT17), .A3(new_n329), .A4(new_n321), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT75), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n311), .A2(KEYINPUT74), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT74), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n293), .A2(KEYINPUT8), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n315), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n336), .A2(new_n339), .A3(new_n297), .ZN(new_n340));
  INV_X1    g0140(.A(new_n223), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n233), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n335), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT15), .B(G87), .Z(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(new_n233), .A3(G33), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n336), .A2(new_n339), .A3(new_n297), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(KEYINPUT75), .C1(new_n233), .C2(new_n341), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n304), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n286), .A2(new_n287), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G238), .A2(G1698), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(new_n351), .C1(new_n239), .C2(G1698), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n264), .A2(new_n265), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT73), .B(G107), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n259), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n274), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n224), .A2(new_n259), .A3(new_n270), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n356), .A2(G190), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n327), .B1(new_n356), .B2(new_n357), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n320), .ZN(new_n361));
  INV_X1    g0161(.A(G77), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n223), .A2(new_n318), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n349), .A2(new_n360), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  AOI211_X1 g0167(.A(new_n363), .B(new_n365), .C1(new_n348), .C2(new_n304), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n356), .A2(new_n357), .ZN(new_n369));
  INV_X1    g0169(.A(G169), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(G179), .B2(new_n369), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n367), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n326), .A2(new_n334), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n233), .B1(new_n295), .B2(new_n211), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(G150), .B2(new_n297), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n233), .A2(G33), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n317), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n318), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n378), .A2(new_n304), .B1(new_n211), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n320), .A2(G50), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT9), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n259), .A2(new_n270), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n280), .B1(new_n384), .B2(new_n212), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT71), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n261), .A2(G222), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n350), .B(new_n387), .C1(new_n260), .C2(new_n261), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n277), .C1(new_n223), .C2(new_n350), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT71), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n280), .B(new_n390), .C1(new_n384), .C2(new_n212), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G200), .ZN(new_n393));
  INV_X1    g0193(.A(G190), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n380), .A2(KEYINPUT9), .A3(new_n381), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n383), .A2(new_n393), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT10), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n395), .A2(KEYINPUT76), .A3(new_n393), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n396), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n382), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n395), .A2(new_n393), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(KEYINPUT76), .C2(KEYINPUT10), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n392), .A2(G179), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n380), .A2(new_n381), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n392), .A2(new_n370), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n400), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(KEYINPUT79), .A2(KEYINPUT14), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n239), .A2(G1698), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n411), .B1(G226), .B2(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G97), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT77), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT77), .B1(new_n412), .B2(new_n413), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n415), .A2(new_n416), .A3(new_n259), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n259), .A2(G238), .A3(new_n270), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT78), .B1(new_n280), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n280), .A2(new_n418), .A3(KEYINPUT78), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT13), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n416), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(new_n277), .A3(new_n414), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT13), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n420), .A4(new_n421), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n410), .B1(new_n428), .B2(G169), .ZN(new_n429));
  INV_X1    g0229(.A(new_n410), .ZN(new_n430));
  AOI211_X1 g0230(.A(new_n370), .B(new_n430), .C1(new_n423), .C2(new_n427), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n423), .A2(new_n427), .A3(G179), .ZN(new_n432));
  NAND2_X1  g0232(.A1(KEYINPUT79), .A2(KEYINPUT14), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n429), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n297), .A2(G50), .B1(G20), .B2(new_n284), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n362), .B2(new_n377), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n304), .ZN(new_n438));
  XOR2_X1   g0238(.A(new_n438), .B(KEYINPUT11), .Z(new_n439));
  NOR2_X1   g0239(.A1(new_n361), .A2(new_n284), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n269), .A2(new_n284), .A3(G13), .A4(G20), .ZN(new_n441));
  XOR2_X1   g0241(.A(new_n441), .B(KEYINPUT12), .Z(new_n442));
  NOR3_X1   g0242(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n435), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n428), .A2(G200), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n443), .C1(new_n394), .C2(new_n428), .ZN(new_n447));
  AND4_X1   g0247(.A1(new_n374), .A2(new_n409), .A3(new_n445), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G1), .ZN(new_n450));
  AND2_X1   g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(G270), .A3(new_n259), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT84), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n450), .B(G274), .C1(new_n452), .C2(new_n451), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n261), .A2(G257), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G264), .A2(G1698), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n459), .C1(new_n264), .C2(new_n265), .ZN(new_n460));
  INV_X1    g0260(.A(G303), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n286), .A2(new_n461), .A3(new_n287), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n277), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n453), .A2(KEYINPUT84), .A3(G270), .A4(new_n259), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n456), .A2(new_n457), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT85), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n463), .A2(new_n457), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT85), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(new_n456), .A4(new_n464), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n466), .A2(KEYINPUT21), .A3(new_n469), .A4(G169), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n465), .A2(new_n272), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n269), .A2(G33), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n318), .A2(new_n473), .A3(new_n232), .A4(new_n303), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n251), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT20), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n251), .A2(G20), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n304), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT86), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n304), .A2(new_n480), .A3(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n483), .B(new_n233), .C1(G33), .C2(new_n217), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT87), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n476), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT87), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n484), .B(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(KEYINPUT20), .A3(new_n479), .A4(new_n481), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n475), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n477), .A2(G1), .A3(new_n206), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n472), .A2(new_n493), .ZN(new_n494));
  AOI211_X1 g0294(.A(new_n491), .B(new_n475), .C1(new_n486), .C2(new_n489), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n466), .A2(G200), .A3(new_n469), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n466), .A2(new_n469), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(new_n394), .ZN(new_n498));
  XOR2_X1   g0298(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n499));
  NAND3_X1  g0299(.A1(new_n466), .A2(G169), .A3(new_n469), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n494), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(KEYINPUT73), .A2(G107), .ZN(new_n503));
  NOR2_X1   g0303(.A1(KEYINPUT73), .A2(G107), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n215), .B(new_n217), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n413), .A2(new_n233), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n505), .A2(KEYINPUT19), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n350), .A2(new_n233), .A3(G68), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT19), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n413), .B2(G20), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n304), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n344), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n379), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n474), .A2(KEYINPUT81), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n474), .A2(KEYINPUT81), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n344), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n512), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G238), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n261), .ZN(new_n520));
  INV_X1    g0320(.A(G244), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G1698), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n522), .C1(new_n264), .C2(new_n265), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n257), .A2(new_n251), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n277), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT82), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n216), .B1(new_n449), .B2(G1), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n269), .A2(new_n273), .A3(G45), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n259), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n259), .B1(new_n523), .B2(new_n525), .ZN(new_n533));
  INV_X1    g0333(.A(new_n531), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT82), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n532), .A2(new_n535), .A3(new_n370), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n518), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n528), .B1(new_n527), .B2(new_n531), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT82), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n272), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT83), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n532), .A2(new_n535), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT83), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n543), .A3(new_n272), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n537), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT23), .B1(new_n249), .B2(G20), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n354), .B2(KEYINPUT23), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n233), .B2(G107), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n547), .A2(new_n233), .B1(new_n549), .B2(new_n524), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n233), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT22), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n350), .A2(KEYINPUT22), .A3(new_n233), .A4(G87), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n550), .A2(KEYINPUT24), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n549), .A2(new_n524), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT23), .B1(new_n503), .B2(new_n504), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n549), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n559), .B2(G20), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n553), .A2(new_n554), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n555), .A2(new_n562), .A3(new_n304), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n515), .A2(G107), .A3(new_n516), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n318), .A2(G107), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n565), .B(KEYINPUT25), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n216), .A2(new_n261), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n218), .A2(G1698), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n264), .C2(new_n265), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G294), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n277), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n453), .A2(G264), .A3(new_n259), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n573), .A2(new_n457), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT89), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n453), .A2(KEYINPUT89), .A3(G264), .A4(new_n259), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n577), .A2(new_n573), .A3(new_n457), .A4(new_n578), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n575), .A2(new_n370), .B1(new_n579), .B2(new_n272), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n567), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n327), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n573), .A2(new_n394), .A3(new_n457), .A4(new_n574), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(new_n564), .A3(new_n566), .A4(new_n563), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n515), .A2(G87), .A3(new_n516), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n512), .A2(new_n514), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n542), .A2(G190), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n532), .A2(new_n535), .A3(G200), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n545), .A2(new_n581), .A3(new_n585), .A4(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n354), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n306), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n297), .A2(G77), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n249), .A2(KEYINPUT6), .A3(G97), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n217), .A2(new_n249), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G97), .A2(G107), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n599), .B2(KEYINPUT6), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G20), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n594), .A2(new_n595), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n304), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n379), .A2(new_n217), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n515), .A2(G97), .A3(new_n516), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n453), .A2(new_n259), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n457), .B1(new_n607), .B2(new_n218), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n216), .B1(new_n286), .B2(new_n287), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT4), .ZN(new_n610));
  OAI21_X1  g0410(.A(G1698), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n483), .ZN(new_n612));
  OAI21_X1  g0412(.A(G244), .B1(new_n264), .B2(new_n265), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(new_n610), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n350), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n611), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n608), .B1(new_n616), .B2(new_n277), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(G169), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n272), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n606), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n277), .ZN(new_n622));
  INV_X1    g0422(.A(new_n608), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G200), .ZN(new_n625));
  INV_X1    g0425(.A(new_n605), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n602), .B2(new_n304), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n617), .A2(G190), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n625), .A2(new_n627), .A3(new_n604), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n502), .A2(new_n592), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n448), .A2(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n408), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n310), .A2(new_n321), .ZN(new_n634));
  INV_X1    g0434(.A(new_n282), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n324), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n322), .A2(KEYINPUT18), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n429), .A2(new_n431), .A3(new_n434), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n443), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n349), .A2(new_n364), .A3(new_n366), .ZN(new_n642));
  INV_X1    g0442(.A(new_n372), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n447), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n639), .B1(new_n646), .B2(new_n334), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n400), .A2(new_n404), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n633), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n606), .A2(new_n619), .A3(new_n620), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(new_n591), .A3(new_n545), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT26), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n533), .A2(new_n534), .ZN(new_n653));
  OR3_X1    g0453(.A1(new_n653), .A2(KEYINPUT90), .A3(G169), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT90), .B1(new_n653), .B2(G169), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n540), .A2(new_n654), .A3(new_n518), .A4(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n653), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G200), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n588), .A2(new_n589), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n656), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(new_n650), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n652), .A2(new_n656), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n581), .A2(KEYINPUT91), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT91), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n567), .A2(new_n666), .A3(new_n580), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n665), .A2(new_n494), .A3(new_n501), .A4(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n621), .A2(new_n629), .A3(new_n585), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n668), .A2(new_n661), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n448), .B1(new_n664), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n649), .A2(new_n671), .ZN(G369));
  NOR3_X1   g0472(.A1(new_n206), .A2(G1), .A3(G20), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT27), .ZN(new_n674));
  OR3_X1    g0474(.A1(new_n673), .A2(KEYINPUT92), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G213), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n673), .B2(new_n674), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT92), .B1(new_n673), .B2(new_n674), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n499), .ZN(new_n682));
  INV_X1    g0482(.A(new_n500), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(new_n493), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n493), .B(new_n681), .C1(new_n684), .C2(new_n472), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n493), .A2(new_n681), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n494), .A2(new_n498), .A3(new_n501), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n567), .A2(new_n681), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n581), .A2(new_n689), .A3(new_n585), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n567), .A2(new_n580), .A3(new_n681), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(G330), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n581), .A2(new_n585), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n681), .B1(new_n494), .B2(new_n501), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n665), .A2(new_n667), .ZN(new_n697));
  INV_X1    g0497(.A(new_n681), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n695), .A2(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n693), .A2(new_n699), .ZN(G399));
  NOR2_X1   g0500(.A1(new_n207), .A2(G41), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n505), .A2(G116), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n701), .A2(new_n269), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n236), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  INV_X1    g0505(.A(new_n620), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n618), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n656), .A3(new_n659), .A4(new_n606), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT26), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n709), .B(new_n656), .C1(new_n651), .C2(KEYINPUT26), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n621), .A2(new_n585), .A3(new_n629), .A4(new_n659), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n495), .B1(new_n471), .B2(new_n470), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n684), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n711), .B1(new_n713), .B2(new_n581), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT29), .B(new_n698), .C1(new_n710), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n543), .B1(new_n542), .B2(new_n272), .ZN(new_n716));
  AOI211_X1 g0516(.A(KEYINPUT83), .B(G179), .C1(new_n532), .C2(new_n535), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n587), .B1(G190), .B2(new_n542), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n718), .A2(new_n537), .B1(new_n590), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n662), .B1(new_n720), .B2(new_n650), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n656), .B1(new_n708), .B2(KEYINPUT26), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n668), .A2(new_n661), .A3(new_n669), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n681), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n715), .B1(new_n725), .B2(KEYINPUT29), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT93), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n577), .A2(new_n573), .A3(new_n578), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n542), .A2(new_n617), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n729), .B2(new_n471), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT30), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n727), .B(new_n732), .C1(new_n729), .C2(new_n471), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n579), .A2(new_n272), .A3(new_n657), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n497), .A2(new_n624), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n731), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n681), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n494), .A2(new_n498), .A3(new_n501), .ZN(new_n739));
  AND4_X1   g0539(.A1(new_n581), .A2(new_n545), .A3(new_n585), .A4(new_n591), .ZN(new_n740));
  INV_X1    g0540(.A(new_n630), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n739), .A2(new_n740), .A3(new_n741), .A4(new_n698), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n738), .B1(new_n742), .B2(KEYINPUT31), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT94), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n736), .A2(KEYINPUT94), .A3(KEYINPUT31), .A4(new_n681), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(G330), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n726), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n705), .B1(new_n750), .B2(new_n269), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT95), .ZN(G364));
  NOR2_X1   g0552(.A1(new_n206), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n269), .B1(new_n753), .B2(G45), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n207), .B2(G41), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT96), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n232), .B1(G20), .B2(new_n370), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n233), .A2(new_n272), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT98), .Z(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(G190), .A3(new_n327), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n762), .A2(KEYINPUT99), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(KEYINPUT99), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n350), .B1(new_n766), .B2(new_n293), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n233), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n394), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G50), .A2(new_n769), .B1(new_n772), .B2(G107), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n394), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n233), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT100), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G190), .A2(G200), .ZN(new_n777));
  AND3_X1   g0577(.A1(new_n761), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n776), .B1(new_n761), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n773), .B1(new_n217), .B2(new_n775), .C1(new_n780), .C2(new_n341), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n770), .A2(new_n777), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G159), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n767), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n760), .A2(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n786), .B1(new_n284), .B2(new_n789), .C1(new_n215), .C2(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n769), .A2(G326), .ZN(new_n792));
  INV_X1    g0592(.A(G294), .ZN(new_n793));
  INV_X1    g0593(.A(new_n790), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n794), .A2(KEYINPUT101), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(KEYINPUT101), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n353), .B1(new_n793), .B2(new_n775), .C1(new_n797), .C2(new_n461), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n792), .B(new_n798), .C1(new_n788), .C2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n765), .A2(G322), .B1(G329), .B2(new_n783), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n802), .B1(new_n803), .B2(new_n771), .C1(new_n804), .C2(new_n780), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n759), .B1(new_n791), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G13), .A2(G33), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n758), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n207), .A2(new_n350), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(G45), .B2(new_n235), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT97), .ZN(new_n813));
  INV_X1    g0613(.A(new_n255), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n449), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n207), .A2(new_n353), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G355), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(G116), .C2(new_n208), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n757), .B(new_n806), .C1(new_n810), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n809), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n688), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n756), .B1(new_n688), .B2(G330), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(G330), .B2(new_n688), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NOR2_X1   g0625(.A1(new_n368), .A2(new_n698), .ZN(new_n826));
  OAI21_X1  g0626(.A(KEYINPUT103), .B1(new_n373), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n642), .A2(new_n681), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT103), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n644), .A2(new_n828), .A3(new_n829), .A4(new_n367), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n645), .A2(new_n681), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OR3_X1    g0633(.A1(new_n725), .A2(KEYINPUT104), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G330), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n742), .A2(KEYINPUT31), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n737), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n746), .A2(new_n747), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n827), .A2(new_n830), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(new_n698), .C1(new_n670), .C2(new_n664), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT104), .B1(new_n725), .B2(new_n833), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n834), .A2(new_n839), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n757), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT105), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n834), .A2(new_n841), .A3(new_n842), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n749), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n772), .A2(G68), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n765), .A2(G143), .B1(G150), .B2(new_n788), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n769), .A2(G137), .ZN(new_n852));
  INV_X1    g0652(.A(G159), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n780), .ZN(new_n854));
  XOR2_X1   g0654(.A(KEYINPUT102), .B(KEYINPUT34), .Z(new_n855));
  OAI221_X1 g0655(.A(new_n850), .B1(new_n293), .B2(new_n775), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n350), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n859), .B1(new_n211), .B2(new_n797), .C1(new_n860), .C2(new_n782), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n353), .B1(new_n768), .B2(new_n461), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n771), .A2(new_n215), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(G283), .B2(new_n788), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n864), .B1(new_n217), .B2(new_n775), .C1(new_n804), .C2(new_n782), .ZN(new_n865));
  INV_X1    g0665(.A(new_n797), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n862), .B(new_n865), .C1(G107), .C2(new_n866), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n867), .B1(new_n251), .B2(new_n780), .C1(new_n793), .C2(new_n766), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n759), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n758), .A2(new_n807), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n757), .B(new_n869), .C1(new_n362), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n833), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n807), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n849), .A2(new_n874), .ZN(G384));
  AOI21_X1  g0675(.A(new_n251), .B1(new_n600), .B2(KEYINPUT35), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n876), .B(new_n234), .C1(KEYINPUT35), .C2(new_n600), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT36), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n236), .B1(new_n293), .B2(new_n284), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n879), .A2(new_n341), .B1(G50), .B2(new_n284), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(G1), .A3(new_n206), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n308), .A2(new_n300), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n321), .ZN(new_n885));
  INV_X1    g0685(.A(new_n679), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n332), .A2(new_n333), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n639), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n885), .B1(new_n635), .B2(new_n886), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n330), .ZN(new_n892));
  INV_X1    g0692(.A(new_n330), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n679), .B1(new_n310), .B2(new_n321), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n893), .A2(new_n322), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n892), .B1(new_n895), .B2(new_n890), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n883), .B1(new_n889), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n887), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n326), .B2(new_n334), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n634), .A2(new_n886), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n636), .A2(new_n900), .A3(new_n890), .A4(new_n330), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n891), .A2(new_n330), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n901), .B1(new_n902), .B2(new_n890), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n897), .A2(KEYINPUT106), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT106), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n906), .B(new_n883), .C1(new_n889), .C2(new_n896), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n882), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n445), .A2(new_n681), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n636), .A2(new_n900), .A3(new_n330), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n912), .A2(new_n901), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n900), .B1(new_n639), .B2(new_n888), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n883), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT39), .B1(new_n915), .B2(new_n904), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n908), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n644), .A2(new_n681), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n841), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n444), .A2(new_n681), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n447), .B(new_n921), .C1(new_n640), .C2(new_n443), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n435), .A2(new_n444), .A3(new_n681), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n905), .A2(new_n907), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n925), .A2(new_n926), .B1(new_n639), .B2(new_n886), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n917), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT107), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n448), .B(new_n715), .C1(KEYINPUT29), .C2(new_n725), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n649), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT31), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n631), .B2(new_n698), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n744), .B1(new_n934), .B2(new_n738), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n922), .A2(new_n923), .B1(new_n831), .B2(new_n832), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n905), .A2(new_n935), .A3(new_n907), .A4(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  INV_X1    g0738(.A(new_n744), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n743), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n924), .A2(new_n833), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n938), .B1(new_n915), .B2(new_n904), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n937), .A2(new_n938), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT108), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n935), .A2(new_n448), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(G330), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n932), .A2(new_n948), .B1(new_n269), .B2(new_n753), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT109), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n932), .A2(new_n948), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n878), .B(new_n881), .C1(new_n950), .C2(new_n951), .ZN(G367));
  INV_X1    g0752(.A(new_n811), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n810), .B1(new_n208), .B2(new_n513), .C1(new_n246), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n756), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT114), .Z(new_n956));
  NAND2_X1  g0756(.A1(new_n587), .A2(new_n681), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n661), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n656), .B2(new_n957), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n772), .A2(G97), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n789), .B2(new_n793), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT46), .B1(new_n797), .B2(new_n251), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n790), .A2(KEYINPUT46), .A3(new_n251), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n350), .B1(new_n783), .B2(G317), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n804), .B2(new_n768), .ZN(new_n966));
  INV_X1    g0766(.A(new_n775), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n966), .B1(new_n593), .B2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n964), .B(new_n968), .C1(new_n803), .C2(new_n780), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G303), .B2(new_n765), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n350), .B1(new_n341), .B2(new_n771), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT115), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n971), .A2(new_n972), .B1(G137), .B2(new_n783), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n972), .B2(new_n971), .C1(new_n853), .C2(new_n789), .ZN(new_n974));
  INV_X1    g0774(.A(new_n780), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n975), .A2(G50), .B1(G68), .B2(new_n967), .ZN(new_n976));
  INV_X1    g0776(.A(G150), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n976), .B1(new_n766), .B2(new_n977), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n974), .B(new_n978), .C1(G58), .C2(new_n794), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n769), .A2(G143), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT47), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n956), .B1(new_n820), .B2(new_n959), .C1(new_n982), .C2(new_n759), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT112), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n696), .A2(new_n695), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n698), .B1(new_n684), .B2(new_n712), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n986), .A2(new_n690), .A3(new_n691), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n985), .A2(new_n987), .B1(new_n688), .B2(G330), .ZN(new_n988));
  INV_X1    g0788(.A(new_n693), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n726), .A2(new_n749), .A3(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT111), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n726), .A2(new_n749), .A3(new_n990), .A4(KEYINPUT111), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n567), .A2(new_n666), .A3(new_n580), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n666), .B1(new_n567), .B2(new_n580), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n698), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n985), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n606), .A2(new_n681), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n621), .A2(new_n629), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n707), .A2(new_n606), .A3(new_n681), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT44), .B1(new_n699), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT45), .B1(new_n699), .B2(new_n1004), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1004), .B(new_n997), .C1(new_n986), .C2(new_n694), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT45), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1003), .B(new_n1005), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n989), .A2(KEYINPUT110), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n993), .A2(new_n994), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n750), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n701), .B(KEYINPUT41), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n984), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1017), .ZN(new_n1019));
  AOI211_X1 g0819(.A(KEYINPUT112), .B(new_n1019), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n754), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT113), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n985), .A2(new_n1001), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT42), .Z(new_n1025));
  OAI21_X1  g0825(.A(new_n621), .B1(new_n1001), .B2(new_n581), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1026), .A2(new_n698), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1023), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n989), .A2(new_n1004), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1028), .B(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n1021), .A2(new_n1022), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1022), .B1(new_n1021), .B2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n983), .B1(new_n1034), .B2(new_n1035), .ZN(G387));
  AND2_X1   g0836(.A1(new_n336), .A2(new_n339), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n211), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT116), .Z(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT50), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n284), .A2(new_n362), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1040), .A2(G45), .A3(new_n1041), .A4(new_n702), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n953), .B1(new_n242), .B2(G45), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n702), .B2(new_n816), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1042), .A2(new_n1044), .B1(G107), .B2(new_n208), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n757), .B1(new_n1045), .B2(new_n810), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n692), .B2(new_n820), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n782), .A2(new_n977), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n967), .A2(new_n344), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n341), .A2(new_n790), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n975), .B2(G68), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1049), .B(new_n1051), .C1(new_n766), .C2(new_n211), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1048), .B(new_n1052), .C1(G159), .C2(new_n769), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n788), .A2(new_n316), .A3(new_n313), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1053), .A2(new_n350), .A3(new_n960), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n765), .A2(G317), .B1(G311), .B2(new_n788), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n769), .A2(G322), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n461), .C2(new_n780), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT48), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n803), .B2(new_n775), .C1(new_n793), .C2(new_n790), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n772), .A2(G116), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n783), .A2(G326), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1062), .A2(new_n353), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1055), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1047), .B1(new_n1067), .B2(new_n758), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n754), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n990), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n993), .A2(new_n994), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n701), .C1(new_n1015), .C2(new_n990), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(G393));
  XNOR2_X1  g0873(.A(new_n1010), .B(new_n989), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1075), .A2(new_n701), .A3(new_n1014), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n765), .A2(G311), .B1(G317), .B2(new_n769), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT52), .Z(new_n1078));
  NAND2_X1  g0878(.A1(new_n975), .A2(G294), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n783), .A2(G322), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1078), .A2(new_n353), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n789), .A2(new_n461), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n790), .A2(new_n803), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n775), .A2(new_n251), .B1(new_n771), .B2(new_n249), .ZN(new_n1084));
  NOR4_X1   g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n353), .B1(new_n975), .B2(new_n1037), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n775), .A2(new_n362), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n863), .B(new_n1087), .C1(G50), .C2(new_n788), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(new_n284), .C2(new_n790), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n765), .A2(G159), .B1(G150), .B2(new_n769), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n1091));
  XNOR2_X1  g0891(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1089), .B(new_n1092), .C1(G143), .C2(new_n783), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n758), .B1(new_n1085), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n252), .A2(new_n811), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n810), .C1(new_n217), .C2(new_n208), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n756), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1004), .A2(new_n820), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT117), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1097), .A2(new_n1099), .B1(new_n1074), .B2(new_n754), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1076), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  OAI21_X1  g0902(.A(new_n353), .B1(new_n768), .B2(new_n803), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1087), .B1(new_n593), .B2(new_n788), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1104), .B(new_n850), .C1(new_n793), .C2(new_n782), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(G87), .C2(new_n866), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n217), .B2(new_n780), .C1(new_n251), .C2(new_n766), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n353), .B1(new_n772), .B2(G50), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT119), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n765), .A2(G132), .B1(G128), .B2(new_n769), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT120), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(G125), .C2(new_n783), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n788), .A2(G137), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n967), .A2(G159), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT54), .B(G143), .Z(new_n1116));
  AOI22_X1  g0916(.A1(new_n975), .A2(new_n1116), .B1(new_n1109), .B2(new_n1108), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n794), .A2(G150), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT53), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1107), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n757), .B1(new_n1121), .B2(new_n758), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n317), .A2(new_n870), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n916), .B1(new_n926), .B2(KEYINPUT39), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(new_n1123), .C1(new_n808), .C2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n909), .B1(new_n915), .B2(new_n904), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n710), .A2(new_n714), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1127), .A2(new_n681), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n918), .B1(new_n1128), .B2(new_n840), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n924), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n909), .B1(new_n920), .B2(new_n924), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n1124), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n935), .A2(G330), .A3(new_n936), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n839), .A2(new_n833), .A3(new_n924), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1131), .B(new_n1137), .C1(new_n1124), .C2(new_n1132), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1125), .B1(new_n1139), .B2(new_n754), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n935), .A2(new_n448), .A3(G330), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n649), .A2(new_n930), .A3(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(G330), .B(new_n833), .C1(new_n743), .C2(new_n748), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1130), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1134), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n920), .ZN(new_n1146));
  OAI211_X1 g0946(.A(G330), .B(new_n833), .C1(new_n743), .C2(new_n939), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1130), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1137), .A2(new_n1129), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1142), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1136), .A2(new_n1150), .A3(new_n1138), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1151), .A2(new_n701), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1150), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1139), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1140), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(G378));
  NAND2_X1  g0956(.A1(new_n937), .A2(new_n938), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n942), .A2(new_n943), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(G330), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1124), .A2(new_n909), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n926), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1130), .B1(new_n841), .B2(new_n919), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1161), .A2(new_n1162), .B1(new_n326), .B2(new_n679), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1159), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(G330), .B(new_n944), .C1(new_n917), .C2(new_n927), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n409), .B(KEYINPUT55), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n679), .B1(new_n380), .B2(new_n381), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1169), .B(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1166), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1164), .A2(new_n1165), .A3(new_n1172), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n1069), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n211), .B1(new_n264), .B2(G41), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n975), .A2(G137), .B1(G125), .B2(new_n769), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n967), .A2(G150), .B1(new_n794), .B2(new_n1116), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(G128), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n766), .C1(new_n860), .C2(new_n789), .ZN(new_n1182));
  AOI21_X1  g0982(.A(G33), .B1(new_n1182), .B2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n772), .A2(G159), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT121), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(G124), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(G124), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n783), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1183), .A2(new_n258), .A3(new_n1184), .A4(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1177), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n788), .A2(G97), .B1(G283), .B2(new_n783), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n251), .B2(new_n768), .ZN(new_n1193));
  OR4_X1    g0993(.A1(G41), .A2(new_n1193), .A3(new_n350), .A4(new_n1050), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n344), .B2(new_n975), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n967), .A2(G68), .B1(new_n772), .B2(G58), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n249), .C2(new_n766), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT58), .Z(new_n1198));
  OAI21_X1  g0998(.A(new_n758), .B1(new_n1191), .B2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT122), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n757), .B1(new_n211), .B2(new_n870), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n1172), .C2(new_n808), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1176), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1142), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1151), .A2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1205), .A2(new_n1174), .A3(KEYINPUT57), .A4(new_n1175), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n701), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1164), .A2(new_n1165), .A3(new_n1172), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1172), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT57), .B1(new_n1210), .B2(new_n1205), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1203), .B1(new_n1207), .B2(new_n1211), .ZN(G375));
  NOR2_X1   g1012(.A1(new_n782), .A2(new_n1181), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n765), .A2(G137), .B1(G159), .B2(new_n866), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n788), .A2(new_n1116), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n293), .B2(new_n771), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n353), .B(new_n1216), .C1(G132), .C2(new_n769), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1214), .B(new_n1217), .C1(new_n977), .C2(new_n780), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1213), .B(new_n1218), .C1(G50), .C2(new_n967), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1049), .B1(new_n780), .B2(new_n354), .C1(new_n766), .C2(new_n803), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n789), .A2(new_n251), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n797), .A2(new_n217), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n353), .B1(new_n771), .B2(new_n362), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT124), .Z(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n793), .B2(new_n768), .C1(new_n461), .C2(new_n782), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n758), .B1(new_n1219), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n870), .A2(new_n284), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n756), .A3(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n924), .A2(new_n808), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1232), .B2(new_n1069), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1232), .A2(new_n1204), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(new_n1019), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1234), .B1(new_n1236), .B2(new_n1153), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(G381));
  NAND2_X1  g1038(.A1(new_n1176), .A2(new_n1202), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1206), .A2(new_n701), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1210), .A2(new_n1205), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT57), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1239), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1155), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1070), .A2(new_n824), .A3(new_n1072), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n983), .B(new_n1101), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1248), .A2(G384), .A3(G381), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(G407));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT63), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n680), .A2(G213), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1203), .B(new_n1155), .C1(new_n1019), .C2(new_n1241), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(new_n1244), .C2(new_n1155), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1146), .A2(new_n1149), .A3(KEYINPUT60), .A4(new_n1142), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1257), .B(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1232), .B2(new_n1204), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n701), .A3(new_n1153), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1233), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(G384), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G384), .B(new_n1233), .C1(new_n1259), .C2(new_n1262), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n680), .A2(G213), .A3(G2897), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1268), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1253), .B1(new_n1256), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G375), .A2(G378), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1267), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1252), .B1(new_n1273), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1246), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1248), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT112), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1016), .A2(new_n984), .A3(new_n1017), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1069), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(KEYINPUT113), .B1(new_n1287), .B2(new_n1032), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1021), .A2(new_n1022), .A3(new_n1033), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1101), .B1(new_n1290), .B2(new_n983), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1281), .B1(new_n1283), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G387), .A2(G390), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1293), .A2(new_n1282), .A3(new_n1248), .A4(new_n1280), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1292), .B(new_n1294), .C1(new_n1253), .C2(new_n1276), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1278), .A2(new_n1295), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(G375), .A2(G378), .B1(G213), .B2(new_n680), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT62), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1275), .A4(new_n1255), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1300), .A2(new_n1252), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n1276), .A2(KEYINPUT62), .B1(new_n1256), .B2(new_n1272), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1297), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT127), .B1(new_n1296), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1276), .A2(KEYINPUT62), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1256), .A2(new_n1272), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1305), .A2(new_n1306), .A3(new_n1252), .A4(new_n1300), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1309), .B(new_n1310), .C1(new_n1295), .C2(new_n1278), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1304), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(new_n1245), .A2(new_n1274), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1292), .A2(new_n1313), .A3(new_n1294), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1316), .B(new_n1267), .ZN(G402));
endmodule


