//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  OR2_X1    g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n453), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G2105), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT68), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G137), .A4(new_n468), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n470), .A2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n473), .A2(KEYINPUT69), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n473), .A2(KEYINPUT69), .ZN(new_n482));
  OAI21_X1  g057(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n480), .B1(new_n484), .B2(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n468), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NOR2_X1   g065(.A1(new_n468), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT70), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n494), .A2(new_n496), .A3(new_n497), .A4(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n463), .B2(new_n464), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n503), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n473), .A2(new_n505), .A3(new_n501), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n473), .A2(G126), .A3(G2105), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n499), .A2(new_n504), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(new_n521), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n520), .A2(new_n526), .ZN(G166));
  INV_X1    g102(.A(new_n524), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XOR2_X1   g108(.A(KEYINPUT73), .B(G51), .Z(new_n534));
  NAND2_X1  g109(.A1(new_n522), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n529), .A2(new_n530), .A3(new_n533), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n522), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n524), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT75), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n519), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AOI22_X1  g120(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n519), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n517), .A2(G81), .A3(new_n521), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n522), .A2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n522), .A2(new_n560), .A3(G53), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n521), .A2(G53), .A3(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT77), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n528), .A2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n515), .A2(new_n516), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n561), .A2(new_n572), .A3(new_n563), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n565), .A2(new_n566), .A3(new_n571), .A4(new_n573), .ZN(G299));
  OR2_X1    g149(.A1(new_n520), .A2(new_n526), .ZN(G303));
  NAND2_X1  g150(.A1(new_n528), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n522), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n515), .A2(G61), .A3(new_n516), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n515), .A2(G86), .A3(new_n516), .A4(new_n521), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n568), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(KEYINPUT78), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(KEYINPUT78), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n528), .A2(G85), .B1(G47), .B2(new_n522), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G290));
  NAND3_X1  g173(.A1(new_n528), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n524), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT81), .Z(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n568), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G54), .B2(new_n522), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT80), .B1(new_n610), .B2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  MUX2_X1   g187(.A(KEYINPUT80), .B(new_n611), .S(new_n612), .Z(G284));
  MUX2_X1   g188(.A(KEYINPUT80), .B(new_n611), .S(new_n612), .Z(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n610), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n610), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n554), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT82), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n473), .A2(new_n469), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n631));
  INV_X1    g206(.A(G135), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n631), .B1(new_n486), .B2(new_n632), .C1(new_n633), .C2(new_n483), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n635), .A3(new_n636), .ZN(G156));
  XOR2_X1   g212(.A(KEYINPUT15), .B(G2435), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT85), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT84), .B(KEYINPUT14), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n641), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n649), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT86), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n669), .A2(new_n670), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n673), .A3(new_n671), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n678), .C1(new_n673), .C2(new_n677), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G32), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n484), .A2(G129), .ZN(new_n688));
  NAND3_X1  g263(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT26), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  AOI22_X1  g267(.A1(new_n691), .A2(new_n692), .B1(G105), .B2(new_n469), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n487), .A2(G141), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n687), .B1(new_n697), .B2(new_n686), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT27), .ZN(new_n699));
  INV_X1    g274(.A(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G20), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT23), .Z(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G299), .B2(G16), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT102), .B(G1956), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n686), .A2(G26), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  OAI21_X1  g284(.A(KEYINPUT96), .B1(G104), .B2(G2105), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g286(.A1(KEYINPUT96), .A2(G104), .A3(G2105), .ZN(new_n712));
  OAI221_X1 g287(.A(G2104), .B1(G116), .B2(new_n468), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G140), .ZN(new_n714));
  INV_X1    g289(.A(G128), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n713), .B1(new_n486), .B2(new_n714), .C1(new_n715), .C2(new_n483), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n709), .B1(new_n716), .B2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G2067), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n705), .A2(new_n706), .ZN(new_n720));
  NOR4_X1   g295(.A1(new_n701), .A2(new_n707), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n702), .A2(G5), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G171), .B2(new_n702), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT101), .B(G1961), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n686), .A2(G35), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n686), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n554), .A2(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G16), .B2(G19), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT95), .B(G1341), .Z(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI22_X1  g307(.A1(new_n728), .A2(G2090), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G2090), .B2(new_n728), .ZN(new_n734));
  INV_X1    g309(.A(G21), .ZN(new_n735));
  AOI21_X1  g310(.A(KEYINPUT99), .B1(new_n702), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G286), .A2(new_n702), .ZN(new_n737));
  MUX2_X1   g312(.A(new_n736), .B(KEYINPUT99), .S(new_n737), .Z(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT100), .B(G1966), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n738), .B(new_n739), .Z(new_n740));
  AND2_X1   g315(.A1(new_n487), .A2(G139), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  AOI22_X1  g318(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n468), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(new_n686), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n686), .B2(G33), .ZN(new_n748));
  INV_X1    g323(.A(G2072), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT98), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n730), .A2(new_n732), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n686), .A2(G27), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G164), .B2(new_n686), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n748), .A2(new_n749), .B1(G2078), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G160), .A2(new_n686), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n757));
  INV_X1    g332(.A(G34), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n686), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2084), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT31), .B(G11), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n764), .A2(G28), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n686), .B1(new_n764), .B2(G28), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n763), .B1(new_n765), .B2(new_n766), .C1(new_n634), .C2(new_n686), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n754), .A2(G2078), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n752), .A2(new_n755), .A3(new_n762), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G4), .A2(G16), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n610), .B2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1348), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n740), .A2(new_n751), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n721), .A2(new_n725), .A3(new_n734), .A4(new_n774), .ZN(new_n775));
  MUX2_X1   g350(.A(G23), .B(G288), .S(G16), .Z(new_n776));
  XOR2_X1   g351(.A(KEYINPUT33), .B(G1976), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n702), .A2(G22), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT91), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G166), .B2(new_n702), .ZN(new_n781));
  INV_X1    g356(.A(G1971), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n778), .B1(KEYINPUT92), .B2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT34), .ZN(new_n785));
  NOR2_X1   g360(.A1(G6), .A2(G16), .ZN(new_n786));
  INV_X1    g361(.A(G305), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT90), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT32), .B(G1981), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n783), .A2(KEYINPUT92), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n784), .A2(new_n785), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n702), .A2(G24), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT89), .Z(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G290), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1986), .ZN(new_n797));
  NAND2_X1  g372(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n686), .A2(G25), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n487), .A2(G131), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n484), .A2(G119), .ZN(new_n801));
  OR2_X1    g376(.A1(G95), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT88), .Z(new_n804));
  NAND3_X1  g379(.A1(new_n800), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n799), .B1(new_n806), .B2(new_n686), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  AND4_X1   g384(.A1(new_n793), .A2(new_n797), .A3(new_n798), .A4(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n784), .A2(new_n791), .A3(new_n792), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n811), .A2(new_n812), .A3(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT93), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n810), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n816), .A2(new_n818), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n775), .B1(new_n819), .B2(new_n820), .ZN(G311));
  INV_X1    g396(.A(new_n775), .ZN(new_n822));
  INV_X1    g397(.A(new_n820), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n816), .A2(new_n818), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(G150));
  NAND2_X1  g400(.A1(new_n610), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n519), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n522), .A2(G55), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n524), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n553), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n833), .B(new_n547), .C1(new_n551), .C2(new_n552), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n827), .B(new_n837), .Z(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n833), .A2(new_n840), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(G145));
  INV_X1    g420(.A(KEYINPUT104), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n805), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n627), .ZN(new_n848));
  OR2_X1    g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n849), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n850));
  INV_X1    g425(.A(G142), .ZN(new_n851));
  INV_X1    g426(.A(G130), .ZN(new_n852));
  OAI221_X1 g427(.A(new_n850), .B1(new_n486), .B2(new_n851), .C1(new_n852), .C2(new_n483), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n848), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n696), .A2(new_n716), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n696), .A2(new_n716), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(G164), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(G164), .B1(new_n858), .B2(new_n859), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n857), .B(new_n746), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n746), .A2(new_n857), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT103), .B1(new_n741), .B2(new_n745), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n860), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n856), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n854), .A2(new_n863), .A3(new_n867), .A4(new_n855), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n489), .B(new_n634), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G160), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  INV_X1    g450(.A(new_n873), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(new_n876), .A3(new_n870), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g454(.A(G868), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n834), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G303), .B(G288), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n596), .A2(G305), .A3(new_n597), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(G305), .B1(new_n596), .B2(new_n597), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n882), .A3(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(KEYINPUT42), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT42), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n892), .A2(KEYINPUT106), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT106), .B1(new_n892), .B2(new_n893), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n610), .A2(new_n616), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n609), .A2(G299), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT41), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(KEYINPUT105), .A3(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n837), .B(new_n621), .Z(new_n905));
  AND2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n898), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n895), .A2(new_n909), .ZN(new_n910));
  OAI221_X1 g485(.A(KEYINPUT106), .B1(new_n906), .B2(new_n908), .C1(new_n892), .C2(new_n893), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n894), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n881), .B1(new_n912), .B2(new_n880), .ZN(G295));
  OAI21_X1  g488(.A(new_n881), .B1(new_n912), .B2(new_n880), .ZN(G331));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n915));
  AOI21_X1  g490(.A(G301), .B1(new_n835), .B2(new_n836), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n835), .A2(G301), .A3(new_n836), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(G168), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(G286), .B1(new_n920), .B2(new_n916), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n907), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n902), .A2(new_n919), .A3(new_n921), .A4(new_n903), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G37), .B1(new_n925), .B2(new_n891), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n890), .A3(new_n924), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n915), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n899), .A2(new_n901), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n919), .A2(new_n921), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n898), .B1(new_n919), .B2(new_n921), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n891), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND4_X1   g507(.A1(new_n915), .A2(new_n932), .A3(new_n927), .A4(new_n875), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n928), .A2(new_n933), .A3(KEYINPUT44), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n915), .A3(new_n927), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n927), .A3(new_n875), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n935), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n934), .A2(new_n939), .ZN(G397));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT45), .B1(new_n508), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n470), .A2(G40), .A3(new_n476), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NOR3_X1   g521(.A1(G290), .A2(G1986), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n945), .A2(G1986), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(G290), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT107), .Z(new_n950));
  XNOR2_X1  g525(.A(new_n716), .B(new_n718), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(new_n946), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT108), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n696), .B(G1996), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n945), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n806), .A2(new_n808), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n806), .A2(new_n808), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n945), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n950), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1976), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT52), .B1(G288), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n508), .A2(new_n941), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n470), .A2(G40), .A3(new_n476), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n508), .A2(KEYINPUT109), .A3(new_n941), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n576), .A2(G1976), .A3(new_n577), .A4(new_n578), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n962), .A2(G8), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(G8), .A3(new_n969), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT52), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1981), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n583), .A2(new_n586), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n519), .B1(new_n580), .B2(new_n581), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n584), .A2(new_n585), .ZN(new_n978));
  OAI21_X1  g553(.A(G1981), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n975), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n981));
  NAND3_X1  g556(.A1(G305), .A2(KEYINPUT111), .A3(G1981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n981), .B1(new_n980), .B2(new_n982), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n968), .A2(G8), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n973), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  NAND3_X1  g563(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(G166), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT110), .B1(new_n963), .B2(KEYINPUT50), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n995), .B(new_n996), .C1(new_n508), .C2(new_n941), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G2090), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n965), .A2(new_n996), .A3(new_n967), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n966), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n963), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n966), .A3(new_n943), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n782), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n991), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n987), .B(new_n988), .C1(new_n993), .C2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1001), .B(new_n966), .C1(new_n994), .C2(new_n997), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1006), .B1(new_n1009), .B2(G2090), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n993), .B1(new_n1010), .B2(G8), .ZN(new_n1011));
  INV_X1    g586(.A(new_n985), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n972), .B(new_n970), .C1(new_n1014), .C2(new_n984), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT114), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G168), .A2(G8), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n508), .A2(KEYINPUT109), .A3(new_n941), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT109), .B1(new_n508), .B2(new_n941), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n966), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1004), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1021), .B2(new_n966), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n739), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1009), .A2(G2084), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1017), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT63), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n1007), .B2(new_n993), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1008), .A2(new_n1016), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1030), .A2(new_n1028), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(KEYINPUT115), .A3(new_n1008), .A4(new_n1016), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT113), .B(KEYINPUT63), .Z(new_n1036));
  NAND2_X1  g611(.A1(new_n1007), .A2(new_n993), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n508), .A2(new_n996), .A3(new_n941), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n966), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n965), .A2(new_n967), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(KEYINPUT50), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1041), .A2(new_n1000), .B1(new_n1005), .B2(new_n782), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n992), .B(new_n989), .C1(new_n1042), .C2(new_n991), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(new_n1043), .A3(new_n987), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1028), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1036), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1033), .A2(new_n1035), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1037), .ZN(new_n1048));
  OR2_X1    g623(.A1(G288), .A2(G1976), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n975), .B1(new_n986), .B2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1048), .A2(new_n987), .B1(new_n1012), .B2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n528), .A2(G91), .B1(new_n570), .B2(G651), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT57), .B1(new_n561), .B2(new_n563), .ZN(new_n1053));
  AOI22_X1  g628(.A1(G299), .A2(KEYINPUT57), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(new_n749), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1004), .A2(new_n966), .A3(new_n943), .A4(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1054), .B(new_n1057), .C1(new_n1041), .C2(G1956), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n968), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT117), .A4(new_n967), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n718), .ZN(new_n1064));
  INV_X1    g639(.A(G1348), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1009), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n610), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n616), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1057), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT50), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n944), .B1(new_n1003), .B2(new_n996), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1956), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1071), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1059), .B1(new_n1068), .B2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT58), .B(G1341), .Z(new_n1079));
  NAND3_X1  g654(.A1(new_n1061), .A2(new_n1062), .A3(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1004), .A2(new_n700), .A3(new_n966), .A4(new_n943), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT118), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(KEYINPUT118), .A3(new_n1081), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1078), .B1(new_n1085), .B2(new_n554), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT61), .B1(new_n1058), .B2(KEYINPUT120), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1076), .A2(new_n1058), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1076), .B(new_n1058), .C1(KEYINPUT120), .C2(KEYINPUT61), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1080), .A2(KEYINPUT118), .A3(new_n1081), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n554), .B(new_n1078), .C1(new_n1092), .C2(new_n1082), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1086), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1064), .A2(KEYINPUT60), .A3(new_n1066), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n609), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n609), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT60), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1067), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1077), .B1(new_n1095), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1025), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(G2078), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1106), .A2(new_n1004), .A3(new_n1023), .A4(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1005), .B2(G2078), .ZN(new_n1110));
  INV_X1    g685(.A(G1961), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1001), .A2(new_n966), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n998), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1109), .A2(G301), .A3(new_n1110), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1118));
  OR2_X1    g693(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1119));
  NAND2_X1  g694(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1107), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n943), .B2(new_n966), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n942), .A2(new_n944), .A3(KEYINPUT122), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1004), .B(new_n1121), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1113), .A2(new_n1110), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1113), .A2(new_n1110), .A3(new_n1125), .A4(KEYINPUT125), .ZN(new_n1129));
  AND4_X1   g704(.A1(KEYINPUT126), .A2(new_n1128), .A3(G171), .A4(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(G301), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT126), .B1(new_n1131), .B2(new_n1129), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1116), .B(new_n1118), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1026), .A2(G168), .A3(new_n1027), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(G8), .ZN(new_n1135));
  AOI21_X1  g710(.A(G168), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT51), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1134), .A2(new_n1138), .A3(G8), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NOR4_X1   g715(.A1(new_n1024), .A2(new_n1025), .A3(new_n1107), .A4(G2078), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1113), .A2(new_n1110), .ZN(new_n1142));
  OAI21_X1  g717(.A(G171), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1126), .A2(G171), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1044), .B1(new_n1145), .B2(new_n1117), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1133), .A2(new_n1140), .A3(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1047), .B(new_n1051), .C1(new_n1105), .C2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1140), .A2(KEYINPUT62), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1044), .A2(new_n1143), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n960), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT46), .B1(new_n945), .B2(new_n700), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT127), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n696), .B1(KEYINPUT46), .B2(new_n700), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1157), .A2(new_n951), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1158), .B2(new_n946), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT47), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n947), .B(KEYINPUT48), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n959), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n955), .A2(new_n956), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n716), .A2(G2067), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n946), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1154), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g742(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1169));
  NOR2_X1   g743(.A1(G229), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g744(.A(new_n878), .B(new_n1170), .C1(new_n928), .C2(new_n933), .ZN(G225));
  INV_X1    g745(.A(G225), .ZN(G308));
endmodule


