

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771;

  XNOR2_X1 U383 ( .A(n757), .B(n468), .ZN(n548) );
  XNOR2_X1 U384 ( .A(n532), .B(n360), .ZN(n757) );
  XNOR2_X1 U385 ( .A(n391), .B(n466), .ZN(n360) );
  XNOR2_X1 U386 ( .A(n392), .B(G131), .ZN(n521) );
  INV_X1 U387 ( .A(KEYINPUT66), .ZN(n392) );
  NOR2_X2 U388 ( .A1(n692), .A2(n421), .ZN(n693) );
  NOR2_X1 U389 ( .A1(n676), .A2(n700), .ZN(n562) );
  INV_X1 U390 ( .A(G953), .ZN(n760) );
  XNOR2_X2 U391 ( .A(n641), .B(n640), .ZN(n381) );
  XNOR2_X2 U392 ( .A(n477), .B(KEYINPUT15), .ZN(n642) );
  NAND2_X2 U393 ( .A1(n397), .A2(n393), .ZN(n769) );
  AND2_X2 U394 ( .A1(n380), .A2(n400), .ZN(n397) );
  NOR2_X1 U395 ( .A1(n558), .A2(n631), .ZN(n559) );
  AND2_X2 U396 ( .A1(n405), .A2(n404), .ZN(n742) );
  NAND2_X1 U397 ( .A1(n435), .A2(n376), .ZN(n405) );
  AND2_X1 U398 ( .A1(n583), .A2(n433), .ZN(n432) );
  XNOR2_X1 U399 ( .A(n409), .B(n408), .ZN(n770) );
  NAND2_X1 U400 ( .A1(n449), .A2(n417), .ZN(n409) );
  NOR2_X1 U401 ( .A1(n590), .A2(n594), .ZN(n555) );
  XNOR2_X1 U402 ( .A(n578), .B(KEYINPUT109), .ZN(n678) );
  XNOR2_X1 U403 ( .A(KEYINPUT6), .B(n631), .ZN(n619) );
  XNOR2_X1 U404 ( .A(n539), .B(n414), .ZN(n578) );
  XNOR2_X1 U405 ( .A(n472), .B(n471), .ZN(n482) );
  XNOR2_X1 U406 ( .A(n379), .B(KEYINPUT79), .ZN(n487) );
  XNOR2_X1 U407 ( .A(G143), .B(G128), .ZN(n379) );
  INV_X1 U408 ( .A(n561), .ZN(n361) );
  XOR2_X1 U409 ( .A(G122), .B(G116), .Z(n533) );
  NOR2_X1 U410 ( .A1(n628), .A2(n627), .ZN(n455) );
  XNOR2_X1 U411 ( .A(n468), .B(G125), .ZN(n500) );
  XNOR2_X1 U412 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n621) );
  XNOR2_X1 U413 ( .A(n482), .B(n388), .ZN(n387) );
  XNOR2_X1 U414 ( .A(n533), .B(n389), .ZN(n388) );
  INV_X1 U415 ( .A(KEYINPUT16), .ZN(n389) );
  AND2_X1 U416 ( .A1(n450), .A2(n452), .ZN(n449) );
  NAND2_X1 U417 ( .A1(n455), .A2(n454), .ZN(n453) );
  AND2_X1 U418 ( .A1(n382), .A2(n383), .ZN(n582) );
  XOR2_X1 U419 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n517) );
  XNOR2_X1 U420 ( .A(n378), .B(n503), .ZN(n708) );
  XNOR2_X1 U421 ( .A(n507), .B(KEYINPUT25), .ZN(n378) );
  XNOR2_X1 U422 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U423 ( .A(G101), .B(G113), .ZN(n480) );
  XNOR2_X1 U424 ( .A(n521), .B(KEYINPUT67), .ZN(n391) );
  NAND2_X1 U425 ( .A1(n464), .A2(n600), .ZN(n641) );
  XNOR2_X1 U426 ( .A(n565), .B(KEYINPUT1), .ZN(n441) );
  XNOR2_X1 U427 ( .A(KEYINPUT8), .B(KEYINPUT65), .ZN(n496) );
  XNOR2_X1 U428 ( .A(n535), .B(n533), .ZN(n419) );
  XNOR2_X1 U429 ( .A(n524), .B(n523), .ZN(n655) );
  XNOR2_X1 U430 ( .A(n462), .B(n522), .ZN(n523) );
  XNOR2_X1 U431 ( .A(n758), .B(n415), .ZN(n524) );
  XNOR2_X1 U432 ( .A(n490), .B(n752), .ZN(n647) );
  XNOR2_X1 U433 ( .A(n364), .B(KEYINPUT41), .ZN(n728) );
  NOR2_X1 U434 ( .A1(n697), .A2(n386), .ZN(n385) );
  INV_X1 U435 ( .A(n694), .ZN(n386) );
  XNOR2_X1 U436 ( .A(n577), .B(n576), .ZN(n598) );
  NAND2_X1 U437 ( .A1(n428), .A2(n366), .ZN(n577) );
  OR2_X1 U438 ( .A1(n633), .A2(n373), .ZN(n447) );
  INV_X1 U439 ( .A(n445), .ZN(n399) );
  AND2_X1 U440 ( .A1(n444), .A2(n395), .ZN(n394) );
  NOR2_X1 U441 ( .A1(n445), .A2(n410), .ZN(n395) );
  NOR2_X1 U442 ( .A1(n619), .A2(KEYINPUT78), .ZN(n451) );
  NOR2_X1 U443 ( .A1(n561), .A2(n560), .ZN(n580) );
  INV_X1 U444 ( .A(KEYINPUT28), .ZN(n420) );
  INV_X1 U445 ( .A(KEYINPUT104), .ZN(n414) );
  XNOR2_X1 U446 ( .A(n413), .B(n374), .ZN(n624) );
  NOR2_X1 U447 ( .A1(n617), .A2(n424), .ZN(n413) );
  BUF_X1 U448 ( .A(n441), .Z(n439) );
  NAND2_X1 U449 ( .A1(n742), .A2(G472), .ZN(n403) );
  NAND2_X1 U450 ( .A1(G953), .A2(G902), .ZN(n607) );
  INV_X1 U451 ( .A(KEYINPUT44), .ZN(n422) );
  XNOR2_X1 U452 ( .A(n637), .B(n423), .ZN(n456) );
  INV_X1 U453 ( .A(KEYINPUT106), .ZN(n423) );
  XNOR2_X1 U454 ( .A(n518), .B(n370), .ZN(n415) );
  XNOR2_X1 U455 ( .A(G104), .B(KEYINPUT12), .ZN(n516) );
  XNOR2_X1 U456 ( .A(G143), .B(G122), .ZN(n519) );
  XOR2_X1 U457 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n520) );
  XNOR2_X1 U458 ( .A(KEYINPUT4), .B(KEYINPUT76), .ZN(n483) );
  XOR2_X1 U459 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n484) );
  XNOR2_X1 U460 ( .A(G902), .B(KEYINPUT90), .ZN(n477) );
  OR2_X1 U461 ( .A1(G902), .A2(G237), .ZN(n553) );
  NOR2_X1 U462 ( .A1(n627), .A2(n709), .ZN(n515) );
  NAND2_X1 U463 ( .A1(n446), .A2(n616), .ZN(n445) );
  NAND2_X1 U464 ( .A1(n633), .A2(n373), .ZN(n446) );
  INV_X1 U465 ( .A(KEYINPUT35), .ZN(n410) );
  INV_X1 U466 ( .A(n619), .ZN(n454) );
  INV_X1 U467 ( .A(KEYINPUT74), .ZN(n411) );
  NOR2_X1 U468 ( .A1(n709), .A2(n708), .ZN(n706) );
  XNOR2_X1 U469 ( .A(n406), .B(n375), .ZN(n617) );
  NAND2_X1 U470 ( .A1(n612), .A2(n425), .ZN(n424) );
  INV_X1 U471 ( .A(n709), .ZN(n425) );
  XNOR2_X1 U472 ( .A(n481), .B(n416), .ZN(n543) );
  XNOR2_X1 U473 ( .A(n478), .B(KEYINPUT70), .ZN(n416) );
  XNOR2_X1 U474 ( .A(G119), .B(KEYINPUT91), .ZN(n478) );
  XNOR2_X1 U475 ( .A(G116), .B(KEYINPUT97), .ZN(n540) );
  XOR2_X1 U476 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n541) );
  NOR2_X1 U477 ( .A1(G953), .A2(G237), .ZN(n544) );
  XNOR2_X1 U478 ( .A(G110), .B(G119), .ZN(n492) );
  XNOR2_X1 U479 ( .A(G128), .B(G137), .ZN(n491) );
  XNOR2_X1 U480 ( .A(n500), .B(G140), .ZN(n501) );
  XNOR2_X1 U481 ( .A(n548), .B(n474), .ZN(n732) );
  XOR2_X1 U482 ( .A(G140), .B(G101), .Z(n470) );
  NAND2_X1 U483 ( .A1(G234), .A2(G237), .ZN(n511) );
  INV_X1 U484 ( .A(n641), .ZN(n402) );
  NOR2_X1 U485 ( .A1(n630), .A2(n430), .ZN(n428) );
  INV_X1 U486 ( .A(n573), .ZN(n430) );
  INV_X1 U487 ( .A(n439), .ZN(n628) );
  BUF_X1 U488 ( .A(n617), .Z(n633) );
  XNOR2_X1 U489 ( .A(n534), .B(n419), .ZN(n536) );
  XOR2_X1 U490 ( .A(G107), .B(KEYINPUT103), .Z(n531) );
  XNOR2_X1 U491 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X1 U492 ( .A1(n760), .A2(G952), .ZN(n746) );
  XNOR2_X1 U493 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U494 ( .A(n581), .B(n384), .ZN(n383) );
  INV_X1 U495 ( .A(KEYINPUT42), .ZN(n384) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n771) );
  XNOR2_X1 U497 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n437) );
  NAND2_X1 U498 ( .A1(n396), .A2(n394), .ZN(n393) );
  INV_X1 U499 ( .A(KEYINPUT32), .ZN(n408) );
  NOR2_X1 U500 ( .A1(n624), .A2(n619), .ZN(n629) );
  XNOR2_X1 U501 ( .A(n403), .B(n644), .ZN(n645) );
  XOR2_X1 U502 ( .A(KEYINPUT62), .B(n643), .Z(n644) );
  AND2_X1 U503 ( .A1(n611), .A2(n610), .ZN(n362) );
  AND2_X1 U504 ( .A1(n749), .A2(KEYINPUT2), .ZN(n363) );
  AND2_X1 U505 ( .A1(n695), .A2(n385), .ZN(n364) );
  AND2_X1 U506 ( .A1(G210), .A2(n553), .ZN(n365) );
  XNOR2_X1 U507 ( .A(n457), .B(KEYINPUT19), .ZN(n601) );
  AND2_X1 U508 ( .A1(n429), .A2(n695), .ZN(n366) );
  NOR2_X1 U509 ( .A1(n664), .A2(n456), .ZN(n367) );
  AND2_X1 U510 ( .A1(n749), .A2(n436), .ZN(n368) );
  OR2_X1 U511 ( .A1(n592), .A2(n591), .ZN(n369) );
  AND2_X1 U512 ( .A1(n544), .A2(G214), .ZN(n370) );
  NOR2_X1 U513 ( .A1(n730), .A2(n465), .ZN(n371) );
  INV_X1 U514 ( .A(G146), .ZN(n468) );
  AND2_X1 U515 ( .A1(n455), .A2(n451), .ZN(n372) );
  NAND2_X1 U516 ( .A1(n363), .A2(n402), .ZN(n404) );
  XOR2_X1 U517 ( .A(n623), .B(KEYINPUT72), .Z(n373) );
  XOR2_X1 U518 ( .A(n613), .B(KEYINPUT22), .Z(n374) );
  XOR2_X1 U519 ( .A(KEYINPUT89), .B(KEYINPUT0), .Z(n375) );
  OR2_X1 U520 ( .A1(n639), .A2(n638), .ZN(n376) );
  XNOR2_X1 U521 ( .A(n543), .B(n387), .ZN(n752) );
  XOR2_X1 U522 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n377) );
  NOR2_X1 U523 ( .A1(n628), .A2(n556), .ZN(n684) );
  AND2_X1 U524 ( .A1(n564), .A2(n563), .ZN(n434) );
  NAND2_X1 U525 ( .A1(n398), .A2(n410), .ZN(n380) );
  NOR2_X1 U526 ( .A1(n381), .A2(KEYINPUT2), .ZN(n691) );
  NAND2_X1 U527 ( .A1(n368), .A2(n381), .ZN(n435) );
  XNOR2_X1 U528 ( .A(n381), .B(n759), .ZN(n761) );
  INV_X1 U529 ( .A(n771), .ZN(n382) );
  XNOR2_X1 U530 ( .A(n383), .B(G137), .ZN(G39) );
  NAND2_X1 U531 ( .A1(n695), .A2(n694), .ZN(n699) );
  INV_X1 U532 ( .A(n728), .ZN(n719) );
  NAND2_X1 U533 ( .A1(n390), .A2(n712), .ZN(n715) );
  XNOR2_X1 U534 ( .A(n390), .B(n618), .ZN(n620) );
  XNOR2_X2 U535 ( .A(n412), .B(n411), .ZN(n390) );
  INV_X1 U536 ( .A(n401), .ZN(n396) );
  NAND2_X1 U537 ( .A1(n444), .A2(n399), .ZN(n398) );
  NAND2_X1 U538 ( .A1(n401), .A2(n410), .ZN(n400) );
  NOR2_X2 U539 ( .A1(n727), .A2(n447), .ZN(n401) );
  NAND2_X1 U540 ( .A1(n427), .A2(n367), .ZN(n426) );
  NAND2_X1 U541 ( .A1(n601), .A2(n362), .ZN(n406) );
  XNOR2_X1 U542 ( .A(n442), .B(n422), .ZN(n427) );
  BUF_X1 U543 ( .A(n727), .Z(n407) );
  NAND2_X1 U544 ( .A1(n453), .A2(KEYINPUT78), .ZN(n452) );
  XNOR2_X1 U545 ( .A(n559), .B(n420), .ZN(n560) );
  NAND2_X1 U546 ( .A1(n441), .A2(n706), .ZN(n412) );
  XNOR2_X1 U547 ( .A(n431), .B(n377), .ZN(n464) );
  NAND2_X1 U548 ( .A1(n418), .A2(n769), .ZN(n442) );
  NAND2_X1 U549 ( .A1(n448), .A2(n372), .ZN(n417) );
  NOR2_X1 U550 ( .A1(n770), .A2(n443), .ZN(n418) );
  NAND2_X1 U551 ( .A1(n593), .A2(n432), .ZN(n431) );
  XNOR2_X1 U552 ( .A(n691), .B(KEYINPUT84), .ZN(n421) );
  NOR2_X1 U553 ( .A1(n434), .A2(n369), .ZN(n433) );
  XNOR2_X2 U554 ( .A(n426), .B(KEYINPUT45), .ZN(n749) );
  NAND2_X1 U555 ( .A1(n572), .A2(n571), .ZN(n429) );
  AND2_X1 U556 ( .A1(n428), .A2(n429), .ZN(n585) );
  INV_X1 U557 ( .A(n642), .ZN(n436) );
  NAND2_X1 U558 ( .A1(n598), .A2(n578), .ZN(n438) );
  NAND2_X1 U559 ( .A1(n440), .A2(n628), .ZN(n707) );
  INV_X1 U560 ( .A(n706), .ZN(n440) );
  NOR2_X1 U561 ( .A1(n594), .A2(n439), .ZN(n595) );
  NOR2_X1 U562 ( .A1(n615), .A2(n439), .ZN(n664) );
  INV_X1 U563 ( .A(n672), .ZN(n443) );
  NAND2_X1 U564 ( .A1(n727), .A2(n373), .ZN(n444) );
  XNOR2_X2 U565 ( .A(n622), .B(n621), .ZN(n727) );
  NAND2_X1 U566 ( .A1(n624), .A2(KEYINPUT78), .ZN(n450) );
  INV_X1 U567 ( .A(n624), .ZN(n448) );
  NOR2_X1 U568 ( .A1(n749), .A2(KEYINPUT2), .ZN(n690) );
  NAND2_X1 U569 ( .A1(n597), .A2(n694), .ZN(n457) );
  XNOR2_X2 U570 ( .A(n458), .B(n365), .ZN(n597) );
  NAND2_X1 U571 ( .A1(n647), .A2(n642), .ZN(n458) );
  XNOR2_X1 U572 ( .A(n459), .B(n731), .ZN(G75) );
  NAND2_X1 U573 ( .A1(n460), .A2(n371), .ZN(n459) );
  NAND2_X1 U574 ( .A1(n461), .A2(n404), .ZN(n460) );
  XNOR2_X1 U575 ( .A(n693), .B(KEYINPUT80), .ZN(n461) );
  XNOR2_X1 U576 ( .A(n473), .B(n482), .ZN(n474) );
  NOR2_X2 U577 ( .A1(G902), .A2(n732), .ZN(n476) );
  XOR2_X1 U578 ( .A(n520), .B(n519), .Z(n462) );
  AND2_X1 U579 ( .A1(G224), .A2(n760), .ZN(n463) );
  OR2_X1 U580 ( .A1(G953), .A2(n729), .ZN(n465) );
  INV_X1 U581 ( .A(KEYINPUT107), .ZN(n618) );
  INV_X1 U582 ( .A(KEYINPUT3), .ZN(n479) );
  INV_X1 U583 ( .A(n688), .ZN(n599) );
  NOR2_X1 U584 ( .A1(n689), .A2(n599), .ZN(n600) );
  XNOR2_X1 U585 ( .A(n489), .B(n488), .ZN(n490) );
  INV_X1 U586 ( .A(KEYINPUT87), .ZN(n575) );
  XNOR2_X1 U587 ( .A(n575), .B(KEYINPUT39), .ZN(n576) );
  INV_X1 U588 ( .A(KEYINPUT60), .ZN(n662) );
  XOR2_X1 U589 ( .A(KEYINPUT4), .B(G137), .Z(n466) );
  XNOR2_X1 U590 ( .A(G134), .B(n487), .ZN(n532) );
  NAND2_X1 U591 ( .A1(G227), .A2(n760), .ZN(n469) );
  XOR2_X1 U592 ( .A(n470), .B(n469), .Z(n473) );
  XOR2_X1 U593 ( .A(G110), .B(KEYINPUT75), .Z(n472) );
  XNOR2_X1 U594 ( .A(G107), .B(G104), .ZN(n471) );
  XNOR2_X1 U595 ( .A(KEYINPUT69), .B(G469), .ZN(n475) );
  XNOR2_X2 U596 ( .A(n476), .B(n475), .ZN(n565) );
  XNOR2_X1 U597 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U598 ( .A(n484), .B(n483), .ZN(n486) );
  XNOR2_X1 U599 ( .A(n500), .B(n463), .ZN(n485) );
  XNOR2_X1 U600 ( .A(n486), .B(n485), .ZN(n489) );
  INV_X1 U601 ( .A(n487), .ZN(n488) );
  INV_X1 U602 ( .A(n597), .ZN(n590) );
  XOR2_X1 U603 ( .A(n491), .B(KEYINPUT23), .Z(n495) );
  XOR2_X1 U604 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n493) );
  XNOR2_X1 U605 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U606 ( .A(n495), .B(n494), .ZN(n499) );
  NAND2_X1 U607 ( .A1(n760), .A2(G234), .ZN(n497) );
  XNOR2_X1 U608 ( .A(n497), .B(n496), .ZN(n529) );
  NAND2_X1 U609 ( .A1(G221), .A2(n529), .ZN(n498) );
  XNOR2_X1 U610 ( .A(n499), .B(n498), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n501), .B(KEYINPUT10), .ZN(n758) );
  XNOR2_X1 U612 ( .A(n502), .B(n758), .ZN(n744) );
  NOR2_X1 U613 ( .A1(n744), .A2(G902), .ZN(n503) );
  NAND2_X1 U614 ( .A1(n642), .A2(G234), .ZN(n504) );
  XNOR2_X1 U615 ( .A(KEYINPUT20), .B(n504), .ZN(n508) );
  NAND2_X1 U616 ( .A1(n508), .A2(G217), .ZN(n506) );
  INV_X1 U617 ( .A(KEYINPUT94), .ZN(n505) );
  INV_X1 U618 ( .A(n708), .ZN(n627) );
  XOR2_X1 U619 ( .A(KEYINPUT21), .B(KEYINPUT95), .Z(n510) );
  NAND2_X1 U620 ( .A1(n508), .A2(G221), .ZN(n509) );
  XNOR2_X1 U621 ( .A(n510), .B(n509), .ZN(n709) );
  XOR2_X1 U622 ( .A(KEYINPUT14), .B(n511), .Z(n726) );
  NAND2_X1 U623 ( .A1(n760), .A2(G952), .ZN(n602) );
  INV_X1 U624 ( .A(n602), .ZN(n513) );
  NOR2_X1 U625 ( .A1(G900), .A2(n607), .ZN(n512) );
  NOR2_X1 U626 ( .A1(n513), .A2(n512), .ZN(n514) );
  NOR2_X1 U627 ( .A1(n726), .A2(n514), .ZN(n573) );
  NAND2_X1 U628 ( .A1(n515), .A2(n573), .ZN(n558) );
  XNOR2_X1 U629 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U630 ( .A(n521), .B(G113), .ZN(n522) );
  NOR2_X1 U631 ( .A1(n655), .A2(G902), .ZN(n528) );
  XOR2_X1 U632 ( .A(KEYINPUT102), .B(KEYINPUT13), .Z(n526) );
  XNOR2_X1 U633 ( .A(KEYINPUT101), .B(G475), .ZN(n525) );
  XNOR2_X1 U634 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U635 ( .A(n528), .B(n527), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G217), .A2(n529), .ZN(n530) );
  XNOR2_X1 U637 ( .A(n531), .B(n530), .ZN(n537) );
  XOR2_X1 U638 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n535) );
  INV_X1 U639 ( .A(n532), .ZN(n534) );
  XNOR2_X1 U640 ( .A(n537), .B(n536), .ZN(n738) );
  NOR2_X1 U641 ( .A1(n738), .A2(G902), .ZN(n538) );
  XNOR2_X1 U642 ( .A(n538), .B(G478), .ZN(n587) );
  NAND2_X1 U643 ( .A1(n579), .A2(n587), .ZN(n539) );
  INV_X1 U644 ( .A(n678), .ZN(n551) );
  XOR2_X1 U645 ( .A(n541), .B(n540), .Z(n542) );
  XNOR2_X1 U646 ( .A(n543), .B(n542), .ZN(n546) );
  NAND2_X1 U647 ( .A1(n544), .A2(G210), .ZN(n545) );
  XNOR2_X1 U648 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U649 ( .A(n548), .B(n547), .ZN(n643) );
  NOR2_X1 U650 ( .A1(n643), .A2(G902), .ZN(n550) );
  INV_X1 U651 ( .A(G472), .ZN(n549) );
  XNOR2_X1 U652 ( .A(n550), .B(n549), .ZN(n566) );
  INV_X1 U653 ( .A(n566), .ZN(n631) );
  NAND2_X1 U654 ( .A1(n551), .A2(n619), .ZN(n552) );
  NOR2_X1 U655 ( .A1(n558), .A2(n552), .ZN(n554) );
  NAND2_X1 U656 ( .A1(G214), .A2(n553), .ZN(n694) );
  NAND2_X1 U657 ( .A1(n554), .A2(n694), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT36), .B(n555), .Z(n556) );
  INV_X1 U659 ( .A(n684), .ZN(n593) );
  OR2_X1 U660 ( .A1(n579), .A2(n587), .ZN(n557) );
  XNOR2_X1 U661 ( .A(n557), .B(KEYINPUT105), .ZN(n668) );
  NOR2_X1 U662 ( .A1(n668), .A2(n578), .ZN(n700) );
  INV_X1 U663 ( .A(n565), .ZN(n561) );
  NAND2_X1 U664 ( .A1(n580), .A2(n601), .ZN(n676) );
  XOR2_X1 U665 ( .A(n562), .B(KEYINPUT47), .Z(n564) );
  NAND2_X1 U666 ( .A1(n562), .A2(KEYINPUT81), .ZN(n563) );
  NAND2_X1 U667 ( .A1(n361), .A2(n706), .ZN(n630) );
  NAND2_X1 U668 ( .A1(n566), .A2(n694), .ZN(n569) );
  INV_X1 U669 ( .A(n569), .ZN(n568) );
  XOR2_X1 U670 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n570) );
  INV_X1 U671 ( .A(n570), .ZN(n567) );
  NAND2_X1 U672 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U673 ( .A1(n570), .A2(n569), .ZN(n571) );
  INV_X1 U674 ( .A(KEYINPUT38), .ZN(n574) );
  XNOR2_X1 U675 ( .A(n574), .B(n597), .ZN(n695) );
  INV_X1 U676 ( .A(n579), .ZN(n586) );
  NAND2_X1 U677 ( .A1(n586), .A2(n587), .ZN(n697) );
  AND2_X1 U678 ( .A1(n580), .A2(n719), .ZN(n581) );
  XNOR2_X1 U679 ( .A(n582), .B(KEYINPUT46), .ZN(n583) );
  NAND2_X1 U680 ( .A1(n700), .A2(KEYINPUT81), .ZN(n584) );
  NOR2_X1 U681 ( .A1(n676), .A2(n584), .ZN(n592) );
  NOR2_X1 U682 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U683 ( .A(n588), .B(KEYINPUT108), .ZN(n616) );
  NAND2_X1 U684 ( .A1(n585), .A2(n616), .ZN(n589) );
  NOR2_X1 U685 ( .A1(n590), .A2(n589), .ZN(n675) );
  XNOR2_X1 U686 ( .A(KEYINPUT82), .B(n675), .ZN(n591) );
  XNOR2_X1 U687 ( .A(n595), .B(KEYINPUT43), .ZN(n596) );
  NOR2_X1 U688 ( .A1(n597), .A2(n596), .ZN(n689) );
  NAND2_X1 U689 ( .A1(n598), .A2(n668), .ZN(n688) );
  INV_X1 U690 ( .A(n697), .ZN(n612) );
  OR2_X1 U691 ( .A1(G898), .A2(n607), .ZN(n603) );
  NAND2_X1 U692 ( .A1(n603), .A2(n602), .ZN(n605) );
  INV_X1 U693 ( .A(n726), .ZN(n604) );
  NAND2_X1 U694 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U695 ( .A1(KEYINPUT92), .A2(n606), .ZN(n611) );
  NOR2_X1 U696 ( .A1(n726), .A2(n607), .ZN(n609) );
  NOR2_X1 U697 ( .A1(G898), .A2(KEYINPUT92), .ZN(n608) );
  NAND2_X1 U698 ( .A1(n609), .A2(n608), .ZN(n610) );
  INV_X1 U699 ( .A(KEYINPUT73), .ZN(n613) );
  XNOR2_X1 U700 ( .A(n629), .B(KEYINPUT88), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n614), .A2(n627), .ZN(n615) );
  NAND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n622) );
  XNOR2_X1 U703 ( .A(KEYINPUT34), .B(KEYINPUT77), .ZN(n623) );
  INV_X1 U704 ( .A(n631), .ZN(n712) );
  OR2_X1 U705 ( .A1(n712), .A2(n624), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n627), .A2(n625), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n628), .A2(n626), .ZN(n672) );
  XNOR2_X1 U708 ( .A(n700), .B(KEYINPUT81), .ZN(n636) );
  NOR2_X1 U709 ( .A1(n633), .A2(n630), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n669) );
  NOR2_X1 U711 ( .A1(n633), .A2(n715), .ZN(n634) );
  XNOR2_X1 U712 ( .A(KEYINPUT31), .B(n634), .ZN(n681) );
  NAND2_X1 U713 ( .A1(n669), .A2(n681), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n637) );
  INV_X1 U715 ( .A(KEYINPUT2), .ZN(n639) );
  XOR2_X1 U716 ( .A(n642), .B(KEYINPUT85), .Z(n638) );
  INV_X1 U717 ( .A(KEYINPUT86), .ZN(n640) );
  INV_X1 U718 ( .A(n746), .ZN(n660) );
  NAND2_X1 U719 ( .A1(n645), .A2(n660), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U721 ( .A1(n742), .A2(G210), .ZN(n651) );
  XNOR2_X1 U722 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n647), .B(KEYINPUT55), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n652), .A2(n660), .ZN(n654) );
  INV_X1 U726 ( .A(KEYINPUT56), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(G51) );
  NAND2_X1 U728 ( .A1(n742), .A2(G475), .ZN(n659) );
  XOR2_X1 U729 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n657) );
  XNOR2_X1 U730 ( .A(n655), .B(KEYINPUT64), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n659), .B(n658), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(G60) );
  XOR2_X1 U734 ( .A(G101), .B(n664), .Z(G3) );
  NOR2_X1 U735 ( .A1(n678), .A2(n669), .ZN(n665) );
  XOR2_X1 U736 ( .A(G104), .B(n665), .Z(G6) );
  XOR2_X1 U737 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n667) );
  XNOR2_X1 U738 ( .A(G107), .B(KEYINPUT112), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(n671) );
  INV_X1 U740 ( .A(n668), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n682), .A2(n669), .ZN(n670) );
  XOR2_X1 U742 ( .A(n671), .B(n670), .Z(G9) );
  XNOR2_X1 U743 ( .A(n672), .B(G110), .ZN(G12) );
  NOR2_X1 U744 ( .A1(n676), .A2(n682), .ZN(n674) );
  XNOR2_X1 U745 ( .A(G128), .B(KEYINPUT29), .ZN(n673) );
  XNOR2_X1 U746 ( .A(n674), .B(n673), .ZN(G30) );
  XOR2_X1 U747 ( .A(G143), .B(n675), .Z(G45) );
  NOR2_X1 U748 ( .A1(n678), .A2(n676), .ZN(n677) );
  XOR2_X1 U749 ( .A(G146), .B(n677), .Z(G48) );
  NOR2_X1 U750 ( .A1(n678), .A2(n681), .ZN(n680) );
  XNOR2_X1 U751 ( .A(G113), .B(KEYINPUT113), .ZN(n679) );
  XNOR2_X1 U752 ( .A(n680), .B(n679), .ZN(G15) );
  NOR2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U754 ( .A(G116), .B(n683), .Z(G18) );
  XNOR2_X1 U755 ( .A(n684), .B(KEYINPUT37), .ZN(n685) );
  XNOR2_X1 U756 ( .A(n685), .B(KEYINPUT114), .ZN(n686) );
  XNOR2_X1 U757 ( .A(G125), .B(n686), .ZN(G27) );
  XOR2_X1 U758 ( .A(G134), .B(KEYINPUT115), .Z(n687) );
  XNOR2_X1 U759 ( .A(n688), .B(n687), .ZN(G36) );
  XOR2_X1 U760 ( .A(G140), .B(n689), .Z(G42) );
  XOR2_X1 U761 ( .A(KEYINPUT83), .B(n690), .Z(n692) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U764 ( .A(KEYINPUT117), .B(n698), .Z(n703) );
  NOR2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U766 ( .A(KEYINPUT118), .B(n701), .ZN(n702) );
  NOR2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U768 ( .A1(n704), .A2(n407), .ZN(n705) );
  XNOR2_X1 U769 ( .A(n705), .B(KEYINPUT119), .ZN(n722) );
  XNOR2_X1 U770 ( .A(n707), .B(KEYINPUT50), .ZN(n714) );
  NAND2_X1 U771 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U772 ( .A(KEYINPUT49), .B(n710), .ZN(n711) );
  NOR2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U774 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U775 ( .A1(n716), .A2(n715), .ZN(n718) );
  XOR2_X1 U776 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n717) );
  XNOR2_X1 U777 ( .A(n718), .B(n717), .ZN(n720) );
  NAND2_X1 U778 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U779 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U780 ( .A(KEYINPUT52), .B(n723), .ZN(n724) );
  NAND2_X1 U781 ( .A1(n724), .A2(G952), .ZN(n725) );
  NOR2_X1 U782 ( .A1(n726), .A2(n725), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n728), .A2(n407), .ZN(n729) );
  XOR2_X1 U784 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n731) );
  XNOR2_X1 U785 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n734) );
  XNOR2_X1 U786 ( .A(n732), .B(KEYINPUT57), .ZN(n733) );
  XNOR2_X1 U787 ( .A(n734), .B(n733), .ZN(n736) );
  NAND2_X1 U788 ( .A1(n742), .A2(G469), .ZN(n735) );
  XOR2_X1 U789 ( .A(n736), .B(n735), .Z(n737) );
  NOR2_X1 U790 ( .A1(n746), .A2(n737), .ZN(G54) );
  XNOR2_X1 U791 ( .A(n738), .B(KEYINPUT124), .ZN(n740) );
  NAND2_X1 U792 ( .A1(G478), .A2(n742), .ZN(n739) );
  XNOR2_X1 U793 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U794 ( .A1(n746), .A2(n741), .ZN(G63) );
  NAND2_X1 U795 ( .A1(G217), .A2(n742), .ZN(n743) );
  XNOR2_X1 U796 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n746), .A2(n745), .ZN(G66) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n747) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n747), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n748), .A2(G898), .ZN(n751) );
  NAND2_X1 U801 ( .A1(n749), .A2(n760), .ZN(n750) );
  NAND2_X1 U802 ( .A1(n751), .A2(n750), .ZN(n756) );
  XNOR2_X1 U803 ( .A(KEYINPUT125), .B(n752), .ZN(n754) );
  OR2_X1 U804 ( .A1(n760), .A2(G898), .ZN(n753) );
  NAND2_X1 U805 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U806 ( .A(n756), .B(n755), .Z(G69) );
  XNOR2_X1 U807 ( .A(n757), .B(n758), .ZN(n762) );
  INV_X1 U808 ( .A(n762), .ZN(n759) );
  NAND2_X1 U809 ( .A1(n761), .A2(n760), .ZN(n768) );
  XNOR2_X1 U810 ( .A(n762), .B(G227), .ZN(n763) );
  XNOR2_X1 U811 ( .A(n763), .B(KEYINPUT126), .ZN(n764) );
  NAND2_X1 U812 ( .A1(n764), .A2(G900), .ZN(n765) );
  NAND2_X1 U813 ( .A1(G953), .A2(n765), .ZN(n766) );
  XOR2_X1 U814 ( .A(KEYINPUT127), .B(n766), .Z(n767) );
  NAND2_X1 U815 ( .A1(n768), .A2(n767), .ZN(G72) );
  XNOR2_X1 U816 ( .A(n769), .B(G122), .ZN(G24) );
  XOR2_X1 U817 ( .A(n770), .B(G119), .Z(G21) );
  XOR2_X1 U818 ( .A(G131), .B(n771), .Z(G33) );
endmodule

