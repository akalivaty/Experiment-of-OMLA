

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(G2104), .A2(n520), .ZN(n903) );
  NAND2_X2 U555 ( .A1(G160), .A2(G40), .ZN(n714) );
  NOR2_X2 U556 ( .A1(n639), .A2(n544), .ZN(n654) );
  NOR2_X2 U557 ( .A1(n538), .A2(n537), .ZN(G160) );
  NAND2_X1 U558 ( .A1(n521), .A2(n520), .ZN(n522) );
  INV_X1 U559 ( .A(G2104), .ZN(n521) );
  INV_X1 U560 ( .A(KEYINPUT97), .ZN(n742) );
  NOR2_X1 U561 ( .A1(n766), .A2(n874), .ZN(n725) );
  INV_X1 U562 ( .A(n775), .ZN(n755) );
  NAND2_X1 U563 ( .A1(n755), .A2(G8), .ZN(n756) );
  NOR2_X1 U564 ( .A1(n760), .A2(n759), .ZN(n761) );
  INV_X1 U565 ( .A(KEYINPUT99), .ZN(n764) );
  INV_X1 U566 ( .A(KEYINPUT32), .ZN(n773) );
  NAND2_X2 U567 ( .A1(n718), .A2(n717), .ZN(n766) );
  XNOR2_X1 U568 ( .A(n754), .B(KEYINPUT93), .ZN(n808) );
  INV_X1 U569 ( .A(G2105), .ZN(n520) );
  AND2_X2 U570 ( .A1(n520), .A2(G2104), .ZN(n908) );
  XNOR2_X1 U571 ( .A(n566), .B(KEYINPUT71), .ZN(n568) );
  NOR2_X1 U572 ( .A1(G651), .A2(n639), .ZN(n647) );
  NAND2_X1 U573 ( .A1(n568), .A2(n567), .ZN(n968) );
  OR2_X1 U574 ( .A1(n531), .A2(n530), .ZN(n718) );
  INV_X1 U575 ( .A(n718), .ZN(G164) );
  XNOR2_X2 U576 ( .A(n522), .B(KEYINPUT17), .ZN(n906) );
  NAND2_X1 U577 ( .A1(G138), .A2(n906), .ZN(n524) );
  NAND2_X1 U578 ( .A1(G102), .A2(n908), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U580 ( .A(KEYINPUT87), .B(n525), .Z(n531) );
  NAND2_X1 U581 ( .A1(G126), .A2(n903), .ZN(n528) );
  NAND2_X1 U582 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XNOR2_X1 U583 ( .A(n526), .B(KEYINPUT65), .ZN(n607) );
  NAND2_X1 U584 ( .A1(G114), .A2(n607), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U586 ( .A(KEYINPUT86), .B(n529), .ZN(n530) );
  NAND2_X1 U587 ( .A1(n906), .A2(G137), .ZN(n534) );
  NAND2_X1 U588 ( .A1(G101), .A2(n908), .ZN(n532) );
  XOR2_X1 U589 ( .A(KEYINPUT23), .B(n532), .Z(n533) );
  NAND2_X1 U590 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G125), .A2(n903), .ZN(n536) );
  NAND2_X1 U592 ( .A1(G113), .A2(n607), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X2 U594 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U595 ( .A1(G90), .A2(n645), .ZN(n540) );
  XOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .Z(n639) );
  INV_X1 U597 ( .A(G651), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G77), .A2(n654), .ZN(n539) );
  NAND2_X1 U599 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U600 ( .A(n541), .B(KEYINPUT9), .ZN(n543) );
  NAND2_X1 U601 ( .A1(G52), .A2(n647), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n548) );
  NOR2_X1 U603 ( .A1(G543), .A2(n544), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT1), .B(n545), .Z(n558) );
  BUF_X1 U605 ( .A(n558), .Z(n648) );
  NAND2_X1 U606 ( .A1(n648), .A2(G64), .ZN(n546) );
  XOR2_X1 U607 ( .A(KEYINPUT68), .B(n546), .Z(n547) );
  NOR2_X1 U608 ( .A1(n548), .A2(n547), .ZN(G171) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U610 ( .A(G57), .ZN(G237) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  NAND2_X1 U612 ( .A1(G91), .A2(n645), .ZN(n550) );
  NAND2_X1 U613 ( .A1(G65), .A2(n648), .ZN(n549) );
  NAND2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G53), .A2(n647), .ZN(n551) );
  XNOR2_X1 U616 ( .A(KEYINPUT69), .B(n551), .ZN(n552) );
  NOR2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n654), .A2(G78), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(G299) );
  NAND2_X1 U620 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U622 ( .A(G223), .ZN(n834) );
  NAND2_X1 U623 ( .A1(n834), .A2(G567), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  NAND2_X1 U625 ( .A1(n558), .A2(G56), .ZN(n559) );
  XNOR2_X1 U626 ( .A(KEYINPUT14), .B(n559), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n645), .A2(G81), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(KEYINPUT12), .ZN(n562) );
  NAND2_X1 U629 ( .A1(G68), .A2(n654), .ZN(n561) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(KEYINPUT13), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n647), .A2(G43), .ZN(n567) );
  INV_X1 U634 ( .A(n968), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G860), .B(KEYINPUT72), .ZN(n594) );
  NAND2_X1 U636 ( .A1(n569), .A2(n594), .ZN(G153) );
  XNOR2_X1 U637 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U638 ( .A1(G868), .A2(G301), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G92), .A2(n645), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G66), .A2(n648), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G79), .A2(n654), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G54), .A2(n647), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U646 ( .A(KEYINPUT15), .B(n576), .Z(n961) );
  INV_X1 U647 ( .A(n961), .ZN(n597) );
  INV_X1 U648 ( .A(G868), .ZN(n665) );
  NAND2_X1 U649 ( .A1(n597), .A2(n665), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n578), .A2(n577), .ZN(G284) );
  NAND2_X1 U651 ( .A1(n647), .A2(G51), .ZN(n579) );
  XOR2_X1 U652 ( .A(KEYINPUT75), .B(n579), .Z(n581) );
  NAND2_X1 U653 ( .A1(n648), .A2(G63), .ZN(n580) );
  NAND2_X1 U654 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U655 ( .A(KEYINPUT6), .B(n582), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n654), .A2(G76), .ZN(n583) );
  XNOR2_X1 U657 ( .A(KEYINPUT74), .B(n583), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n645), .A2(G89), .ZN(n584) );
  XNOR2_X1 U659 ( .A(KEYINPUT4), .B(n584), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U661 ( .A(n587), .B(KEYINPUT5), .Z(n588) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U663 ( .A(KEYINPUT7), .B(n590), .Z(n591) );
  XNOR2_X1 U664 ( .A(KEYINPUT76), .B(n591), .ZN(G168) );
  XOR2_X1 U665 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U666 ( .A1(G868), .A2(G286), .ZN(n593) );
  NAND2_X1 U667 ( .A1(G299), .A2(n665), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(G297) );
  INV_X1 U669 ( .A(G559), .ZN(n595) );
  NOR2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U672 ( .A(KEYINPUT16), .B(n598), .Z(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n968), .ZN(n601) );
  NAND2_X1 U674 ( .A1(G868), .A2(n961), .ZN(n599) );
  NOR2_X1 U675 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U677 ( .A1(G135), .A2(n906), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT78), .ZN(n606) );
  XOR2_X1 U679 ( .A(KEYINPUT18), .B(KEYINPUT77), .Z(n604) );
  NAND2_X1 U680 ( .A1(G123), .A2(n903), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n604), .B(n603), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G111), .A2(n607), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G99), .A2(n908), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n932) );
  XOR2_X1 U687 ( .A(G2096), .B(n932), .Z(n612) );
  NOR2_X1 U688 ( .A1(G2100), .A2(n612), .ZN(n613) );
  XNOR2_X1 U689 ( .A(KEYINPUT79), .B(n613), .ZN(G156) );
  NAND2_X1 U690 ( .A1(G559), .A2(n961), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n614), .B(KEYINPUT80), .ZN(n663) );
  XNOR2_X1 U692 ( .A(n663), .B(n968), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n615), .A2(G860), .ZN(n623) );
  NAND2_X1 U694 ( .A1(n648), .A2(G67), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G93), .A2(n645), .ZN(n616) );
  XOR2_X1 U696 ( .A(KEYINPUT81), .B(n616), .Z(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G80), .A2(n654), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G55), .A2(n647), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n666) );
  XOR2_X1 U702 ( .A(n623), .B(n666), .Z(G145) );
  NAND2_X1 U703 ( .A1(G75), .A2(n654), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G50), .A2(n647), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G88), .A2(n645), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G62), .A2(n648), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U710 ( .A(n630), .B(KEYINPUT83), .ZN(G303) );
  INV_X1 U711 ( .A(G303), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G86), .A2(n645), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G61), .A2(n648), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n654), .A2(G73), .ZN(n633) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n647), .A2(G48), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U720 ( .A1(G49), .A2(n647), .ZN(n638) );
  XNOR2_X1 U721 ( .A(n638), .B(KEYINPUT82), .ZN(n644) );
  NAND2_X1 U722 ( .A1(G87), .A2(n639), .ZN(n641) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U725 ( .A1(n648), .A2(n642), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(G288) );
  NAND2_X1 U727 ( .A1(G85), .A2(n645), .ZN(n646) );
  XOR2_X1 U728 ( .A(KEYINPUT66), .B(n646), .Z(n653) );
  NAND2_X1 U729 ( .A1(G47), .A2(n647), .ZN(n650) );
  NAND2_X1 U730 ( .A1(G60), .A2(n648), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U732 ( .A(KEYINPUT67), .B(n651), .Z(n652) );
  NOR2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n654), .A2(G72), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n656), .A2(n655), .ZN(G290) );
  XNOR2_X1 U736 ( .A(G166), .B(n968), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n657), .B(G305), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n658), .B(G299), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n659), .B(G288), .ZN(n660) );
  XOR2_X1 U740 ( .A(n666), .B(n660), .Z(n662) );
  XNOR2_X1 U741 ( .A(G290), .B(KEYINPUT19), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n662), .B(n661), .ZN(n917) );
  XOR2_X1 U743 ( .A(n917), .B(n663), .Z(n664) );
  NOR2_X1 U744 ( .A1(n665), .A2(n664), .ZN(n668) );
  NOR2_X1 U745 ( .A1(G868), .A2(n666), .ZN(n667) );
  NOR2_X1 U746 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2084), .A2(G2078), .ZN(n669) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U749 ( .A1(n670), .A2(G2090), .ZN(n671) );
  XNOR2_X1 U750 ( .A(n671), .B(KEYINPUT21), .ZN(n672) );
  XNOR2_X1 U751 ( .A(KEYINPUT84), .B(n672), .ZN(n673) );
  NAND2_X1 U752 ( .A1(G2072), .A2(n673), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U754 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U757 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U758 ( .A1(G96), .A2(n676), .ZN(n838) );
  NAND2_X1 U759 ( .A1(n838), .A2(G2106), .ZN(n680) );
  NAND2_X1 U760 ( .A1(G69), .A2(G120), .ZN(n677) );
  NOR2_X1 U761 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U762 ( .A1(G108), .A2(n678), .ZN(n839) );
  NAND2_X1 U763 ( .A1(n839), .A2(G567), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n680), .A2(n679), .ZN(n853) );
  NAND2_X1 U765 ( .A1(G661), .A2(G483), .ZN(n681) );
  NOR2_X1 U766 ( .A1(n853), .A2(n681), .ZN(n837) );
  NAND2_X1 U767 ( .A1(n837), .A2(G36), .ZN(n682) );
  XOR2_X1 U768 ( .A(KEYINPUT85), .B(n682), .Z(G176) );
  NAND2_X1 U769 ( .A1(G140), .A2(n906), .ZN(n684) );
  NAND2_X1 U770 ( .A1(G104), .A2(n908), .ZN(n683) );
  NAND2_X1 U771 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n685), .ZN(n690) );
  NAND2_X1 U773 ( .A1(G128), .A2(n903), .ZN(n687) );
  NAND2_X1 U774 ( .A1(G116), .A2(n607), .ZN(n686) );
  NAND2_X1 U775 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U776 ( .A(KEYINPUT35), .B(n688), .Z(n689) );
  NOR2_X1 U777 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U778 ( .A(KEYINPUT36), .B(n691), .ZN(n895) );
  XNOR2_X1 U779 ( .A(KEYINPUT37), .B(G2067), .ZN(n826) );
  NOR2_X1 U780 ( .A1(n895), .A2(n826), .ZN(n930) );
  INV_X1 U781 ( .A(G1384), .ZN(n715) );
  AND2_X1 U782 ( .A1(n718), .A2(n715), .ZN(n692) );
  NOR2_X1 U783 ( .A1(n692), .A2(n714), .ZN(n828) );
  NAND2_X1 U784 ( .A1(n930), .A2(n828), .ZN(n825) );
  NAND2_X1 U785 ( .A1(n607), .A2(G107), .ZN(n699) );
  NAND2_X1 U786 ( .A1(G119), .A2(n903), .ZN(n694) );
  NAND2_X1 U787 ( .A1(G95), .A2(n908), .ZN(n693) );
  NAND2_X1 U788 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n906), .A2(G131), .ZN(n695) );
  XOR2_X1 U790 ( .A(KEYINPUT88), .B(n695), .Z(n696) );
  NOR2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U793 ( .A(KEYINPUT89), .B(n700), .ZN(n900) );
  XOR2_X1 U794 ( .A(KEYINPUT90), .B(G1991), .Z(n1018) );
  NOR2_X1 U795 ( .A1(n900), .A2(n1018), .ZN(n711) );
  XOR2_X1 U796 ( .A(KEYINPUT38), .B(KEYINPUT91), .Z(n702) );
  NAND2_X1 U797 ( .A1(G105), .A2(n908), .ZN(n701) );
  XNOR2_X1 U798 ( .A(n702), .B(n701), .ZN(n709) );
  NAND2_X1 U799 ( .A1(G129), .A2(n903), .ZN(n704) );
  NAND2_X1 U800 ( .A1(G117), .A2(n607), .ZN(n703) );
  NAND2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n906), .A2(G141), .ZN(n705) );
  XOR2_X1 U803 ( .A(KEYINPUT92), .B(n705), .Z(n706) );
  NOR2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n899) );
  AND2_X1 U806 ( .A1(n899), .A2(G1996), .ZN(n710) );
  NOR2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n934) );
  INV_X1 U808 ( .A(n828), .ZN(n712) );
  NOR2_X1 U809 ( .A1(n934), .A2(n712), .ZN(n820) );
  INV_X1 U810 ( .A(n820), .ZN(n713) );
  NAND2_X1 U811 ( .A1(n825), .A2(n713), .ZN(n815) );
  INV_X1 U812 ( .A(n714), .ZN(n716) );
  AND2_X1 U813 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X2 U814 ( .A(KEYINPUT95), .B(n766), .ZN(n747) );
  NAND2_X1 U815 ( .A1(n747), .A2(G2072), .ZN(n720) );
  XOR2_X1 U816 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n719) );
  XNOR2_X1 U817 ( .A(n720), .B(n719), .ZN(n739) );
  INV_X1 U818 ( .A(n747), .ZN(n721) );
  NAND2_X1 U819 ( .A1(n721), .A2(G1956), .ZN(n736) );
  NAND2_X1 U820 ( .A1(n739), .A2(n736), .ZN(n722) );
  NAND2_X1 U821 ( .A1(G299), .A2(n722), .ZN(n723) );
  XOR2_X1 U822 ( .A(KEYINPUT28), .B(n723), .Z(n745) );
  INV_X1 U823 ( .A(G1996), .ZN(n874) );
  XOR2_X1 U824 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n724) );
  XNOR2_X1 U825 ( .A(n725), .B(n724), .ZN(n728) );
  AND2_X1 U826 ( .A1(n766), .A2(G1341), .ZN(n726) );
  NOR2_X1 U827 ( .A1(n726), .A2(n968), .ZN(n727) );
  AND2_X2 U828 ( .A1(n728), .A2(n727), .ZN(n733) );
  NAND2_X1 U829 ( .A1(n733), .A2(n961), .ZN(n732) );
  NAND2_X1 U830 ( .A1(G1348), .A2(n766), .ZN(n730) );
  NAND2_X1 U831 ( .A1(G2067), .A2(n747), .ZN(n729) );
  NAND2_X1 U832 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U833 ( .A1(n732), .A2(n731), .ZN(n735) );
  OR2_X1 U834 ( .A1(n961), .A2(n733), .ZN(n734) );
  AND2_X1 U835 ( .A1(n735), .A2(n734), .ZN(n741) );
  INV_X1 U836 ( .A(n736), .ZN(n737) );
  NOR2_X1 U837 ( .A1(G299), .A2(n737), .ZN(n738) );
  AND2_X1 U838 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U839 ( .A1(n741), .A2(n740), .ZN(n743) );
  XNOR2_X1 U840 ( .A(n743), .B(n742), .ZN(n744) );
  NOR2_X1 U841 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U842 ( .A(n746), .B(KEYINPUT29), .ZN(n751) );
  INV_X1 U843 ( .A(G1961), .ZN(n995) );
  NAND2_X1 U844 ( .A1(n995), .A2(n766), .ZN(n749) );
  XNOR2_X1 U845 ( .A(G2078), .B(KEYINPUT25), .ZN(n1006) );
  NAND2_X1 U846 ( .A1(n747), .A2(n1006), .ZN(n748) );
  NAND2_X1 U847 ( .A1(n749), .A2(n748), .ZN(n753) );
  NAND2_X1 U848 ( .A1(G171), .A2(n753), .ZN(n750) );
  NAND2_X1 U849 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U850 ( .A(n752), .B(KEYINPUT98), .ZN(n763) );
  NOR2_X1 U851 ( .A1(G171), .A2(n753), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n766), .A2(G8), .ZN(n754) );
  INV_X1 U853 ( .A(n808), .ZN(n796) );
  NOR2_X1 U854 ( .A1(G1966), .A2(n796), .ZN(n780) );
  NOR2_X1 U855 ( .A1(G2084), .A2(n766), .ZN(n775) );
  OR2_X1 U856 ( .A1(n780), .A2(n756), .ZN(n757) );
  XNOR2_X1 U857 ( .A(KEYINPUT30), .B(n757), .ZN(n758) );
  NOR2_X1 U858 ( .A1(n758), .A2(G168), .ZN(n759) );
  XOR2_X1 U859 ( .A(KEYINPUT31), .B(n761), .Z(n762) );
  NAND2_X1 U860 ( .A1(n763), .A2(n762), .ZN(n778) );
  NAND2_X1 U861 ( .A1(n778), .A2(G286), .ZN(n765) );
  XNOR2_X1 U862 ( .A(n765), .B(n764), .ZN(n771) );
  NOR2_X1 U863 ( .A1(G1971), .A2(n796), .ZN(n768) );
  NOR2_X1 U864 ( .A1(G2090), .A2(n766), .ZN(n767) );
  NOR2_X1 U865 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U866 ( .A1(G303), .A2(n769), .ZN(n770) );
  NAND2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U868 ( .A1(n772), .A2(G8), .ZN(n774) );
  XNOR2_X1 U869 ( .A(n774), .B(n773), .ZN(n791) );
  NAND2_X1 U870 ( .A1(G8), .A2(n775), .ZN(n776) );
  XNOR2_X1 U871 ( .A(n776), .B(KEYINPUT94), .ZN(n777) );
  NAND2_X1 U872 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n787) );
  NOR2_X1 U874 ( .A1(n791), .A2(n787), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G166), .A2(G8), .ZN(n781) );
  NOR2_X1 U876 ( .A1(G2090), .A2(n781), .ZN(n782) );
  NOR2_X1 U877 ( .A1(n783), .A2(n782), .ZN(n785) );
  INV_X1 U878 ( .A(KEYINPUT101), .ZN(n784) );
  XNOR2_X1 U879 ( .A(n785), .B(n784), .ZN(n786) );
  NOR2_X1 U880 ( .A1(n786), .A2(n808), .ZN(n813) );
  NAND2_X1 U881 ( .A1(G1976), .A2(G288), .ZN(n957) );
  INV_X1 U882 ( .A(n957), .ZN(n794) );
  OR2_X2 U883 ( .A1(n787), .A2(n794), .ZN(n788) );
  OR2_X1 U884 ( .A1(n788), .A2(n796), .ZN(n789) );
  XNOR2_X1 U885 ( .A(G1981), .B(G305), .ZN(n970) );
  OR2_X2 U886 ( .A1(n789), .A2(n970), .ZN(n790) );
  NOR2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n802) );
  INV_X1 U888 ( .A(n970), .ZN(n800) );
  NOR2_X1 U889 ( .A1(G1976), .A2(G288), .ZN(n803) );
  NOR2_X1 U890 ( .A1(G1971), .A2(G303), .ZN(n792) );
  NOR2_X1 U891 ( .A1(n803), .A2(n792), .ZN(n965) );
  XNOR2_X1 U892 ( .A(KEYINPUT100), .B(n965), .ZN(n793) );
  OR2_X1 U893 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U894 ( .A1(n796), .A2(n795), .ZN(n798) );
  INV_X1 U895 ( .A(KEYINPUT33), .ZN(n797) );
  NAND2_X1 U896 ( .A1(n798), .A2(n797), .ZN(n799) );
  AND2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n806) );
  AND2_X1 U899 ( .A1(n803), .A2(KEYINPUT33), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n804), .A2(n808), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n811) );
  NOR2_X1 U902 ( .A1(G1981), .A2(G305), .ZN(n807) );
  XNOR2_X1 U903 ( .A(n807), .B(KEYINPUT24), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n817) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n956) );
  NAND2_X1 U909 ( .A1(n956), .A2(n828), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n832) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n899), .ZN(n944) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n818) );
  AND2_X1 U913 ( .A1(n900), .A2(n1018), .ZN(n936) );
  NOR2_X1 U914 ( .A1(n818), .A2(n936), .ZN(n819) );
  NOR2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n944), .A2(n821), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT39), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n823), .B(KEYINPUT102), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n895), .A2(n826), .ZN(n928) );
  NAND2_X1 U921 ( .A1(n827), .A2(n928), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U923 ( .A(KEYINPUT103), .B(n830), .Z(n831) );
  NAND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U925 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U928 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U937 ( .A(G1341), .B(G1348), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n840), .B(G2427), .ZN(n850) );
  XOR2_X1 U939 ( .A(KEYINPUT106), .B(G2430), .Z(n842) );
  XNOR2_X1 U940 ( .A(G2446), .B(G2451), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U942 ( .A(KEYINPUT105), .B(G2435), .Z(n844) );
  XNOR2_X1 U943 ( .A(G2438), .B(G2454), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U945 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U946 ( .A(KEYINPUT104), .B(G2443), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n851), .A2(G14), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n852), .B(KEYINPUT107), .ZN(G401) );
  INV_X1 U951 ( .A(n853), .ZN(G319) );
  XOR2_X1 U952 ( .A(G2678), .B(KEYINPUT110), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2100), .B(KEYINPUT43), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n856), .B(G2096), .Z(n858) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2078), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U958 ( .A(KEYINPUT109), .B(G2090), .Z(n860) );
  XNOR2_X1 U959 ( .A(G2084), .B(G2072), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U961 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U962 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(G227) );
  XOR2_X1 U964 ( .A(G1981), .B(G1961), .Z(n866) );
  XNOR2_X1 U965 ( .A(G1991), .B(G1966), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U967 ( .A(G1986), .B(G1976), .Z(n868) );
  XNOR2_X1 U968 ( .A(G1956), .B(G1971), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U971 ( .A(KEYINPUT111), .B(G2474), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT41), .B(n873), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(G229) );
  NAND2_X1 U975 ( .A1(G124), .A2(n903), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n876), .B(KEYINPUT112), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n877), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G136), .A2(n906), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G112), .A2(n607), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G100), .A2(n908), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(KEYINPUT113), .B(n884), .Z(G162) );
  NAND2_X1 U985 ( .A1(G139), .A2(n906), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G103), .A2(n908), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n891) );
  NAND2_X1 U988 ( .A1(G127), .A2(n903), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G115), .A2(n607), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n939) );
  XOR2_X1 U993 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n893) );
  XNOR2_X1 U994 ( .A(G160), .B(G162), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n939), .B(n894), .ZN(n897) );
  XNOR2_X1 U997 ( .A(G164), .B(n895), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U999 ( .A(n898), .B(n932), .Z(n902) );
  XOR2_X1 U1000 ( .A(n900), .B(n899), .Z(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n915) );
  NAND2_X1 U1002 ( .A1(G130), .A2(n903), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(G118), .A2(n607), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(n906), .A2(G142), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n907), .B(KEYINPUT114), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(G106), .A2(n908), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(KEYINPUT45), .B(n911), .Z(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n916), .ZN(G395) );
  XOR2_X1 U1013 ( .A(KEYINPUT115), .B(n917), .Z(n919) );
  XNOR2_X1 U1014 ( .A(G171), .B(n961), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(n920), .B(G286), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n921), .ZN(G397) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n922) );
  XOR2_X1 U1019 ( .A(KEYINPUT49), .B(n922), .Z(n923) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n923), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G401), .A2(n924), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT116), .B(n925), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G108), .ZN(G238) );
  INV_X1 U1027 ( .A(n928), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n938) );
  XOR2_X1 U1029 ( .A(G2084), .B(G160), .Z(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n949) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n941) );
  INV_X1 U1035 ( .A(G2072), .ZN(n1011) );
  XNOR2_X1 U1036 ( .A(n1011), .B(n939), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(KEYINPUT50), .B(n942), .ZN(n947) );
  XOR2_X1 U1039 ( .A(G2090), .B(G162), .Z(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1041 ( .A(KEYINPUT51), .B(n945), .Z(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT52), .B(n950), .ZN(n952) );
  INV_X1 U1045 ( .A(KEYINPUT55), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n953), .A2(G29), .ZN(n1037) );
  INV_X1 U1048 ( .A(G16), .ZN(n1003) );
  XNOR2_X1 U1049 ( .A(KEYINPUT56), .B(KEYINPUT123), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(n1003), .B(n954), .ZN(n977) );
  XNOR2_X1 U1051 ( .A(G1956), .B(G299), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n967) );
  XNOR2_X1 U1054 ( .A(G171), .B(G1961), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(G1971), .A2(G303), .ZN(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1057 ( .A(n961), .B(G1348), .Z(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n975) );
  XNOR2_X1 U1061 ( .A(n968), .B(G1341), .ZN(n973) );
  XOR2_X1 U1062 ( .A(G1966), .B(G168), .Z(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(KEYINPUT57), .B(n971), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n1005) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G22), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(G23), .B(G1976), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n981) );
  XOR2_X1 U1071 ( .A(G1986), .B(G24), .Z(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n983) );
  XOR2_X1 U1073 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n982) );
  XNOR2_X1 U1074 ( .A(n983), .B(n982), .ZN(n1000) );
  XOR2_X1 U1075 ( .A(G1966), .B(G21), .Z(n994) );
  XOR2_X1 U1076 ( .A(G1348), .B(KEYINPUT59), .Z(n984) );
  XNOR2_X1 U1077 ( .A(G4), .B(n984), .ZN(n991) );
  XOR2_X1 U1078 ( .A(G1981), .B(G6), .Z(n988) );
  XNOR2_X1 U1079 ( .A(G1341), .B(G19), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(G1956), .B(G20), .ZN(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1083 ( .A(KEYINPUT125), .B(n989), .Z(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(KEYINPUT60), .B(n992), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n998) );
  XOR2_X1 U1087 ( .A(G5), .B(n995), .Z(n996) );
  XNOR2_X1 U1088 ( .A(KEYINPUT124), .B(n996), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1091 ( .A(KEYINPUT61), .B(n1001), .Z(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1035) );
  XNOR2_X1 U1094 ( .A(G27), .B(KEYINPUT119), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1007), .B(n1006), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G32), .B(G1996), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT120), .B(n1010), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(G33), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(G28), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(KEYINPUT118), .B(G2067), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G26), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(KEYINPUT117), .B(n1018), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(G25), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1108 ( .A(KEYINPUT53), .B(n1022), .Z(n1026) );
  XNOR2_X1 U1109 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(n1023), .B(G34), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(G2084), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(G35), .B(G2090), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1115 ( .A(n1029), .B(KEYINPUT55), .ZN(n1031) );
  INV_X1 U1116 ( .A(G29), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(G11), .A2(n1032), .ZN(n1033) );
  XNOR2_X1 U1119 ( .A(KEYINPUT122), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1122 ( .A(n1038), .B(KEYINPUT62), .ZN(n1039) );
  XNOR2_X1 U1123 ( .A(KEYINPUT127), .B(n1039), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

