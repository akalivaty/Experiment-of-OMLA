

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714;

  XNOR2_X1 U364 ( .A(n413), .B(G469), .ZN(n524) );
  XNOR2_X2 U365 ( .A(n481), .B(n480), .ZN(n711) );
  XNOR2_X2 U366 ( .A(n467), .B(KEYINPUT35), .ZN(n714) );
  XNOR2_X2 U367 ( .A(n363), .B(G143), .ZN(n460) );
  XNOR2_X2 U368 ( .A(G128), .B(KEYINPUT64), .ZN(n363) );
  AND2_X1 U369 ( .A1(n353), .A2(n345), .ZN(n352) );
  XNOR2_X1 U370 ( .A(n359), .B(KEYINPUT40), .ZN(n552) );
  NAND2_X1 U371 ( .A1(n548), .A2(n526), .ZN(n618) );
  XNOR2_X1 U372 ( .A(n360), .B(n344), .ZN(n474) );
  XNOR2_X1 U373 ( .A(n425), .B(G140), .ZN(n700) );
  INV_X2 U374 ( .A(G953), .ZN(n702) );
  XNOR2_X2 U375 ( .A(n699), .B(n404), .ZN(n364) );
  XNOR2_X2 U376 ( .A(n402), .B(n401), .ZN(n699) );
  OR2_X1 U377 ( .A1(n681), .A2(G902), .ZN(n413) );
  AND2_X1 U378 ( .A1(n474), .A2(n650), .ZN(n430) );
  XNOR2_X1 U379 ( .A(n351), .B(n350), .ZN(n349) );
  INV_X1 U380 ( .A(KEYINPUT81), .ZN(n350) );
  NAND2_X1 U381 ( .A1(n618), .A2(KEYINPUT47), .ZN(n351) );
  XNOR2_X1 U382 ( .A(n355), .B(n482), .ZN(n354) );
  NAND2_X1 U383 ( .A1(n358), .A2(n356), .ZN(n355) );
  AND2_X1 U384 ( .A1(n711), .A2(n357), .ZN(n356) );
  AND2_X1 U385 ( .A1(n531), .A2(n646), .ZN(n431) );
  OR2_X1 U386 ( .A1(n584), .A2(G902), .ZN(n360) );
  XNOR2_X1 U387 ( .A(n424), .B(KEYINPUT10), .ZN(n425) );
  AND2_X1 U388 ( .A1(n524), .A2(n523), .ZN(n548) );
  NAND2_X1 U389 ( .A1(n354), .A2(n366), .ZN(n365) );
  AND2_X1 U390 ( .A1(n501), .A2(n502), .ZN(n366) );
  NOR2_X1 U391 ( .A1(n649), .A2(n518), .ZN(n530) );
  XNOR2_X1 U392 ( .A(n364), .B(n341), .ZN(n589) );
  XNOR2_X1 U393 ( .A(n362), .B(n361), .ZN(n457) );
  INV_X1 U394 ( .A(KEYINPUT8), .ZN(n361) );
  NAND2_X1 U395 ( .A1(n702), .A2(G234), .ZN(n362) );
  XNOR2_X1 U396 ( .A(n377), .B(G146), .ZN(n424) );
  XNOR2_X1 U397 ( .A(n432), .B(KEYINPUT107), .ZN(n433) );
  XNOR2_X1 U398 ( .A(n376), .B(n375), .ZN(n694) );
  XNOR2_X1 U399 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U400 ( .A(n427), .B(n342), .ZN(n584) );
  OR2_X1 U401 ( .A1(n558), .A2(n595), .ZN(n359) );
  XNOR2_X1 U402 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n480) );
  NOR2_X1 U403 ( .A1(n531), .A2(n484), .ZN(n340) );
  XOR2_X1 U404 ( .A(n407), .B(n406), .Z(n341) );
  XOR2_X1 U405 ( .A(n419), .B(n418), .Z(n342) );
  XOR2_X1 U406 ( .A(KEYINPUT23), .B(KEYINPUT70), .Z(n343) );
  XOR2_X1 U407 ( .A(n429), .B(KEYINPUT25), .Z(n344) );
  AND2_X1 U408 ( .A1(n628), .A2(n541), .ZN(n345) );
  NAND2_X1 U409 ( .A1(n665), .A2(KEYINPUT47), .ZN(n346) );
  XNOR2_X1 U410 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n347) );
  NAND2_X1 U411 ( .A1(n530), .A2(n519), .ZN(n522) );
  XNOR2_X2 U412 ( .A(n475), .B(KEYINPUT106), .ZN(n519) );
  XNOR2_X2 U413 ( .A(n348), .B(G472), .ZN(n475) );
  OR2_X2 U414 ( .A1(n589), .A2(G902), .ZN(n348) );
  NAND2_X1 U415 ( .A1(n349), .A2(n346), .ZN(n527) );
  NAND2_X1 U416 ( .A1(n555), .A2(n352), .ZN(n557) );
  XNOR2_X1 U417 ( .A(n529), .B(KEYINPUT80), .ZN(n353) );
  INV_X1 U418 ( .A(n616), .ZN(n357) );
  INV_X1 U419 ( .A(n714), .ZN(n358) );
  INV_X1 U420 ( .A(n552), .ZN(n602) );
  XNOR2_X1 U421 ( .A(n545), .B(KEYINPUT39), .ZN(n558) );
  XNOR2_X1 U422 ( .A(n364), .B(n412), .ZN(n681) );
  INV_X1 U423 ( .A(n567), .ZN(n691) );
  XNOR2_X2 U424 ( .A(n365), .B(n347), .ZN(n567) );
  XNOR2_X2 U425 ( .A(n450), .B(KEYINPUT13), .ZN(n487) );
  XNOR2_X2 U426 ( .A(n494), .B(n408), .ZN(n531) );
  XNOR2_X2 U427 ( .A(n460), .B(KEYINPUT4), .ZN(n402) );
  XNOR2_X1 U428 ( .A(n426), .B(n700), .ZN(n427) );
  XOR2_X1 U429 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n367) );
  XOR2_X1 U430 ( .A(G104), .B(G107), .Z(n368) );
  INV_X1 U431 ( .A(G125), .ZN(n377) );
  INV_X1 U432 ( .A(KEYINPUT30), .ZN(n503) );
  INV_X1 U433 ( .A(KEYINPUT85), .ZN(n535) );
  INV_X1 U434 ( .A(n568), .ZN(n569) );
  XNOR2_X1 U435 ( .A(n535), .B(KEYINPUT36), .ZN(n536) );
  XNOR2_X1 U436 ( .A(n537), .B(n536), .ZN(n538) );
  INV_X1 U437 ( .A(KEYINPUT63), .ZN(n593) );
  AND2_X1 U438 ( .A1(n575), .A2(n574), .ZN(G63) );
  XNOR2_X1 U439 ( .A(G110), .B(KEYINPUT76), .ZN(n369) );
  XNOR2_X1 U440 ( .A(n368), .B(n369), .ZN(n411) );
  INV_X1 U441 ( .A(KEYINPUT3), .ZN(n370) );
  XNOR2_X1 U442 ( .A(n370), .B(G119), .ZN(n372) );
  XNOR2_X1 U443 ( .A(G116), .B(G113), .ZN(n371) );
  XNOR2_X1 U444 ( .A(n372), .B(n371), .ZN(n407) );
  XNOR2_X1 U445 ( .A(n411), .B(n407), .ZN(n376) );
  XOR2_X1 U446 ( .A(KEYINPUT73), .B(G122), .Z(n374) );
  INV_X1 U447 ( .A(KEYINPUT16), .ZN(n373) );
  NAND2_X1 U448 ( .A1(G224), .A2(n702), .ZN(n379) );
  XNOR2_X2 U449 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n378) );
  XNOR2_X1 U450 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U451 ( .A(KEYINPUT67), .B(G101), .ZN(n403) );
  XNOR2_X1 U452 ( .A(n380), .B(n403), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n424), .B(n381), .ZN(n382) );
  XNOR2_X1 U454 ( .A(n382), .B(n402), .ZN(n383) );
  XNOR2_X1 U455 ( .A(n694), .B(n383), .ZN(n605) );
  XNOR2_X1 U456 ( .A(KEYINPUT87), .B(KEYINPUT15), .ZN(n384) );
  INV_X1 U457 ( .A(G902), .ZN(n463) );
  XNOR2_X1 U458 ( .A(n384), .B(n463), .ZN(n568) );
  NAND2_X1 U459 ( .A1(n605), .A2(n568), .ZN(n387) );
  INV_X1 U460 ( .A(G237), .ZN(n385) );
  NAND2_X1 U461 ( .A1(n463), .A2(n385), .ZN(n388) );
  AND2_X1 U462 ( .A1(n388), .A2(G210), .ZN(n386) );
  XNOR2_X2 U463 ( .A(n387), .B(n386), .ZN(n564) );
  NAND2_X1 U464 ( .A1(n388), .A2(G214), .ZN(n660) );
  NAND2_X1 U465 ( .A1(n564), .A2(n660), .ZN(n534) );
  XNOR2_X1 U466 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n389) );
  XNOR2_X1 U467 ( .A(n534), .B(n389), .ZN(n525) );
  NAND2_X1 U468 ( .A1(G237), .A2(G234), .ZN(n390) );
  XNOR2_X1 U469 ( .A(n390), .B(KEYINPUT88), .ZN(n391) );
  XNOR2_X1 U470 ( .A(KEYINPUT14), .B(n391), .ZN(n393) );
  NAND2_X1 U471 ( .A1(n393), .A2(G952), .ZN(n392) );
  XOR2_X1 U472 ( .A(KEYINPUT89), .B(n392), .Z(n673) );
  NOR2_X1 U473 ( .A1(n673), .A2(G953), .ZN(n505) );
  NOR2_X1 U474 ( .A1(G898), .A2(n702), .ZN(n696) );
  NAND2_X1 U475 ( .A1(n393), .A2(G902), .ZN(n394) );
  XOR2_X1 U476 ( .A(KEYINPUT90), .B(n394), .Z(n506) );
  NAND2_X1 U477 ( .A1(n696), .A2(n506), .ZN(n395) );
  XNOR2_X1 U478 ( .A(KEYINPUT91), .B(n395), .ZN(n396) );
  NOR2_X1 U479 ( .A1(n505), .A2(n396), .ZN(n397) );
  NOR2_X1 U480 ( .A1(n525), .A2(n397), .ZN(n398) );
  XNOR2_X1 U481 ( .A(KEYINPUT0), .B(n398), .ZN(n495) );
  INV_X1 U482 ( .A(n495), .ZN(n471) );
  XNOR2_X1 U483 ( .A(G137), .B(G134), .ZN(n400) );
  XNOR2_X1 U484 ( .A(G131), .B(KEYINPUT69), .ZN(n399) );
  XNOR2_X1 U485 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U486 ( .A(n403), .B(G146), .ZN(n404) );
  NOR2_X1 U487 ( .A1(G953), .A2(G237), .ZN(n436) );
  NAND2_X1 U488 ( .A1(n436), .A2(G210), .ZN(n405) );
  XNOR2_X1 U489 ( .A(n405), .B(KEYINPUT5), .ZN(n406) );
  BUF_X2 U490 ( .A(n475), .Z(n494) );
  INV_X1 U491 ( .A(KEYINPUT6), .ZN(n408) );
  NAND2_X1 U492 ( .A1(G227), .A2(n702), .ZN(n409) );
  XNOR2_X1 U493 ( .A(G140), .B(n409), .ZN(n410) );
  XNOR2_X1 U494 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X2 U495 ( .A(n524), .B(KEYINPUT1), .ZN(n646) );
  XOR2_X1 U496 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n415) );
  NAND2_X1 U497 ( .A1(G234), .A2(n568), .ZN(n414) );
  XNOR2_X1 U498 ( .A(n415), .B(n414), .ZN(n428) );
  NAND2_X1 U499 ( .A1(G221), .A2(n428), .ZN(n417) );
  INV_X1 U500 ( .A(KEYINPUT21), .ZN(n416) );
  XNOR2_X1 U501 ( .A(n417), .B(n416), .ZN(n650) );
  XOR2_X1 U502 ( .A(G137), .B(G119), .Z(n419) );
  XNOR2_X1 U503 ( .A(G128), .B(G110), .ZN(n418) );
  XNOR2_X1 U504 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n420) );
  XNOR2_X1 U505 ( .A(n343), .B(n420), .ZN(n421) );
  XNOR2_X1 U506 ( .A(n421), .B(n367), .ZN(n423) );
  NAND2_X1 U507 ( .A1(G221), .A2(n457), .ZN(n422) );
  XNOR2_X1 U508 ( .A(n423), .B(n422), .ZN(n426) );
  NAND2_X1 U509 ( .A1(n428), .A2(G217), .ZN(n429) );
  XNOR2_X2 U510 ( .A(n430), .B(KEYINPUT68), .ZN(n645) );
  AND2_X1 U511 ( .A1(n431), .A2(n645), .ZN(n434) );
  INV_X1 U512 ( .A(KEYINPUT33), .ZN(n432) );
  XNOR2_X1 U513 ( .A(n434), .B(n433), .ZN(n675) );
  NOR2_X1 U514 ( .A1(n471), .A2(n675), .ZN(n435) );
  XNOR2_X1 U515 ( .A(n435), .B(KEYINPUT34), .ZN(n466) );
  XOR2_X1 U516 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n438) );
  NAND2_X1 U517 ( .A1(n436), .A2(G214), .ZN(n437) );
  XNOR2_X1 U518 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U519 ( .A(KEYINPUT99), .B(KEYINPUT101), .Z(n440) );
  XNOR2_X1 U520 ( .A(G113), .B(KEYINPUT11), .ZN(n439) );
  XNOR2_X1 U521 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U522 ( .A(n442), .B(n441), .Z(n447) );
  XOR2_X1 U523 ( .A(G131), .B(G122), .Z(n444) );
  XNOR2_X1 U524 ( .A(G143), .B(G104), .ZN(n443) );
  XNOR2_X1 U525 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U526 ( .A(n700), .B(n445), .ZN(n446) );
  XNOR2_X1 U527 ( .A(n447), .B(n446), .ZN(n576) );
  NOR2_X1 U528 ( .A1(G902), .A2(n576), .ZN(n448) );
  XNOR2_X1 U529 ( .A(G475), .B(n448), .ZN(n449) );
  INV_X1 U530 ( .A(n449), .ZN(n450) );
  XOR2_X1 U531 ( .A(G134), .B(G122), .Z(n452) );
  XNOR2_X1 U532 ( .A(G107), .B(G116), .ZN(n451) );
  XNOR2_X1 U533 ( .A(n452), .B(n451), .ZN(n456) );
  XOR2_X1 U534 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n454) );
  XNOR2_X1 U535 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n453) );
  XNOR2_X1 U536 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U537 ( .A(n456), .B(n455), .Z(n459) );
  NAND2_X1 U538 ( .A1(G217), .A2(n457), .ZN(n458) );
  XNOR2_X1 U539 ( .A(n459), .B(n458), .ZN(n462) );
  INV_X1 U540 ( .A(n460), .ZN(n461) );
  XNOR2_X1 U541 ( .A(n462), .B(n461), .ZN(n571) );
  NAND2_X1 U542 ( .A1(n571), .A2(n463), .ZN(n465) );
  XOR2_X1 U543 ( .A(KEYINPUT104), .B(G478), .Z(n464) );
  XNOR2_X1 U544 ( .A(n465), .B(n464), .ZN(n485) );
  NOR2_X1 U545 ( .A1(n487), .A2(n485), .ZN(n513) );
  NAND2_X1 U546 ( .A1(n466), .A2(n513), .ZN(n467) );
  INV_X1 U547 ( .A(n650), .ZN(n468) );
  NAND2_X1 U548 ( .A1(n485), .A2(n487), .ZN(n663) );
  NOR2_X1 U549 ( .A1(n468), .A2(n663), .ZN(n469) );
  XNOR2_X1 U550 ( .A(n469), .B(KEYINPUT105), .ZN(n470) );
  NOR2_X2 U551 ( .A1(n471), .A2(n470), .ZN(n473) );
  XOR2_X1 U552 ( .A(KEYINPUT72), .B(KEYINPUT22), .Z(n472) );
  XNOR2_X1 U553 ( .A(n473), .B(n472), .ZN(n477) );
  NOR2_X1 U554 ( .A1(n477), .A2(n646), .ZN(n483) );
  BUF_X1 U555 ( .A(n474), .Z(n649) );
  NOR2_X1 U556 ( .A1(n649), .A2(n519), .ZN(n476) );
  AND2_X1 U557 ( .A1(n483), .A2(n476), .ZN(n616) );
  NOR2_X1 U558 ( .A1(n649), .A2(n477), .ZN(n479) );
  INV_X1 U559 ( .A(n646), .ZN(n488) );
  NOR2_X1 U560 ( .A1(n488), .A2(n531), .ZN(n478) );
  NAND2_X1 U561 ( .A1(n479), .A2(n478), .ZN(n481) );
  NOR2_X1 U562 ( .A1(KEYINPUT44), .A2(KEYINPUT71), .ZN(n482) );
  NAND2_X1 U563 ( .A1(KEYINPUT44), .A2(KEYINPUT71), .ZN(n502) );
  NAND2_X1 U564 ( .A1(n483), .A2(n649), .ZN(n484) );
  INV_X1 U565 ( .A(n485), .ZN(n486) );
  NOR2_X1 U566 ( .A1(n487), .A2(n486), .ZN(n622) );
  AND2_X1 U567 ( .A1(n487), .A2(n486), .ZN(n624) );
  NOR2_X1 U568 ( .A1(n622), .A2(n624), .ZN(n665) );
  NAND2_X1 U569 ( .A1(n645), .A2(n494), .ZN(n489) );
  NOR2_X1 U570 ( .A1(n489), .A2(n488), .ZN(n656) );
  NAND2_X1 U571 ( .A1(n656), .A2(n495), .ZN(n490) );
  XNOR2_X1 U572 ( .A(n490), .B(KEYINPUT31), .ZN(n491) );
  XNOR2_X1 U573 ( .A(KEYINPUT98), .B(n491), .ZN(n625) );
  NAND2_X1 U574 ( .A1(n645), .A2(n524), .ZN(n493) );
  INV_X1 U575 ( .A(KEYINPUT96), .ZN(n492) );
  XNOR2_X2 U576 ( .A(n493), .B(n492), .ZN(n511) );
  INV_X1 U577 ( .A(n511), .ZN(n497) );
  INV_X1 U578 ( .A(n494), .ZN(n652) );
  NAND2_X1 U579 ( .A1(n495), .A2(n652), .ZN(n496) );
  NOR2_X1 U580 ( .A1(n497), .A2(n496), .ZN(n498) );
  XOR2_X1 U581 ( .A(KEYINPUT97), .B(n498), .Z(n611) );
  NOR2_X1 U582 ( .A1(n625), .A2(n611), .ZN(n499) );
  NOR2_X1 U583 ( .A1(n665), .A2(n499), .ZN(n500) );
  NOR2_X1 U584 ( .A1(n340), .A2(n500), .ZN(n501) );
  NAND2_X1 U585 ( .A1(n519), .A2(n660), .ZN(n504) );
  XNOR2_X1 U586 ( .A(n504), .B(n503), .ZN(n510) );
  INV_X1 U587 ( .A(n505), .ZN(n509) );
  NAND2_X1 U588 ( .A1(G953), .A2(n506), .ZN(n507) );
  OR2_X1 U589 ( .A1(n507), .A2(G900), .ZN(n508) );
  NAND2_X1 U590 ( .A1(n509), .A2(n508), .ZN(n517) );
  AND2_X1 U591 ( .A1(n510), .A2(n517), .ZN(n512) );
  NAND2_X1 U592 ( .A1(n512), .A2(n511), .ZN(n544) );
  INV_X1 U593 ( .A(n544), .ZN(n515) );
  AND2_X1 U594 ( .A1(n513), .A2(n564), .ZN(n514) );
  NAND2_X1 U595 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U596 ( .A(n516), .B(KEYINPUT109), .ZN(n598) );
  XNOR2_X1 U597 ( .A(n598), .B(KEYINPUT82), .ZN(n528) );
  NAND2_X1 U598 ( .A1(n517), .A2(n650), .ZN(n518) );
  INV_X1 U599 ( .A(KEYINPUT110), .ZN(n520) );
  XNOR2_X1 U600 ( .A(n520), .B(KEYINPUT28), .ZN(n521) );
  XNOR2_X1 U601 ( .A(n522), .B(n521), .ZN(n523) );
  INV_X1 U602 ( .A(n525), .ZN(n526) );
  NOR2_X1 U603 ( .A1(n528), .A2(n527), .ZN(n529) );
  AND2_X1 U604 ( .A1(n530), .A2(n622), .ZN(n532) );
  NAND2_X1 U605 ( .A1(n532), .A2(n531), .ZN(n559) );
  XNOR2_X1 U606 ( .A(n559), .B(KEYINPUT112), .ZN(n533) );
  NOR2_X1 U607 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U608 ( .A1(n538), .A2(n646), .ZN(n628) );
  OR2_X1 U609 ( .A1(n665), .A2(KEYINPUT47), .ZN(n539) );
  OR2_X1 U610 ( .A1(n618), .A2(n539), .ZN(n540) );
  XNOR2_X1 U611 ( .A(n540), .B(KEYINPUT74), .ZN(n541) );
  XNOR2_X1 U612 ( .A(KEYINPUT75), .B(KEYINPUT38), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n564), .B(n542), .ZN(n661) );
  INV_X1 U614 ( .A(n661), .ZN(n543) );
  NOR2_X1 U615 ( .A1(n544), .A2(n543), .ZN(n545) );
  INV_X1 U616 ( .A(n622), .ZN(n595) );
  NAND2_X1 U617 ( .A1(n661), .A2(n660), .ZN(n664) );
  NOR2_X1 U618 ( .A1(n664), .A2(n663), .ZN(n546) );
  XNOR2_X1 U619 ( .A(KEYINPUT41), .B(n546), .ZN(n674) );
  INV_X1 U620 ( .A(n674), .ZN(n547) );
  NAND2_X1 U621 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U622 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n549) );
  XNOR2_X1 U623 ( .A(n550), .B(n549), .ZN(n713) );
  INV_X1 U624 ( .A(n713), .ZN(n551) );
  NAND2_X1 U625 ( .A1(n552), .A2(n551), .ZN(n554) );
  INV_X1 U626 ( .A(KEYINPUT46), .ZN(n553) );
  XNOR2_X1 U627 ( .A(n554), .B(n553), .ZN(n555) );
  INV_X1 U628 ( .A(KEYINPUT48), .ZN(n556) );
  XNOR2_X1 U629 ( .A(n557), .B(n556), .ZN(n566) );
  INV_X1 U630 ( .A(n624), .ZN(n617) );
  OR2_X1 U631 ( .A1(n558), .A2(n617), .ZN(n600) );
  XOR2_X1 U632 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n562) );
  NOR2_X1 U633 ( .A1(n646), .A2(n559), .ZN(n560) );
  NAND2_X1 U634 ( .A1(n660), .A2(n560), .ZN(n561) );
  XNOR2_X1 U635 ( .A(n562), .B(n561), .ZN(n563) );
  OR2_X1 U636 ( .A1(n564), .A2(n563), .ZN(n631) );
  AND2_X1 U637 ( .A1(n600), .A2(n631), .ZN(n565) );
  AND2_X2 U638 ( .A1(n566), .A2(n565), .ZN(n701) );
  NAND2_X2 U639 ( .A1(n567), .A2(n701), .ZN(n634) );
  XNOR2_X2 U640 ( .A(n634), .B(KEYINPUT2), .ZN(n570) );
  AND2_X4 U641 ( .A1(n570), .A2(n569), .ZN(n603) );
  NAND2_X1 U642 ( .A1(n603), .A2(G478), .ZN(n572) );
  XNOR2_X1 U643 ( .A(n572), .B(n571), .ZN(n575) );
  INV_X1 U644 ( .A(G952), .ZN(n573) );
  AND2_X1 U645 ( .A1(n573), .A2(G953), .ZN(n687) );
  INV_X1 U646 ( .A(n687), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n603), .A2(G475), .ZN(n580) );
  XOR2_X1 U648 ( .A(KEYINPUT59), .B(KEYINPUT121), .Z(n578) );
  XNOR2_X1 U649 ( .A(n576), .B(KEYINPUT65), .ZN(n577) );
  XNOR2_X1 U650 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U651 ( .A(n580), .B(n579), .ZN(n581) );
  NOR2_X2 U652 ( .A1(n581), .A2(n687), .ZN(n583) );
  XNOR2_X1 U653 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n583), .B(n582), .ZN(G60) );
  NAND2_X1 U655 ( .A1(n603), .A2(G217), .ZN(n585) );
  XNOR2_X1 U656 ( .A(n585), .B(n584), .ZN(n586) );
  NOR2_X2 U657 ( .A1(n586), .A2(n687), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT122), .ZN(G66) );
  NAND2_X1 U659 ( .A1(n603), .A2(G472), .ZN(n591) );
  XNOR2_X1 U660 ( .A(KEYINPUT86), .B(KEYINPUT62), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n591), .B(n590), .ZN(n592) );
  NOR2_X2 U663 ( .A1(n592), .A2(n687), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n594), .B(n593), .ZN(G57) );
  XOR2_X1 U665 ( .A(G146), .B(KEYINPUT115), .Z(n597) );
  NOR2_X1 U666 ( .A1(n618), .A2(n595), .ZN(n596) );
  XOR2_X1 U667 ( .A(n597), .B(n596), .Z(G48) );
  XOR2_X1 U668 ( .A(G143), .B(n598), .Z(G45) );
  XOR2_X1 U669 ( .A(G134), .B(KEYINPUT117), .Z(n599) );
  XNOR2_X1 U670 ( .A(n600), .B(n599), .ZN(G36) );
  XNOR2_X1 U671 ( .A(G131), .B(KEYINPUT127), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n602), .B(n601), .ZN(G33) );
  NAND2_X1 U673 ( .A1(n603), .A2(G210), .ZN(n607) );
  XNOR2_X1 U674 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n605), .B(n604), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n607), .B(n606), .ZN(n608) );
  NOR2_X2 U677 ( .A1(n608), .A2(n687), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n609), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U679 ( .A(G101), .B(n340), .Z(G3) );
  NAND2_X1 U680 ( .A1(n611), .A2(n622), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n610), .B(G104), .ZN(G6) );
  XOR2_X1 U682 ( .A(KEYINPUT113), .B(KEYINPUT26), .Z(n613) );
  NAND2_X1 U683 ( .A1(n611), .A2(n624), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n613), .B(n612), .ZN(n615) );
  XOR2_X1 U685 ( .A(G107), .B(KEYINPUT27), .Z(n614) );
  XNOR2_X1 U686 ( .A(n615), .B(n614), .ZN(G9) );
  XOR2_X1 U687 ( .A(G110), .B(n616), .Z(G12) );
  XOR2_X1 U688 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n620) );
  NOR2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U690 ( .A(n620), .B(n619), .Z(n621) );
  XNOR2_X1 U691 ( .A(G128), .B(n621), .ZN(G30) );
  NAND2_X1 U692 ( .A1(n625), .A2(n622), .ZN(n623) );
  XNOR2_X1 U693 ( .A(n623), .B(G113), .ZN(G15) );
  NAND2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U695 ( .A(n626), .B(KEYINPUT116), .ZN(n627) );
  XNOR2_X1 U696 ( .A(G116), .B(n627), .ZN(G18) );
  INV_X1 U697 ( .A(n628), .ZN(n629) );
  XNOR2_X1 U698 ( .A(G125), .B(n629), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n630), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U700 ( .A(n631), .ZN(n632) );
  XOR2_X1 U701 ( .A(G140), .B(n632), .Z(n633) );
  XNOR2_X1 U702 ( .A(KEYINPUT118), .B(n633), .ZN(G42) );
  BUF_X1 U703 ( .A(n634), .Z(n635) );
  INV_X1 U704 ( .A(n635), .ZN(n636) );
  NAND2_X1 U705 ( .A1(n636), .A2(KEYINPUT2), .ZN(n638) );
  XNOR2_X1 U706 ( .A(KEYINPUT79), .B(KEYINPUT2), .ZN(n639) );
  NAND2_X1 U707 ( .A1(n691), .A2(n639), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n643) );
  INV_X1 U709 ( .A(n701), .ZN(n640) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(KEYINPUT83), .ZN(n642) );
  NOR2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U713 ( .A1(G953), .A2(n644), .ZN(n679) );
  NOR2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U715 ( .A(KEYINPUT119), .B(n647), .Z(n648) );
  XNOR2_X1 U716 ( .A(n648), .B(KEYINPUT50), .ZN(n655) );
  NOR2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U718 ( .A(n651), .B(KEYINPUT49), .ZN(n653) );
  NAND2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n657) );
  NOR2_X1 U721 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U722 ( .A(KEYINPUT51), .B(n658), .Z(n659) );
  NOR2_X1 U723 ( .A1(n674), .A2(n659), .ZN(n670) );
  NOR2_X1 U724 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U725 ( .A1(n663), .A2(n662), .ZN(n667) );
  NOR2_X1 U726 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U727 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U728 ( .A1(n668), .A2(n675), .ZN(n669) );
  NOR2_X1 U729 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U730 ( .A(n671), .B(KEYINPUT52), .ZN(n672) );
  NOR2_X1 U731 ( .A1(n673), .A2(n672), .ZN(n677) );
  NOR2_X1 U732 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U733 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U734 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U735 ( .A(KEYINPUT53), .B(n680), .Z(G75) );
  NAND2_X1 U736 ( .A1(n603), .A2(G469), .ZN(n685) );
  XOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n683) );
  XNOR2_X1 U738 ( .A(n681), .B(KEYINPUT120), .ZN(n682) );
  XNOR2_X1 U739 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U740 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U741 ( .A1(n687), .A2(n686), .ZN(G54) );
  NAND2_X1 U742 ( .A1(G953), .A2(G224), .ZN(n688) );
  XNOR2_X1 U743 ( .A(KEYINPUT61), .B(n688), .ZN(n689) );
  NAND2_X1 U744 ( .A1(n689), .A2(G898), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n690), .B(KEYINPUT123), .ZN(n693) );
  NOR2_X1 U746 ( .A1(G953), .A2(n691), .ZN(n692) );
  NOR2_X1 U747 ( .A1(n693), .A2(n692), .ZN(n698) );
  XOR2_X1 U748 ( .A(n694), .B(G101), .Z(n695) );
  NOR2_X1 U749 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U750 ( .A(n698), .B(n697), .Z(G69) );
  XNOR2_X1 U751 ( .A(n699), .B(n700), .ZN(n704) );
  XNOR2_X1 U752 ( .A(n701), .B(n704), .ZN(n703) );
  NAND2_X1 U753 ( .A1(n703), .A2(n702), .ZN(n709) );
  XOR2_X1 U754 ( .A(G227), .B(n704), .Z(n705) );
  NAND2_X1 U755 ( .A1(n705), .A2(G900), .ZN(n706) );
  XNOR2_X1 U756 ( .A(KEYINPUT124), .B(n706), .ZN(n707) );
  NAND2_X1 U757 ( .A1(n707), .A2(G953), .ZN(n708) );
  NAND2_X1 U758 ( .A1(n709), .A2(n708), .ZN(G72) );
  XOR2_X1 U759 ( .A(G119), .B(KEYINPUT125), .Z(n710) );
  XNOR2_X1 U760 ( .A(n711), .B(n710), .ZN(G21) );
  XOR2_X1 U761 ( .A(G137), .B(KEYINPUT126), .Z(n712) );
  XNOR2_X1 U762 ( .A(n713), .B(n712), .ZN(G39) );
  XOR2_X1 U763 ( .A(G122), .B(n714), .Z(G24) );
endmodule

