//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT81), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n191), .B(new_n193), .Z(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(G107), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n197), .A2(new_n200), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n196), .A2(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n199), .A2(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(G101), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n211), .B1(G143), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n210), .B1(new_n213), .B2(KEYINPUT82), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n209), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n215), .A2(new_n221), .A3(new_n211), .A4(G128), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n208), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT10), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(KEYINPUT83), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT83), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n215), .A2(new_n221), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n213), .A2(KEYINPUT82), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT82), .B(KEYINPUT1), .C1(new_n220), .C2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G128), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n228), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n207), .B1(new_n232), .B2(new_n222), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n227), .B1(new_n233), .B2(KEYINPUT10), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n228), .B1(new_n213), .B2(new_n210), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n222), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n208), .A2(KEYINPUT10), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  OR2_X1    g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n228), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n209), .A2(KEYINPUT0), .A3(G128), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n197), .A2(new_n200), .A3(new_n202), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G101), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(new_n248), .A3(G101), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n238), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G134), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT11), .B1(new_n252), .B2(G137), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G134), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT64), .B1(new_n255), .B2(G134), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n252), .A3(G137), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(G131), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n253), .A2(new_n256), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n263), .A2(new_n264), .A3(new_n258), .A4(new_n260), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(KEYINPUT65), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n267), .B(G131), .C1(new_n257), .C2(new_n261), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n235), .A2(new_n251), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n269), .B1(new_n235), .B2(new_n251), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n195), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n235), .A2(new_n251), .A3(new_n269), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n208), .A2(new_n237), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(new_n233), .ZN(new_n275));
  OR3_X1    g089(.A1(new_n275), .A2(KEYINPUT12), .A3(new_n269), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT12), .B1(new_n275), .B2(new_n269), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n273), .A2(new_n276), .A3(new_n194), .A4(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n272), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n189), .B1(new_n279), .B2(new_n187), .ZN(new_n280));
  OR3_X1    g094(.A1(new_n270), .A2(new_n271), .A3(new_n195), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n273), .A2(new_n277), .A3(new_n276), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n195), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n280), .B1(new_n187), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G221), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT9), .B(G234), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n288), .B2(new_n188), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G214), .B1(G237), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G210), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G125), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n236), .A2(new_n297), .A3(new_n222), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n241), .B2(new_n242), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n192), .A2(G224), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT88), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT89), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n301), .B(new_n304), .Z(new_n305));
  INV_X1    g119(.A(G116), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT68), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G116), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n309), .A3(G119), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT67), .ZN(new_n311));
  INV_X1    g125(.A(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(KEYINPUT67), .A2(G119), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(G116), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G113), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT2), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G113), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n310), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT69), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n310), .A2(new_n315), .A3(new_n323), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n310), .A2(new_n315), .ZN(new_n326));
  INV_X1    g140(.A(new_n320), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT84), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n250), .A3(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n322), .A2(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n247), .A2(new_n249), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT84), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n315), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(new_n316), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n310), .A2(new_n315), .A3(new_n335), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n325), .A3(new_n208), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n331), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G122), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(KEYINPUT86), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n345), .B1(new_n341), .B2(new_n343), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n332), .A2(new_n333), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n338), .A2(new_n337), .B1(new_n322), .B2(new_n324), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n350), .A2(new_n330), .B1(new_n208), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n352), .A2(new_n353), .A3(new_n342), .A4(new_n334), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n331), .A2(new_n334), .A3(new_n342), .A4(new_n340), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT87), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n356), .A3(KEYINPUT6), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n305), .B1(new_n349), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n355), .B(new_n353), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n303), .A2(KEYINPUT7), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n299), .B2(new_n300), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n243), .A2(G125), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(KEYINPUT7), .A3(new_n298), .A4(new_n303), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n339), .A2(new_n325), .A3(new_n207), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n342), .B(KEYINPUT8), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n337), .B1(new_n368), .B2(new_n326), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n207), .B1(new_n369), .B2(new_n325), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n364), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT90), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n364), .B(KEYINPUT90), .C1(new_n367), .C2(new_n370), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n188), .B1(new_n359), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n296), .B1(new_n358), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n305), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n354), .A2(KEYINPUT6), .A3(new_n356), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n341), .A2(new_n343), .ZN(new_n380));
  INV_X1    g194(.A(new_n345), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n346), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n378), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n373), .A2(new_n374), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n354), .A2(new_n356), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n387), .A3(new_n295), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n294), .B1(new_n377), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(G237), .A2(G953), .ZN(new_n390));
  AOI21_X1  g204(.A(G143), .B1(new_n390), .B2(G214), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(G143), .A3(G214), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT18), .A3(G131), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n212), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT18), .A2(G131), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n392), .A2(new_n393), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n401));
  OR3_X1    g215(.A1(new_n297), .A2(KEYINPUT16), .A3(G140), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(G146), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT75), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n401), .A2(KEYINPUT75), .A3(G146), .A4(new_n402), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n401), .A2(new_n402), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n405), .B(new_n406), .C1(G146), .C2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n394), .A2(KEYINPUT17), .A3(G131), .ZN(new_n409));
  INV_X1    g223(.A(new_n393), .ZN(new_n410));
  OAI21_X1  g224(.A(G131), .B1(new_n410), .B2(new_n391), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n392), .A2(new_n264), .A3(new_n393), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n409), .B1(new_n413), .B2(KEYINPUT17), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n400), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(new_n196), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n417), .B(new_n400), .C1(new_n408), .C2(new_n414), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n188), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G475), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n396), .B(KEYINPUT19), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n212), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT78), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n403), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n401), .A2(KEYINPUT78), .A3(G146), .A4(new_n402), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n425), .A2(new_n413), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n400), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n418), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n420), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n432), .A2(KEYINPUT91), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n431), .B2(new_n420), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT91), .B1(new_n437), .B2(new_n433), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n423), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n220), .A2(G128), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n210), .A2(G143), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(G134), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT92), .B1(new_n306), .B2(G122), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT92), .ZN(new_n446));
  INV_X1    g260(.A(G122), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G116), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n307), .A2(new_n309), .A3(G122), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n199), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n450), .A2(KEYINPUT14), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n449), .B1(new_n450), .B2(KEYINPUT14), .ZN(new_n454));
  OAI21_X1  g268(.A(G107), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT93), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n449), .A2(new_n450), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G107), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n451), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT13), .B1(new_n210), .B2(G143), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n443), .B1(new_n252), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT13), .A4(G134), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n457), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n449), .A2(new_n450), .A3(new_n199), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n199), .B1(new_n449), .B2(new_n450), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n464), .B(new_n457), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n456), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT74), .B(G217), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n288), .A2(new_n192), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT94), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n472), .A2(new_n473), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n470), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT93), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n478), .A2(new_n468), .B1(new_n455), .B2(new_n452), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n473), .A3(new_n472), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n480), .A3(new_n188), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n481), .B(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G952), .ZN(new_n485));
  AOI211_X1 g299(.A(G953), .B(new_n485), .C1(G234), .C2(G237), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n188), .B(new_n192), .C1(G234), .C2(G237), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT21), .B(G898), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n440), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n292), .A2(new_n389), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n266), .A2(new_n244), .A3(new_n268), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n255), .A2(G134), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n252), .A2(G137), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n264), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n496), .A2(KEYINPUT66), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(KEYINPUT66), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n237), .A2(new_n497), .A3(new_n265), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n332), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(new_n499), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT30), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n493), .A2(new_n503), .A3(new_n499), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT70), .B1(new_n505), .B2(new_n329), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n493), .A2(new_n503), .A3(new_n499), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n503), .B1(new_n493), .B2(new_n499), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT70), .B(new_n329), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n500), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT72), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n390), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT27), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(G101), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n512), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n500), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n329), .B1(new_n507), .B2(new_n508), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT70), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n519), .B1(new_n522), .B2(new_n509), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT72), .B1(new_n523), .B2(new_n516), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n332), .B1(new_n493), .B2(new_n499), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT28), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n519), .A2(KEYINPUT28), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT29), .B1(new_n529), .B2(new_n516), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n518), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n528), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n526), .A2(KEYINPUT73), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n516), .A2(KEYINPUT29), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n537), .A2(new_n188), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n500), .A2(new_n516), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n506), .B2(new_n510), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n522), .A2(new_n509), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT31), .A3(new_n543), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n517), .B1(new_n527), .B2(new_n528), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n541), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g365(.A1(G472), .A2(new_n539), .B1(new_n551), .B2(KEYINPUT32), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n553));
  INV_X1    g367(.A(new_n550), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n546), .B2(new_n548), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n555), .B2(new_n541), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT32), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT31), .B1(new_n547), .B2(new_n543), .ZN(new_n558));
  AOI211_X1 g372(.A(new_n545), .B(new_n542), .C1(new_n522), .C2(new_n509), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n550), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(KEYINPUT71), .A3(new_n540), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n552), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n427), .A2(new_n428), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n396), .A2(new_n212), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n313), .A2(new_n314), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(G128), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT76), .B(G110), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n312), .A2(new_n210), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n568), .B2(new_n210), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n569), .B(new_n570), .C1(new_n572), .C2(new_n567), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT24), .B(G110), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT77), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n573), .A2(new_n576), .A3(KEYINPUT77), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n566), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n569), .B1(new_n572), .B2(new_n567), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n583), .A2(G110), .B1(new_n575), .B2(new_n572), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n408), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT22), .B(G137), .ZN(new_n586));
  INV_X1    g400(.A(G234), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n286), .A2(new_n587), .A3(G953), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n586), .B(new_n588), .Z(new_n589));
  NAND3_X1  g403(.A1(new_n582), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n589), .ZN(new_n591));
  INV_X1    g405(.A(new_n585), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n581), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n471), .B1(new_n587), .B2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n188), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT79), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT25), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n590), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n598), .A2(new_n599), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n595), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n597), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n492), .B1(new_n563), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n605), .ZN(new_n607));
  AOI211_X1 g421(.A(KEYINPUT80), .B(new_n607), .C1(new_n552), .C2(new_n562), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n491), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT95), .B(G101), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G3));
  AND2_X1   g425(.A1(new_n556), .A2(new_n561), .ZN(new_n612));
  INV_X1    g426(.A(G472), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n560), .B2(new_n188), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n291), .A2(new_n607), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n358), .A2(new_n376), .A3(new_n296), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n295), .B1(new_n384), .B2(new_n387), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n293), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n472), .A2(KEYINPUT96), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n479), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n470), .A2(KEYINPUT96), .A3(new_n472), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT97), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n476), .A2(new_n480), .A3(new_n622), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT97), .B1(new_n624), .B2(new_n625), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n482), .A2(G902), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT98), .B1(new_n481), .B2(new_n482), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n481), .A2(KEYINPUT98), .A3(new_n482), .ZN(new_n634));
  OAI22_X1  g448(.A1(new_n630), .A2(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n489), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n440), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT99), .B1(new_n621), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n634), .A2(new_n633), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n629), .A2(new_n628), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n632), .B1(new_n640), .B2(new_n626), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n440), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n389), .A2(new_n644), .A3(new_n645), .A4(new_n636), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n638), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n618), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  INV_X1    g464(.A(new_n484), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n437), .A2(new_n433), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n437), .A2(new_n433), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n423), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n621), .A2(new_n489), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n618), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NAND2_X1  g473(.A1(new_n612), .A2(new_n615), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n582), .A2(new_n585), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n591), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n596), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n603), .A2(new_n604), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n292), .A2(new_n389), .A3(new_n490), .A4(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT37), .B(G110), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT100), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n668), .B(new_n670), .ZN(G12));
  NAND3_X1  g485(.A1(new_n666), .A2(new_n285), .A3(new_n290), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT101), .B(G900), .Z(new_n674));
  AOI21_X1  g488(.A(new_n486), .B1(new_n487), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n423), .B(new_n676), .C1(new_n653), .C2(new_n652), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n651), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n389), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n563), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT102), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n672), .B1(new_n552), .B2(new_n562), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n679), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  NAND2_X1  g500(.A1(new_n511), .A2(new_n516), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n519), .A2(new_n525), .ZN(new_n688));
  AOI21_X1  g502(.A(G902), .B1(new_n688), .B2(new_n517), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n613), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n551), .B2(KEYINPUT32), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n562), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT103), .Z(new_n693));
  AND2_X1   g507(.A1(new_n440), .A2(new_n484), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n665), .A2(new_n694), .A3(new_n293), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n675), .B(KEYINPUT39), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n292), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n695), .B1(new_n697), .B2(KEYINPUT40), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n377), .A2(new_n388), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT38), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n693), .A2(new_n698), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT104), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  OAI211_X1 g518(.A(new_n440), .B(new_n676), .C1(new_n639), .C2(new_n641), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT105), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n635), .A2(new_n707), .A3(new_n440), .A4(new_n676), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n621), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n682), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  XNOR2_X1  g526(.A(new_n279), .B(new_n187), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n289), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n605), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n647), .A2(new_n563), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  AND3_X1   g533(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n539), .A2(G472), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n551), .A2(KEYINPUT32), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n656), .B(new_n716), .C1(new_n720), .C2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n715), .B1(new_n552), .B2(new_n562), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(KEYINPUT106), .A3(new_n656), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  INV_X1    g544(.A(new_n714), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n621), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n666), .A2(new_n490), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n563), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  NOR2_X1   g549(.A1(new_n731), .A2(new_n489), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n517), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n541), .B1(new_n549), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n614), .A2(new_n607), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n389), .A2(KEYINPUT107), .A3(new_n694), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT107), .B1(new_n389), .B2(new_n694), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n736), .B(new_n740), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  OR3_X1    g559(.A1(new_n614), .A2(new_n739), .A3(new_n665), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n709), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n732), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NAND2_X1  g563(.A1(new_n283), .A2(KEYINPUT108), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n282), .A2(new_n751), .A3(new_n195), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n750), .A2(G469), .A3(new_n281), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n289), .B1(new_n280), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n293), .A3(new_n377), .A4(new_n388), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n709), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n557), .B1(new_n555), .B2(new_n541), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n721), .A2(new_n722), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n605), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT42), .ZN(new_n760));
  INV_X1    g574(.A(new_n755), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n709), .A2(KEYINPUT42), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n563), .A2(new_n761), .A3(new_n762), .A4(new_n605), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n264), .ZN(G33));
  NAND4_X1  g579(.A1(new_n563), .A2(new_n761), .A3(new_n605), .A4(new_n678), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  NOR2_X1   g581(.A1(new_n642), .A2(new_n440), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT43), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n660), .A2(new_n666), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(KEYINPUT109), .Z(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n187), .B1(new_n284), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n750), .A2(new_n281), .A3(new_n752), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n776), .B2(new_n774), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n777), .B1(new_n187), .B2(new_n188), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(KEYINPUT46), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n279), .A2(new_n187), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n779), .B2(KEYINPUT46), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n290), .B(new_n696), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n377), .A2(new_n388), .A3(new_n293), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(new_n770), .B2(new_n771), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n773), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  OAI21_X1  g602(.A(new_n290), .B1(new_n780), .B2(new_n782), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT47), .ZN(new_n790));
  OR4_X1    g604(.A1(new_n563), .A2(new_n605), .A3(new_n709), .A4(new_n785), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NOR2_X1   g607(.A1(new_n693), .A2(new_n607), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n713), .A2(KEYINPUT49), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n713), .A2(KEYINPUT49), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n289), .A2(new_n294), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n768), .A3(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n700), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n727), .A2(KEYINPUT106), .A3(new_n656), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT106), .B1(new_n727), .B2(new_n656), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n717), .A2(new_n734), .A3(new_n744), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT110), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n644), .B1(new_n643), .B2(new_n484), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n807), .A2(new_n621), .A3(new_n489), .ZN(new_n808));
  OAI22_X1  g622(.A1(new_n808), .A2(new_n617), .B1(new_n660), .B2(new_n667), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n606), .A2(new_n608), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n491), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n760), .A2(new_n763), .A3(new_n766), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n747), .A2(new_n761), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n677), .A2(new_n484), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n377), .A2(new_n814), .A3(new_n388), .A4(new_n293), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT111), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n682), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n717), .A2(new_n734), .A3(new_n744), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n729), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n806), .A2(new_n811), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n754), .A2(new_n665), .A3(new_n676), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n562), .B2(new_n691), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n699), .A2(new_n293), .A3(new_n694), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT107), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n741), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n710), .A2(new_n682), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n682), .A2(new_n683), .A3(new_n679), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n683), .B1(new_n682), .B2(new_n679), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n830), .B(new_n748), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n685), .A2(new_n835), .A3(new_n748), .A4(new_n830), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n801), .B1(new_n823), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n747), .A2(new_n761), .B1(new_n682), .B2(new_n816), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(new_n760), .A3(new_n763), .A4(new_n766), .ZN(new_n840));
  INV_X1    g654(.A(new_n609), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n840), .A2(new_n841), .A3(new_n809), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n804), .A2(new_n801), .A3(new_n805), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n836), .A3(new_n843), .A4(new_n834), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(KEYINPUT54), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n820), .A2(new_n729), .A3(new_n821), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n821), .B1(new_n820), .B2(new_n729), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n836), .A3(new_n834), .A4(new_n842), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(new_n801), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n846), .B1(new_n851), .B2(KEYINPUT54), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n790), .B1(new_n290), .B2(new_n713), .ZN(new_n853));
  INV_X1    g667(.A(new_n785), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n769), .A2(new_n486), .A3(new_n740), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n731), .A2(new_n785), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n486), .B1(new_n857), .B2(KEYINPUT113), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(KEYINPUT113), .B2(new_n857), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n794), .A2(new_n859), .A3(new_n643), .A4(new_n642), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n769), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(new_n746), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT112), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n294), .B1(new_n863), .B2(KEYINPUT50), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n700), .A2(new_n731), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n855), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(KEYINPUT50), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n856), .A2(new_n860), .A3(new_n862), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n607), .B1(new_n552), .B2(new_n757), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n859), .A2(new_n873), .A3(new_n769), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT48), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n794), .A2(new_n859), .A3(new_n644), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n485), .B(G953), .C1(new_n855), .C2(new_n732), .ZN(new_n879));
  XOR2_X1   g693(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n852), .A2(new_n871), .A3(new_n872), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n800), .B1(new_n883), .B2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n192), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n805), .B1(new_n726), .B2(new_n728), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n811), .A2(new_n888), .A3(new_n819), .A4(KEYINPUT53), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n837), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n850), .B2(new_n801), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n188), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT56), .B1(new_n892), .B2(G210), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n379), .A2(new_n383), .A3(new_n378), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n358), .ZN(new_n895));
  XOR2_X1   g709(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n896));
  XNOR2_X1  g710(.A(new_n895), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n887), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n893), .B2(new_n897), .ZN(G51));
  NAND2_X1  g713(.A1(new_n272), .A2(new_n278), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n891), .B(KEYINPUT54), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n189), .B(KEYINPUT57), .Z(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n777), .B(KEYINPUT116), .Z(new_n904));
  NAND2_X1  g718(.A1(new_n892), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n886), .B1(new_n903), .B2(new_n905), .ZN(G54));
  AND3_X1   g720(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n887), .B1(new_n907), .B2(new_n432), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n432), .B2(new_n907), .ZN(G60));
  XOR2_X1   g723(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n910));
  NOR2_X1   g724(.A1(new_n482), .A2(new_n188), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n630), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n887), .B1(new_n901), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n915), .A2(KEYINPUT118), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n630), .B1(new_n852), .B2(new_n912), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(KEYINPUT118), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G63));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n921));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT60), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n891), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n923), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n845), .A2(KEYINPUT119), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n924), .A2(new_n594), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n887), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT119), .B1(new_n845), .B2(new_n925), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n921), .B(new_n923), .C1(new_n838), .C2(new_n844), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n663), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT120), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n933), .B(new_n663), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n928), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n920), .B1(new_n935), .B2(KEYINPUT61), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n929), .A2(new_n930), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n886), .B1(new_n937), .B2(new_n594), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n924), .A2(new_n926), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n933), .B1(new_n939), .B2(new_n663), .ZN(new_n940));
  INV_X1    g754(.A(new_n934), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(KEYINPUT121), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n936), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(KEYINPUT61), .B(new_n938), .C1(new_n940), .C2(new_n941), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n932), .A2(new_n934), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(KEYINPUT122), .A3(KEYINPUT61), .A4(new_n938), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n945), .A2(new_n951), .ZN(G66));
  INV_X1    g766(.A(new_n488), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n192), .B1(new_n953), .B2(G224), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n849), .A2(new_n811), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT123), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n954), .B1(new_n957), .B2(new_n192), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n349), .B(new_n357), .C1(G898), .C2(new_n192), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n958), .B(new_n959), .Z(G69));
  XOR2_X1   g774(.A(new_n505), .B(new_n424), .Z(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(G900), .B2(G953), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n685), .A2(new_n711), .A3(new_n748), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n784), .A2(new_n829), .A3(new_n873), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n787), .A2(new_n792), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n812), .B(KEYINPUT126), .Z(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT127), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n962), .B1(new_n968), .B2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n787), .A2(new_n792), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n697), .A2(new_n807), .A3(new_n785), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n810), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n703), .A2(new_n963), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n972), .A2(new_n974), .A3(new_n978), .A4(new_n975), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n961), .B(KEYINPUT124), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n969), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n968), .B2(new_n957), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n517), .A3(new_n523), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n518), .A2(new_n524), .A3(new_n544), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n989), .A2(new_n986), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n886), .B1(new_n851), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n977), .A2(new_n956), .A3(new_n979), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n687), .B1(new_n993), .B2(new_n986), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n992), .A2(new_n994), .ZN(G57));
endmodule


