//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n201), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n209), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n224));
  OR2_X1    g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(new_n203), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(new_n223), .B2(new_n224), .ZN(new_n233));
  AND4_X1   g0033(.A1(new_n219), .A2(new_n220), .A3(new_n225), .A4(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G68), .Z(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  AOI21_X1  g0049(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G1698), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n257), .A2(G222), .B1(G77), .B2(new_n256), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT66), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT66), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n262), .A3(G1698), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n260), .A2(G223), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n251), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT65), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G33), .A3(G41), .ZN(new_n274));
  INV_X1    g0074(.A(new_n226), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n267), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n270), .B1(new_n277), .B2(new_n211), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n265), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G200), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT68), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n226), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(new_n266), .B2(G20), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n284), .B1(new_n287), .B2(G50), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n227), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(G20), .B2(new_n204), .ZN(new_n295));
  INV_X1    g0095(.A(new_n286), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n288), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XOR2_X1   g0097(.A(new_n297), .B(KEYINPUT9), .Z(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(G190), .B2(new_n279), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n282), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n282), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n283), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n203), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT12), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n292), .A2(G50), .ZN(new_n308));
  INV_X1    g0108(.A(G77), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n308), .B1(new_n227), .B2(G68), .C1(new_n309), .C2(new_n290), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(KEYINPUT11), .A3(new_n286), .ZN(new_n311));
  INV_X1    g0111(.A(new_n287), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n307), .B(new_n311), .C1(new_n203), .C2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT11), .B1(new_n310), .B2(new_n286), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n253), .A2(new_n255), .A3(G232), .A4(G1698), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n253), .A2(new_n255), .A3(G226), .A4(new_n259), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n250), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n276), .A2(KEYINPUT69), .A3(new_n267), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G238), .ZN(new_n323));
  INV_X1    g0123(.A(G41), .ZN(new_n324));
  INV_X1    g0124(.A(G45), .ZN(new_n325));
  AOI21_X1  g0125(.A(G1), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n226), .B1(KEYINPUT65), .B2(new_n271), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(new_n274), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(KEYINPUT69), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n270), .B(new_n321), .C1(new_n323), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT13), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n269), .B1(new_n320), .B2(new_n250), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n332), .B(new_n333), .C1(new_n329), .C2(new_n323), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n331), .A2(G179), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n331), .B2(new_n334), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT14), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI211_X1 g0139(.A(KEYINPUT14), .B(new_n336), .C1(new_n331), .C2(new_n334), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n316), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n331), .A2(new_n334), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G200), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n315), .C1(new_n344), .C2(new_n342), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n280), .A2(new_n336), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n279), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n347), .A2(new_n297), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G232), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n256), .A2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n259), .B1(G107), .B2(new_n256), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n260), .A2(G238), .A3(new_n263), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n251), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G244), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n270), .B1(new_n277), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(G200), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n289), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n292), .B1(G20), .B2(G77), .ZN(new_n361));
  XOR2_X1   g0161(.A(KEYINPUT15), .B(G87), .Z(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(new_n227), .A3(G33), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n296), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n305), .A2(new_n309), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n312), .B2(new_n309), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n368), .A2(KEYINPUT67), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n356), .A2(new_n358), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G190), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n368), .B2(KEYINPUT67), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n348), .ZN(new_n374));
  INV_X1    g0174(.A(new_n367), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n336), .B1(new_n356), .B2(new_n358), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n304), .A2(new_n346), .A3(new_n351), .A4(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT71), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n269), .B1(new_n328), .B2(G232), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n253), .A2(new_n255), .A3(G226), .A4(G1698), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n253), .A2(new_n255), .A3(G223), .A4(new_n259), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G87), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n250), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n382), .A2(new_n387), .A3(new_n344), .ZN(new_n388));
  AOI21_X1  g0188(.A(G200), .B1(new_n382), .B2(new_n387), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n381), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G200), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n386), .A2(new_n250), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n270), .B1(new_n277), .B2(new_n352), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n382), .A2(new_n387), .A3(new_n344), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(KEYINPUT71), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT7), .B1(new_n256), .B2(new_n227), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n398), .B(G20), .C1(new_n253), .C2(new_n255), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n230), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G20), .ZN(new_n403));
  INV_X1    g0203(.A(G159), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT70), .B1(new_n293), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT70), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n292), .A2(new_n406), .A3(G159), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n400), .A2(new_n409), .A3(KEYINPUT16), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n398), .B1(new_n261), .B2(G20), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n254), .A2(G33), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT7), .B(new_n227), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n203), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n411), .B1(new_n416), .B2(new_n408), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n410), .A2(new_n417), .A3(new_n286), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n360), .A2(new_n305), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n312), .B2(new_n360), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n390), .A2(new_n396), .A3(new_n418), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT72), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n400), .A2(new_n409), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n296), .B1(new_n424), .B2(new_n411), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n420), .B1(new_n425), .B2(new_n410), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT72), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n426), .A2(new_n427), .A3(new_n396), .A4(new_n390), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(KEYINPUT17), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n418), .A2(new_n421), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n382), .A2(new_n387), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G169), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n348), .B2(new_n431), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n430), .A2(KEYINPUT18), .A3(new_n433), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n422), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n429), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n380), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n253), .A2(new_n255), .A3(G250), .A4(new_n259), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n253), .A2(new_n255), .A3(G257), .A4(G1698), .ZN(new_n444));
  INV_X1    g0244(.A(G294), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n443), .B(new_n444), .C1(new_n252), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n250), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n325), .A2(G1), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G41), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n451), .A4(G274), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n276), .A2(new_n453), .A3(G264), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n447), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT81), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT81), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n447), .A2(new_n457), .A3(new_n452), .A4(new_n454), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n344), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n391), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT74), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n266), .A2(G33), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n296), .A2(new_n462), .A3(new_n283), .A4(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n283), .A2(new_n463), .A3(new_n226), .A4(new_n285), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT74), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G107), .ZN(new_n468));
  INV_X1    g0268(.A(G107), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n305), .B(new_n469), .C1(KEYINPUT80), .C2(KEYINPUT25), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT80), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT25), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(new_n283), .C2(G107), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n470), .B(new_n473), .C1(new_n471), .C2(new_n472), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT23), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n227), .B2(G107), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n469), .A2(KEYINPUT23), .A3(G20), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n227), .A2(G33), .A3(G116), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n261), .A2(new_n227), .A3(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n261), .A2(new_n484), .A3(new_n227), .A4(G87), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n481), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n286), .B1(new_n486), .B2(KEYINPUT24), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(KEYINPUT24), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n475), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n461), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n489), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n468), .B(new_n474), .C1(new_n492), .C2(new_n487), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n336), .B1(new_n456), .B2(new_n458), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n455), .A2(new_n348), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT82), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT82), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n491), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n276), .A2(new_n453), .A3(G270), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n502), .A2(new_n452), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n253), .A2(new_n255), .A3(G257), .A4(new_n259), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n253), .A2(new_n255), .A3(G264), .A4(G1698), .ZN(new_n505));
  INV_X1    g0305(.A(G303), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(new_n261), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n250), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G116), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n465), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n305), .A2(new_n510), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n285), .A2(new_n226), .B1(G20), .B2(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G283), .ZN(new_n514));
  INV_X1    g0314(.A(G97), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n514), .B(new_n227), .C1(G33), .C2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT20), .B1(new_n513), .B2(new_n516), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n511), .B(new_n512), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n509), .A2(new_n520), .A3(G169), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n520), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n503), .A2(new_n508), .A3(G190), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n502), .A2(new_n452), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n250), .B2(new_n507), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n524), .B(new_n525), .C1(new_n527), .C2(new_n391), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n509), .A2(new_n520), .A3(KEYINPUT21), .A4(G169), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(G179), .A3(new_n520), .ZN(new_n530));
  AND4_X1   g0330(.A1(new_n523), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n253), .A2(new_n255), .A3(G238), .A4(new_n259), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n253), .A2(new_n255), .A3(G244), .A4(G1698), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n532), .B(new_n533), .C1(new_n252), .C2(new_n510), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n250), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n325), .A2(new_n268), .A3(G1), .ZN(new_n536));
  OAI21_X1  g0336(.A(G250), .B1(new_n325), .B2(G1), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n276), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n348), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT78), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n535), .A2(new_n539), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n336), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n467), .A2(new_n362), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n206), .A2(new_n212), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT79), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT79), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n206), .A2(new_n547), .A3(new_n212), .ZN(new_n548));
  NAND3_X1  g0348(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n546), .A2(new_n548), .B1(new_n227), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n253), .A2(new_n255), .A3(new_n227), .A4(G68), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n290), .A2(new_n515), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(KEYINPUT19), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n286), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n362), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n305), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n544), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT78), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n535), .A2(new_n558), .A3(new_n348), .A4(new_n539), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n541), .A2(new_n543), .A3(new_n557), .A4(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n554), .A2(new_n556), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n542), .A2(G200), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n535), .A2(G190), .A3(new_n539), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n467), .A2(G87), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n292), .A2(G77), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT6), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT73), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n571), .B2(new_n206), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n207), .A2(KEYINPUT73), .A3(new_n568), .A4(new_n570), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n568), .C2(G97), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n567), .B1(new_n574), .B2(new_n227), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n469), .B1(new_n412), .B2(new_n415), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n286), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n467), .A2(G97), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n283), .A2(G97), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT75), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n515), .B1(new_n464), .B2(new_n466), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT75), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n582), .A2(new_n583), .A3(new_n579), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n577), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n253), .A2(new_n255), .A3(G244), .A4(new_n259), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT76), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT4), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n253), .A2(new_n255), .A3(G250), .A4(G1698), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n589), .A2(new_n514), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n250), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n276), .A2(new_n453), .A3(G257), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT77), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n276), .A2(new_n453), .A3(KEYINPUT77), .A4(G257), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n452), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n594), .A2(new_n600), .A3(new_n348), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n592), .A2(new_n514), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(KEYINPUT4), .B2(new_n588), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n251), .B1(new_n603), .B2(new_n591), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n336), .B1(new_n604), .B2(new_n599), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n585), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(G200), .B1(new_n604), .B2(new_n599), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n594), .A2(new_n600), .A3(G190), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n578), .A2(KEYINPUT75), .A3(new_n580), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n583), .B1(new_n582), .B2(new_n579), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n607), .A2(new_n608), .A3(new_n577), .A4(new_n611), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n531), .A2(new_n566), .A3(new_n606), .A4(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n442), .A2(new_n501), .A3(new_n613), .ZN(G372));
  INV_X1    g0414(.A(KEYINPUT84), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT83), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n539), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n537), .B1(new_n327), .B2(new_n274), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT83), .B1(new_n618), .B2(new_n536), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(G169), .B1(new_n620), .B2(new_n535), .ZN(new_n621));
  INV_X1    g0421(.A(new_n540), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n615), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n617), .A2(new_n619), .B1(new_n250), .B2(new_n534), .ZN(new_n624));
  OAI211_X1 g0424(.A(KEYINPUT84), .B(new_n540), .C1(new_n624), .C2(G169), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n623), .A2(new_n625), .B1(new_n561), .B2(new_n544), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n563), .A2(new_n564), .A3(new_n556), .A4(new_n554), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT85), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n624), .B2(new_n391), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n539), .A2(new_n616), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n618), .A2(KEYINPUT83), .A3(new_n536), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n535), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(KEYINPUT85), .A3(G200), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n627), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n606), .A2(new_n612), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n493), .B1(new_n459), .B2(new_n460), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n496), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n626), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n627), .A2(new_n633), .A3(new_n629), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n626), .A2(new_n641), .A3(new_n606), .ZN(new_n642));
  INV_X1    g0442(.A(new_n606), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n566), .ZN(new_n644));
  XOR2_X1   g0444(.A(KEYINPUT86), .B(KEYINPUT26), .Z(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n642), .A2(KEYINPUT26), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n442), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n341), .A2(new_n377), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n429), .A2(new_n440), .A3(new_n345), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n438), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n350), .B1(new_n652), .B2(new_n304), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(G13), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G20), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n266), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n501), .B1(new_n490), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n496), .B2(new_n663), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n520), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n531), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n638), .B2(new_n666), .ZN(new_n668));
  XOR2_X1   g0468(.A(KEYINPUT87), .B(G330), .Z(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n638), .A2(new_n662), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n501), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n496), .A2(new_n662), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(G399));
  NAND3_X1  g0477(.A1(new_n546), .A2(new_n510), .A3(new_n548), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n221), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n679), .A2(new_n682), .A3(G1), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n231), .B2(new_n682), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n662), .B1(new_n640), .B2(new_n647), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n642), .A2(KEYINPUT26), .B1(new_n644), .B2(new_n646), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n632), .A2(new_n336), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT84), .B1(new_n688), .B2(new_n540), .ZN(new_n689));
  INV_X1    g0489(.A(new_n625), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n557), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n491), .A2(new_n606), .A3(new_n612), .A4(new_n634), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n496), .A2(new_n638), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n663), .B1(new_n687), .B2(new_n694), .ZN(new_n695));
  MUX2_X1   g0495(.A(new_n686), .B(new_n695), .S(KEYINPUT29), .Z(new_n696));
  NAND4_X1  g0496(.A1(new_n613), .A2(new_n498), .A3(new_n500), .A4(new_n663), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT88), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n509), .B2(new_n348), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n527), .A2(KEYINPUT88), .A3(G179), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n542), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n447), .A2(new_n454), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n594), .A2(new_n704), .A3(new_n705), .A4(new_n600), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n699), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n447), .A2(new_n535), .A3(new_n454), .A4(new_n539), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n708), .A2(new_n604), .A3(new_n599), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(KEYINPUT30), .A3(new_n701), .A4(new_n702), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n594), .A2(new_n600), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT89), .B1(new_n711), .B2(new_n455), .ZN(new_n712));
  OAI211_X1 g0512(.A(KEYINPUT89), .B(new_n455), .C1(new_n604), .C2(new_n599), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n632), .A2(new_n348), .A3(new_n509), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n707), .B(new_n710), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n698), .B1(new_n717), .B2(new_n662), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n697), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n698), .A3(new_n662), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n720), .A2(new_n669), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n696), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n685), .B1(new_n723), .B2(G1), .ZN(G364));
  AOI21_X1  g0524(.A(new_n266), .B1(new_n656), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n681), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(G355), .A2(new_n221), .A3(new_n261), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n248), .A2(new_n325), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n680), .A2(new_n261), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G45), .B2(new_n231), .ZN(new_n732));
  OAI221_X1 g0532(.A(new_n729), .B1(G116), .B2(new_n221), .C1(new_n730), .C2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G13), .A2(G33), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n226), .B1(G20), .B2(new_n336), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT90), .Z(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n728), .B1(new_n733), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT91), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n227), .A2(new_n344), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n348), .A2(new_n391), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n348), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n745), .A2(new_n201), .B1(new_n747), .B2(new_n202), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n227), .A2(G190), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n746), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n748), .B1(G77), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT92), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n391), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n469), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n256), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n743), .A2(new_n754), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n212), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n744), .A2(new_n749), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n759), .B1(G68), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G179), .A2(G200), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n227), .B1(new_n763), .B2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G97), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n749), .A2(new_n763), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G159), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n766), .B1(new_n769), .B2(KEYINPUT32), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(KEYINPUT32), .B2(new_n769), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n753), .A2(new_n757), .A3(new_n762), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT93), .ZN(new_n773));
  INV_X1    g0573(.A(G326), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n745), .A2(new_n774), .B1(new_n758), .B2(new_n506), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n261), .B(new_n775), .C1(G329), .C2(new_n768), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  INV_X1    g0577(.A(new_n755), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n761), .A2(new_n777), .B1(new_n778), .B2(G283), .ZN(new_n779));
  INV_X1    g0579(.A(new_n747), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G322), .A2(new_n780), .B1(new_n751), .B2(G311), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n765), .A2(G294), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n776), .A2(new_n779), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(KEYINPUT94), .B1(new_n773), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n737), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n773), .A2(KEYINPUT94), .A3(new_n783), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n742), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n736), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n668), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n671), .A2(new_n727), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n669), .B2(new_n668), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n790), .A2(new_n792), .ZN(G396));
  NOR2_X1   g0593(.A1(new_n377), .A2(new_n662), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n369), .A2(new_n372), .B1(new_n367), .B2(new_n663), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(new_n795), .B2(new_n377), .ZN(new_n796));
  AOI21_X1  g0596(.A(KEYINPUT96), .B1(new_n686), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n686), .A2(new_n796), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n797), .B(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n722), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n728), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT97), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n801), .A2(new_n802), .B1(new_n800), .B2(new_n799), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G143), .A2(new_n780), .B1(new_n761), .B2(G150), .ZN(new_n806));
  INV_X1    g0606(.A(new_n745), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G137), .B1(new_n751), .B2(G159), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n261), .B1(new_n758), .B2(new_n201), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n755), .A2(new_n203), .B1(new_n767), .B2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n812), .B(new_n814), .C1(G58), .C2(new_n765), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n810), .A2(new_n811), .A3(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n761), .A2(KEYINPUT95), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n761), .A2(KEYINPUT95), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n212), .A2(new_n755), .B1(new_n750), .B2(new_n510), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n261), .B(new_n822), .C1(G294), .C2(new_n780), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n745), .A2(new_n506), .B1(new_n767), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n758), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(G107), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n821), .A2(new_n766), .A3(new_n823), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n816), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n737), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n737), .A2(new_n734), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n728), .B1(new_n309), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n830), .B(new_n832), .C1(new_n796), .C2(new_n735), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n805), .A2(new_n833), .ZN(G384));
  INV_X1    g0634(.A(KEYINPUT35), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n510), .B(new_n229), .C1(new_n574), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n835), .B2(new_n574), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT36), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n401), .A2(G77), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n231), .A2(new_n841), .B1(G50), .B2(new_n203), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(G1), .A3(new_n655), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n839), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT98), .Z(new_n845));
  NAND2_X1  g0645(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n717), .B2(new_n662), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n707), .A2(new_n710), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT89), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n604), .A2(new_n599), .ZN(new_n851));
  INV_X1    g0651(.A(new_n455), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n716), .B1(new_n853), .B2(new_n713), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n662), .B(new_n847), .C1(new_n849), .C2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n697), .B1(new_n848), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n796), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n316), .A2(new_n662), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n341), .A2(new_n345), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n316), .B(new_n662), .C1(new_n339), .C2(new_n340), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n860), .A2(KEYINPUT99), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT99), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT102), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n418), .A2(KEYINPUT100), .A3(new_n421), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT100), .B1(new_n418), .B2(new_n421), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n867), .A2(new_n868), .A3(new_n660), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n441), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n423), .A2(new_n428), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n431), .A2(new_n348), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G169), .B2(new_n431), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n873), .A2(new_n660), .B1(new_n418), .B2(new_n421), .ZN(new_n874));
  XNOR2_X1  g0674(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n867), .A2(new_n868), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n660), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n423), .A2(new_n428), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n870), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n870), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n866), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n870), .A2(new_n882), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n870), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(KEYINPUT102), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n865), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n426), .A2(new_n660), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n441), .A2(KEYINPUT104), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT104), .B1(new_n441), .B2(new_n893), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n422), .B(new_n434), .C1(new_n426), .C2(new_n660), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n875), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n877), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g0700(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n889), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n858), .A2(new_n864), .A3(new_n892), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n891), .A2(new_n892), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n442), .A2(new_n857), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n669), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n696), .A2(new_n442), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n653), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n341), .A2(new_n662), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n914), .B(new_n889), .C1(new_n900), .C2(new_n902), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT39), .B1(new_n883), .B2(new_n884), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n691), .A2(new_n643), .A3(new_n634), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT26), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n560), .A2(new_n565), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n606), .A2(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n918), .A2(new_n919), .B1(new_n921), .B2(new_n645), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n663), .B(new_n796), .C1(new_n922), .C2(new_n694), .ZN(new_n923));
  INV_X1    g0723(.A(new_n794), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n860), .A2(new_n861), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT99), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n860), .A2(KEYINPUT99), .A3(new_n861), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n923), .A2(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n885), .A2(new_n890), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n436), .A2(new_n437), .A3(new_n660), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n917), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n912), .A2(new_n934), .B1(new_n266), .B2(new_n656), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n912), .A2(new_n934), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n845), .B1(new_n935), .B2(new_n936), .ZN(G367));
  NAND2_X1  g0737(.A1(new_n561), .A2(new_n564), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n662), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n691), .A2(new_n634), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n691), .B2(new_n939), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT43), .B1(new_n941), .B2(KEYINPUT106), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(KEYINPUT106), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n643), .A2(new_n662), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n585), .A2(new_n662), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n606), .A2(new_n612), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n501), .A2(new_n673), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n606), .B1(new_n948), .B2(new_n496), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n950), .A2(KEYINPUT42), .B1(new_n663), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(KEYINPUT42), .B2(new_n950), .ZN(new_n953));
  MUX2_X1   g0753(.A(new_n943), .B(new_n945), .S(new_n953), .Z(new_n954));
  AOI21_X1  g0754(.A(new_n672), .B1(new_n948), .B2(new_n946), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n681), .B(KEYINPUT41), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n676), .A2(new_n949), .ZN(new_n960));
  XOR2_X1   g0760(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n676), .A2(new_n949), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n963));
  AOI22_X1  g0763(.A1(new_n960), .A2(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n676), .C2(new_n949), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n962), .A2(new_n963), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n672), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n964), .A2(new_n966), .A3(new_n672), .A4(new_n965), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n674), .B1(new_n665), .B2(new_n673), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT109), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n972), .A3(new_n671), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n670), .B(KEYINPUT109), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n973), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n969), .A2(new_n723), .A3(new_n970), .A4(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n959), .B1(new_n976), .B2(new_n723), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n956), .B(new_n957), .C1(new_n977), .C2(new_n726), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n740), .B1(new_n221), .B2(new_n555), .ZN(new_n979));
  INV_X1    g0779(.A(new_n731), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n241), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n727), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT110), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n758), .B2(new_n510), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n820), .A2(G294), .B1(KEYINPUT46), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(KEYINPUT46), .B2(new_n984), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n807), .A2(G311), .B1(new_n778), .B2(G97), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G283), .A2(new_n751), .B1(new_n768), .B2(G317), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n765), .A2(G107), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n261), .B1(new_n780), .B2(G303), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n807), .A2(G143), .B1(new_n778), .B2(G77), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n256), .B1(new_n826), .B2(G58), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n203), .C2(new_n764), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G150), .A2(new_n780), .B1(new_n751), .B2(G50), .ZN(new_n995));
  INV_X1    g0795(.A(G137), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(new_n996), .B2(new_n767), .C1(new_n819), .C2(new_n404), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n986), .A2(new_n991), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT47), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n785), .B1(new_n998), .B2(new_n999), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n982), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n941), .B2(new_n789), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n978), .A2(new_n1003), .ZN(G387));
  OR2_X1    g0804(.A1(new_n665), .A2(new_n789), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n678), .A2(new_n221), .A3(new_n261), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(G107), .B2(new_n221), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n980), .B1(new_n238), .B2(G45), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n679), .A2(KEYINPUT111), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n679), .A2(KEYINPUT111), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n289), .A2(G50), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g0812(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1007), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n727), .B1(new_n1015), .B2(new_n739), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n261), .B1(new_n768), .B2(G326), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n807), .A2(G322), .B1(new_n751), .B2(G303), .ZN(new_n1018));
  INV_X1    g0818(.A(G317), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n747), .C1(new_n819), .C2(new_n824), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT48), .Z(new_n1021));
  INV_X1    g0821(.A(G283), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n758), .A2(new_n445), .B1(new_n764), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1017), .B1(new_n510), .B2(new_n755), .C1(new_n1024), .C2(KEYINPUT49), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1024), .A2(KEYINPUT49), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n745), .A2(KEYINPUT112), .A3(new_n404), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT112), .B1(new_n745), .B2(new_n404), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n555), .C2(new_n764), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n758), .A2(new_n309), .B1(new_n767), .B2(new_n291), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n256), .B(new_n1030), .C1(G97), .C2(new_n778), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G50), .A2(new_n780), .B1(new_n751), .B2(G68), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n289), .C2(new_n760), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1025), .A2(new_n1026), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1016), .B1(new_n1034), .B2(new_n737), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n975), .A2(new_n726), .B1(new_n1005), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n975), .A2(new_n723), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n681), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n975), .A2(new_n723), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(G393));
  OAI21_X1  g0840(.A(new_n740), .B1(new_n515), .B2(new_n221), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n245), .A2(new_n980), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n727), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n820), .A2(G50), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n745), .A2(new_n291), .B1(new_n747), .B2(new_n404), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n758), .A2(new_n203), .B1(new_n750), .B2(new_n289), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G143), .B2(new_n768), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n764), .A2(new_n309), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n256), .B(new_n1049), .C1(G87), .C2(new_n778), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1044), .A2(new_n1046), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G283), .A2(new_n826), .B1(new_n768), .B2(G322), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT113), .Z(new_n1053));
  AOI211_X1 g0853(.A(new_n261), .B(new_n756), .C1(G294), .C2(new_n751), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n510), .C2(new_n764), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT52), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n745), .A2(new_n1019), .B1(new_n747), .B2(new_n824), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n820), .A2(G303), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1051), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1043), .B1(new_n1060), .B2(new_n737), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n949), .B2(new_n789), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n969), .A2(new_n970), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(new_n1037), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n976), .A2(new_n681), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1062), .B1(new_n725), .B2(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(G390));
  OAI22_X1  g0866(.A1(new_n918), .A2(new_n919), .B1(new_n921), .B2(new_n645), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n662), .B1(new_n640), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n795), .A2(new_n377), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n794), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n913), .B1(new_n1070), .B2(new_n864), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n441), .A2(new_n893), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT104), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n441), .A2(KEYINPUT104), .A3(new_n893), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n1075), .A3(new_n898), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n883), .B1(new_n1076), .B2(new_n901), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT114), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n913), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1069), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n924), .B1(new_n695), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n927), .A2(new_n928), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT114), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n903), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1078), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n722), .A2(new_n796), .A3(new_n1082), .ZN(new_n1087));
  OAI21_X1  g0887(.A(KEYINPUT115), .B1(new_n929), .B2(new_n1079), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT115), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n794), .B1(new_n686), .B2(new_n796), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1089), .B(new_n913), .C1(new_n1090), .C2(new_n864), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1088), .A2(new_n1091), .A3(new_n915), .A4(new_n916), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1086), .A2(new_n1087), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n442), .A2(G330), .A3(new_n857), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n910), .A2(new_n1094), .A3(new_n653), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1082), .A2(G330), .A3(new_n796), .A4(new_n857), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n719), .A2(new_n721), .A3(new_n796), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n864), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1090), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(G330), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n864), .B1(new_n858), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n1087), .A3(new_n1070), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1095), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT116), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n915), .A2(new_n916), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1107), .A2(new_n1108), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1093), .B1(new_n1105), .B2(new_n1106), .C1(new_n1109), .C2(new_n1096), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1093), .B1(new_n1109), .B2(new_n1096), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1105), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(KEYINPUT116), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1110), .A2(new_n1113), .A3(new_n681), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1111), .A2(new_n725), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1108), .A2(new_n734), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n831), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n727), .B1(new_n360), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n820), .A2(G137), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n745), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(G125), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n747), .A2(new_n813), .B1(new_n767), .B2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT54), .B(G143), .Z(new_n1124));
  AOI211_X1 g0924(.A(new_n1121), .B(new_n1123), .C1(new_n751), .C2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n758), .A2(new_n291), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n261), .B1(new_n755), .B2(new_n201), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G159), .B2(new_n765), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1119), .A2(new_n1125), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n819), .A2(new_n469), .B1(new_n515), .B2(new_n750), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT117), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n807), .A2(G283), .B1(new_n778), .B2(G68), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G116), .A2(new_n780), .B1(new_n768), .B2(G294), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n759), .A2(new_n1049), .A3(new_n261), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1131), .A2(KEYINPUT117), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1130), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1118), .B1(new_n1138), .B2(new_n737), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1116), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1115), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1114), .A2(new_n1141), .ZN(G378));
  INV_X1    g0942(.A(KEYINPUT57), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n891), .A2(new_n892), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n904), .A2(new_n903), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(G330), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n933), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n905), .B(G330), .C1(new_n917), .C2(new_n932), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n304), .A2(new_n351), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n660), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n297), .A2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1150), .B(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1153), .B(new_n1154), .Z(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1149), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1147), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1143), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1093), .B(new_n1105), .C1(new_n1109), .C2(new_n1096), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1095), .B(KEYINPUT122), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n682), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT121), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1147), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1155), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1157), .A2(KEYINPUT121), .A3(new_n1158), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1164), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1163), .B1(new_n1170), .B2(KEYINPUT57), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n725), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n727), .B1(G50), .B2(new_n1117), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n1120), .A2(new_n747), .B1(new_n760), .B2(new_n813), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n826), .A2(new_n1124), .B1(new_n751), .B2(G137), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n1122), .B2(new_n745), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1174), .B(new_n1176), .C1(G150), .C2(new_n765), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT59), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(G33), .A2(G41), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT118), .Z(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G159), .A2(new_n778), .B1(new_n768), .B2(G124), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1179), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G41), .B(new_n261), .C1(new_n768), .C2(G283), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n202), .B2(new_n755), .C1(new_n309), .C2(new_n758), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT119), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n745), .A2(new_n510), .B1(new_n747), .B2(new_n469), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n555), .A2(new_n750), .B1(new_n515), .B2(new_n760), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(G68), .C2(new_n765), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(KEYINPUT58), .A3(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1181), .B(new_n201), .C1(G41), .C2(new_n261), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1185), .A2(new_n1192), .A3(new_n1193), .A4(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1173), .B1(new_n1197), .B2(new_n737), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1156), .B2(new_n735), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT120), .Z(new_n1200));
  NOR2_X1   g1000(.A1(new_n1172), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1171), .A2(new_n1201), .ZN(G375));
  AND2_X1   g1002(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1095), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT123), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT123), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1203), .A2(new_n1206), .A3(new_n1095), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(new_n958), .A3(new_n1112), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT124), .Z(new_n1210));
  AOI21_X1  g1010(.A(new_n728), .B1(new_n203), .B2(new_n831), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G283), .A2(new_n780), .B1(new_n768), .B2(G303), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n515), .B2(new_n758), .C1(new_n819), .C2(new_n510), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n555), .A2(new_n764), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n256), .B1(new_n755), .B2(new_n309), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n745), .A2(new_n445), .B1(new_n750), .B2(new_n469), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n820), .A2(new_n1124), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n813), .B2(new_n745), .C1(new_n996), .C2(new_n747), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT125), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n261), .B1(new_n755), .B2(new_n202), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G50), .B2(new_n765), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G159), .A2(new_n826), .B1(new_n751), .B2(G150), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n1120), .C2(new_n767), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1219), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1224), .A2(new_n1220), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1217), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1211), .B1(new_n785), .B2(new_n1227), .C1(new_n1082), .C2(new_n735), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n1203), .B2(new_n725), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT126), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1229), .B(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1210), .A2(new_n1231), .ZN(G381));
  OR2_X1    g1032(.A1(G393), .A2(G396), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(G378), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1171), .A2(new_n1235), .A3(new_n1201), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1234), .A2(G381), .A3(new_n1236), .ZN(G407));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G343), .C2(new_n1236), .ZN(G409));
  INV_X1    g1038(.A(G390), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(G387), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G390), .A2(new_n1003), .A3(new_n978), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  XOR2_X1   g1042(.A(G393), .B(G396), .Z(new_n1243));
  XNOR2_X1  g1043(.A(new_n1242), .B(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT61), .ZN(new_n1246));
  INV_X1    g1046(.A(G384), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n681), .B1(new_n1204), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1112), .A2(KEYINPUT60), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1208), .B2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1229), .B(KEYINPUT126), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1247), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1205), .A2(new_n1207), .B1(new_n1112), .B2(KEYINPUT60), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1231), .B(G384), .C1(new_n1254), .C2(new_n1249), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n661), .A2(G213), .A3(G2897), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1253), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1235), .B1(new_n1171), .B2(new_n1201), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n661), .A2(G213), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n959), .B(new_n1164), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n726), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1114), .A2(new_n1141), .A3(new_n1199), .A4(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1261), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1259), .B1(new_n1260), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1260), .A2(new_n1267), .A3(new_n1265), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1246), .B(new_n1266), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1245), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1265), .B1(G378), .B2(G375), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1267), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT63), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1266), .A2(new_n1246), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G375), .A2(G378), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1265), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(KEYINPUT63), .A3(new_n1279), .A4(new_n1274), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1244), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT127), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1246), .B(new_n1266), .C1(new_n1268), .C2(KEYINPUT63), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1244), .A2(new_n1280), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT127), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1272), .B1(new_n1282), .B2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(new_n1278), .A2(new_n1236), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(new_n1274), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(new_n1244), .ZN(G402));
endmodule


