//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT66), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n215), .B1(new_n218), .B2(new_n220), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT68), .Z(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n239), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G68), .ZN(new_n249));
  INV_X1    g0049(.A(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n248), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT71), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT71), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n258), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n216), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT72), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT72), .A4(new_n216), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n262), .A2(KEYINPUT73), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT73), .B1(new_n262), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XOR2_X1   g0066(.A(KEYINPUT8), .B(G58), .Z(new_n267));
  NAND2_X1  g0067(.A1(new_n210), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n267), .A2(new_n269), .B1(G150), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(new_n204), .B2(new_n210), .ZN(new_n272));
  INV_X1    g0072(.A(G13), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n273), .A2(new_n210), .A3(G1), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n266), .A2(new_n272), .B1(new_n202), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT73), .ZN(new_n276));
  AND2_X1   g0076(.A1(G1), .A2(G13), .ZN(new_n277));
  AND3_X1   g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n258), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT72), .B1(new_n279), .B2(new_n257), .ZN(new_n280));
  INV_X1    g0080(.A(new_n263), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n262), .A2(KEYINPUT73), .A3(new_n263), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n274), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n210), .A2(G1), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(G50), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n275), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT9), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT9), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n275), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT69), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT69), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G1698), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G222), .ZN(new_n299));
  INV_X1    g0099(.A(G223), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n294), .B1(KEYINPUT70), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(KEYINPUT70), .B2(new_n300), .ZN(new_n302));
  OR2_X1    g0102(.A1(KEYINPUT3), .A2(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT3), .A2(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n299), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n306), .B(new_n307), .C1(G77), .C2(new_n305), .ZN(new_n308));
  INV_X1    g0108(.A(G274), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G41), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(new_n277), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G41), .ZN(new_n312));
  INV_X1    g0112(.A(G45), .ZN(new_n313));
  AOI21_X1  g0113(.A(G1), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n277), .A2(new_n310), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n316), .B1(G226), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n308), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G200), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(G190), .B2(new_n322), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n292), .A2(new_n293), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n293), .B1(new_n292), .B2(new_n325), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g0131(.A(new_n331), .B(KEYINPUT74), .Z(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n288), .C1(G169), .C2(new_n322), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n319), .A2(KEYINPUT77), .ZN(new_n336));
  INV_X1    g0136(.A(G238), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n319), .B2(KEYINPUT77), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n316), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  AND2_X1   g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NOR2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n295), .A2(new_n297), .A3(G226), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G232), .A2(G1698), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n307), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n339), .A2(new_n340), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT79), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n339), .A2(new_n349), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT13), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n339), .A2(KEYINPUT79), .A3(new_n340), .A4(new_n349), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n352), .A2(new_n354), .A3(G190), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n274), .A2(new_n250), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT12), .ZN(new_n358));
  INV_X1    g0158(.A(new_n274), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n280), .B2(new_n281), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n286), .A2(G68), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT80), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n269), .A2(G77), .B1(G20), .B2(new_n250), .ZN(new_n364));
  INV_X1    g0164(.A(new_n270), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n202), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n282), .A2(new_n283), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT11), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n356), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT78), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n350), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n339), .A2(KEYINPUT78), .A3(new_n340), .A4(new_n349), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n354), .A3(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n373), .A2(G200), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(G169), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT14), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n352), .A2(new_n354), .A3(G179), .A4(new_n355), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT14), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n373), .A2(new_n379), .A3(G169), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n363), .A2(new_n368), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n375), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G58), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n250), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n385), .B2(new_n201), .ZN(new_n386));
  INV_X1    g0186(.A(G159), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n365), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n303), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n304), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT81), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n305), .B2(G20), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT81), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n343), .A2(new_n393), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n388), .B1(new_n395), .B2(G68), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n280), .A2(new_n281), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n250), .B1(new_n392), .B2(new_n389), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(new_n388), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n267), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n359), .B1(new_n403), .B2(new_n285), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n284), .B2(new_n403), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n315), .B1(new_n319), .B2(new_n241), .ZN(new_n407));
  OAI211_X1 g0207(.A(G226), .B(G1698), .C1(new_n341), .C2(new_n342), .ZN(new_n408));
  INV_X1    g0208(.A(G33), .ZN(new_n409));
  INV_X1    g0209(.A(G87), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n295), .B(new_n297), .C1(new_n341), .C2(new_n342), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n408), .B1(new_n409), .B2(new_n410), .C1(new_n411), .C2(new_n300), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n407), .B1(new_n412), .B2(new_n307), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n413), .A2(G179), .ZN(new_n414));
  INV_X1    g0214(.A(G169), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n406), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT18), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n406), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G190), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n413), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G200), .B2(new_n413), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(new_n402), .A3(new_n405), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n424), .A2(new_n402), .A3(new_n405), .A4(KEYINPUT17), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n419), .A2(new_n421), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n316), .B1(G244), .B2(new_n320), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n294), .B1(new_n303), .B2(new_n304), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G238), .ZN(new_n432));
  INV_X1    g0232(.A(G107), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n305), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT75), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n411), .B2(new_n241), .ZN(new_n436));
  INV_X1    g0236(.A(new_n411), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(KEYINPUT75), .A3(G232), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n434), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n430), .B1(new_n439), .B2(new_n317), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n415), .ZN(new_n441));
  OR3_X1    g0241(.A1(new_n360), .A2(new_n205), .A3(new_n285), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT15), .B(G87), .ZN(new_n443));
  OR3_X1    g0243(.A1(new_n443), .A2(KEYINPUT76), .A3(new_n268), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n267), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT76), .B1(new_n443), .B2(new_n268), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(new_n398), .B1(new_n205), .B2(new_n274), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n441), .A2(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n440), .A2(G179), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n440), .A2(G200), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n453), .B(new_n454), .C1(new_n422), .C2(new_n440), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n429), .A2(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n335), .A2(new_n383), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n409), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n210), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT23), .B1(new_n433), .B2(G20), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n463), .A2(new_n210), .A3(G107), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n461), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT88), .B(KEYINPUT22), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n305), .A2(new_n466), .A3(new_n210), .A4(G87), .ZN(new_n467));
  INV_X1    g0267(.A(new_n466), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n210), .B(G87), .C1(new_n341), .C2(new_n342), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n465), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI211_X1 g0273(.A(KEYINPUT24), .B(new_n465), .C1(new_n467), .C2(new_n470), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n398), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n282), .A2(new_n283), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n409), .A2(G1), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n476), .A2(G107), .A3(new_n359), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n274), .A2(new_n433), .ZN(new_n480));
  XOR2_X1   g0280(.A(new_n480), .B(KEYINPUT25), .Z(new_n481));
  NAND3_X1  g0281(.A1(new_n475), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(G257), .B(G1698), .C1(new_n341), .C2(new_n342), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G294), .ZN(new_n484));
  INV_X1    g0284(.A(G250), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(new_n484), .C1(new_n411), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n307), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n313), .A2(G1), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n488), .A2(new_n489), .B1(new_n277), .B2(new_n310), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n209), .A2(G45), .ZN(new_n491));
  NOR2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n490), .A2(G264), .B1(new_n311), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(G179), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n415), .B2(new_n497), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n482), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT89), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n487), .A2(new_n496), .A3(new_n501), .A4(new_n422), .ZN(new_n502));
  AND2_X1   g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n489), .B1(new_n503), .B2(new_n492), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(G264), .A3(new_n317), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n311), .A2(new_n489), .A3(new_n488), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n307), .B2(new_n486), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n502), .B1(new_n508), .B2(G200), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n501), .B1(new_n508), .B2(new_n422), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n475), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n479), .A2(new_n481), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT90), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n479), .A2(new_n481), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT90), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT89), .B1(new_n497), .B2(G190), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n497), .A2(new_n323), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n502), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n514), .A2(new_n515), .A3(new_n518), .A4(new_n475), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n500), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n298), .A2(G257), .A3(new_n305), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n431), .A2(G264), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n343), .A2(G303), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n307), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n504), .A2(G270), .A3(new_n317), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n506), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n415), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n360), .A2(new_n459), .A3(new_n477), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n273), .A2(G1), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(G20), .A3(new_n459), .ZN(new_n532));
  AOI21_X1  g0332(.A(G20), .B1(G33), .B2(G283), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n409), .A2(G97), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(G20), .B2(new_n459), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n260), .A2(KEYINPUT20), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT20), .B1(new_n260), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n529), .B(KEYINPUT21), .C1(new_n530), .C2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n527), .B1(new_n524), .B2(new_n307), .ZN(new_n540));
  OAI211_X1 g0340(.A(G179), .B(new_n540), .C1(new_n530), .C2(new_n538), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT21), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n530), .A2(new_n538), .ZN(new_n544));
  INV_X1    g0344(.A(new_n529), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n540), .A2(G190), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n544), .B(new_n547), .C1(new_n323), .C2(new_n540), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n542), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  AOI211_X1 g0349(.A(new_n274), .B(new_n477), .C1(new_n282), .C2(new_n283), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n210), .B1(new_n347), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(G97), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n410), .A2(new_n553), .A3(new_n433), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n210), .B(G68), .C1(new_n341), .C2(new_n342), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n551), .B1(new_n268), .B2(new_n553), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(new_n262), .A3(new_n263), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n443), .A2(new_n274), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n561), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT87), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n550), .A2(G87), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n311), .A2(new_n489), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT85), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n311), .A2(KEYINPUT85), .A3(new_n489), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT86), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n491), .A2(G250), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n307), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n317), .A2(KEYINPUT86), .A3(G250), .A4(new_n491), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n411), .A2(new_n337), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n460), .B1(new_n431), .B2(G244), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n317), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n323), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n568), .A2(new_n569), .B1(new_n573), .B2(new_n574), .ZN(new_n582));
  OAI211_X1 g0382(.A(G244), .B(G1698), .C1(new_n341), .C2(new_n342), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n409), .B2(new_n459), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n307), .B1(new_n584), .B2(new_n577), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n422), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n359), .B(new_n478), .C1(new_n264), .C2(new_n265), .ZN(new_n588));
  INV_X1    g0388(.A(new_n562), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n588), .A2(new_n443), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n582), .A2(new_n330), .A3(new_n585), .ZN(new_n592));
  AOI21_X1  g0392(.A(G169), .B1(new_n582), .B2(new_n585), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n565), .A2(new_n587), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(G244), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n411), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT4), .ZN(new_n598));
  OAI211_X1 g0398(.A(G250), .B(G1698), .C1(new_n341), .C2(new_n342), .ZN(new_n599));
  INV_X1    g0399(.A(G283), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n409), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT4), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n411), .B2(new_n596), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n598), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n307), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n504), .A2(G257), .A3(new_n317), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n607), .A2(KEYINPUT83), .A3(new_n506), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT83), .B1(new_n607), .B2(new_n506), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT84), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(new_n506), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT83), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n607), .A2(new_n506), .A3(KEYINPUT83), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT84), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n606), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n476), .A2(G97), .A3(new_n359), .A4(new_n478), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT7), .B1(new_n343), .B2(new_n210), .ZN(new_n620));
  INV_X1    g0420(.A(new_n389), .ZN(new_n621));
  OAI21_X1  g0421(.A(G107), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n553), .A2(new_n433), .A3(KEYINPUT6), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT6), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G97), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n433), .A2(KEYINPUT82), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT82), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G107), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n623), .A2(new_n625), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n623), .A2(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n630));
  OAI21_X1  g0430(.A(G20), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n270), .A2(G77), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n622), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n633), .A2(new_n398), .B1(new_n553), .B2(new_n274), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n619), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n601), .B1(KEYINPUT4), .B2(new_n597), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n317), .B1(new_n636), .B2(new_n604), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n614), .A2(new_n615), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n637), .A2(new_n638), .A3(new_n422), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n618), .A2(new_n635), .A3(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n330), .B(new_n606), .C1(new_n611), .C2(new_n616), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n619), .A2(new_n634), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n415), .B1(new_n637), .B2(new_n638), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n595), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n458), .A2(new_n520), .A3(new_n549), .A4(new_n647), .ZN(G372));
  AND3_X1   g0448(.A1(new_n406), .A2(new_n417), .A3(new_n420), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n420), .B1(new_n406), .B2(new_n417), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n380), .A2(new_n378), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n379), .B1(new_n373), .B2(G169), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n382), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(new_n452), .ZN(new_n655));
  INV_X1    g0455(.A(new_n375), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n427), .A2(new_n428), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n651), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT93), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n328), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(new_n333), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n513), .A2(new_n519), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT91), .B1(new_n664), .B2(new_n646), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n610), .B1(new_n608), .B2(new_n609), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n614), .A2(KEYINPUT84), .A3(new_n615), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n323), .B1(new_n668), .B2(new_n606), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n669), .A2(new_n643), .A3(new_n639), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n513), .A2(new_n519), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT91), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n672), .A2(new_n673), .A3(new_n674), .A4(new_n595), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n542), .A2(new_n546), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n482), .A2(new_n499), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n678), .A2(KEYINPUT92), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(KEYINPUT92), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n665), .A2(new_n675), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n591), .A2(new_n594), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT26), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n564), .A2(new_n562), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n284), .A2(G87), .A3(new_n478), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n587), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n685), .B1(new_n689), .B2(new_n645), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n595), .A2(new_n671), .A3(KEYINPUT26), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n684), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n682), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n458), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n663), .A2(new_n694), .ZN(G369));
  NAND2_X1  g0495(.A1(new_n531), .A2(new_n210), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n544), .A2(new_n702), .ZN(new_n703));
  MUX2_X1   g0503(.A(new_n549), .B(new_n676), .S(new_n703), .Z(new_n704));
  INV_X1    g0504(.A(KEYINPUT94), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n482), .A2(new_n701), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n520), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n500), .A2(new_n701), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n706), .A2(G330), .A3(new_n711), .ZN(new_n712));
  OR3_X1    g0512(.A1(new_n679), .A2(new_n680), .A3(new_n701), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n520), .A2(new_n676), .A3(new_n702), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n213), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n554), .A2(G116), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n220), .B2(new_n720), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n540), .A2(G179), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT95), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n637), .A2(new_n638), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n540), .A2(KEYINPUT95), .A3(G179), .ZN(new_n730));
  AND4_X1   g0530(.A1(new_n487), .A2(new_n582), .A3(new_n505), .A4(new_n585), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n732), .A2(KEYINPUT96), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n733), .B1(new_n732), .B2(KEYINPUT96), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n540), .A2(G179), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n508), .B1(new_n585), .B2(new_n582), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n617), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n734), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n725), .B1(new_n739), .B2(new_n702), .ZN(new_n740));
  INV_X1    g0540(.A(new_n734), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n732), .A2(KEYINPUT96), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n738), .B1(new_n742), .B2(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n647), .A2(new_n520), .A3(new_n549), .A4(new_n702), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n740), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT29), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT97), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n693), .B2(new_n702), .ZN(new_n752));
  AOI211_X1 g0552(.A(KEYINPUT97), .B(new_n701), .C1(new_n682), .C2(new_n692), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n542), .A2(new_n678), .A3(new_n546), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n672), .A2(new_n673), .A3(new_n595), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n692), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(KEYINPUT29), .A3(new_n702), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n749), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n724), .B1(new_n759), .B2(G1), .ZN(G364));
  NOR2_X1   g0560(.A1(new_n273), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n209), .B1(new_n761), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n719), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n706), .B2(G330), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G330), .B2(new_n706), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT98), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n704), .A2(G20), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n718), .A2(new_n343), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n773), .A2(G355), .B1(new_n459), .B2(new_n718), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n718), .A2(new_n305), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G45), .B2(new_n220), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n254), .A2(new_n313), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n771), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n216), .B1(G20), .B2(new_n415), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n764), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n210), .A2(new_n422), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n323), .A2(G179), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G87), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT99), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n330), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n210), .A2(G190), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n792), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n793), .A2(new_n384), .B1(new_n795), .B2(new_n205), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G179), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(KEYINPUT32), .A3(G159), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT32), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n798), .B2(new_n387), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n791), .A2(new_n796), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n790), .B(new_n803), .C1(new_n791), .C2(new_n796), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n794), .A2(new_n785), .ZN(new_n805));
  NOR4_X1   g0605(.A1(new_n210), .A2(new_n330), .A3(new_n422), .A4(new_n323), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n305), .B1(new_n805), .B2(new_n433), .C1(new_n807), .C2(new_n202), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n210), .B1(new_n797), .B2(G190), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n553), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n210), .A2(new_n330), .A3(new_n323), .A4(G190), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n250), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n804), .A2(new_n808), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT101), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n789), .A2(G303), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n343), .B1(new_n795), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT33), .B(G317), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n811), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n809), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n806), .A2(G326), .B1(new_n822), .B2(G294), .ZN(new_n823));
  INV_X1    g0623(.A(G322), .ZN(new_n824));
  INV_X1    g0624(.A(G329), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n793), .A2(new_n824), .B1(new_n798), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n805), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(G283), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n817), .A2(new_n821), .A3(new_n823), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n815), .A2(KEYINPUT101), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n816), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n782), .B(new_n783), .C1(new_n831), .C2(new_n780), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n768), .A2(new_n769), .B1(new_n772), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n449), .A2(new_n701), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n455), .A2(new_n835), .B1(new_n450), .B2(new_n451), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT104), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n450), .A2(new_n451), .A3(new_n702), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n839), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT104), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n752), .B2(new_n753), .ZN(new_n845));
  INV_X1    g0645(.A(new_n693), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n452), .A2(new_n455), .A3(new_n702), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n764), .B1(new_n848), .B2(new_n748), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n748), .B2(new_n848), .ZN(new_n850));
  INV_X1    g0650(.A(new_n793), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G294), .ZN(new_n852));
  INV_X1    g0652(.A(new_n795), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G116), .A2(new_n853), .B1(new_n827), .B2(G87), .ZN(new_n854));
  INV_X1    g0654(.A(new_n789), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n852), .B(new_n854), .C1(new_n855), .C2(new_n433), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n343), .B1(new_n798), .B2(new_n818), .ZN(new_n857));
  INV_X1    g0657(.A(G303), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n807), .A2(new_n858), .B1(new_n812), .B2(new_n600), .ZN(new_n859));
  NOR4_X1   g0659(.A1(new_n856), .A2(new_n810), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT102), .ZN(new_n861));
  XOR2_X1   g0661(.A(KEYINPUT103), .B(G143), .Z(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n851), .A2(new_n863), .B1(new_n853), .B2(G159), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  INV_X1    g0665(.A(G150), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n864), .B1(new_n865), .B2(new_n807), .C1(new_n866), .C2(new_n812), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT34), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n855), .A2(new_n202), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n343), .B1(new_n827), .B2(G68), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n872), .B1(new_n384), .B2(new_n809), .C1(new_n873), .C2(new_n798), .ZN(new_n874));
  NOR4_X1   g0674(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n780), .B1(new_n861), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n780), .A2(new_n770), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n783), .B1(new_n205), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n837), .A2(new_n839), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n876), .B(new_n878), .C1(new_n880), .C2(new_n771), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n850), .A2(new_n881), .ZN(G384));
  NOR2_X1   g0682(.A1(new_n629), .A2(new_n630), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n459), .B(new_n218), .C1(new_n884), .C2(KEYINPUT35), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(KEYINPUT35), .B2(new_n884), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT36), .Z(new_n887));
  OR3_X1    g0687(.A1(new_n220), .A2(new_n205), .A3(new_n385), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n209), .B(G13), .C1(new_n888), .C2(new_n249), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n699), .B1(new_n649), .B2(new_n650), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n382), .A2(new_n701), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n654), .A2(new_n656), .A3(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n382), .B(new_n701), .C1(new_n381), .C2(new_n375), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n847), .B1(new_n682), .B2(new_n692), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n841), .ZN(new_n897));
  INV_X1    g0697(.A(new_n699), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n476), .B1(KEYINPUT16), .B2(new_n396), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n405), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n429), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT105), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n359), .B1(new_n264), .B2(new_n265), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n267), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n900), .A2(new_n899), .B1(new_n906), .B2(new_n404), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n425), .B1(new_n907), .B2(new_n699), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n414), .A2(new_n416), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n904), .B(KEYINPUT37), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n406), .A2(new_n898), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n418), .A2(new_n912), .A3(new_n913), .A4(new_n425), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n902), .A2(new_n898), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n902), .A2(new_n417), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n917), .A3(new_n425), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n904), .B1(new_n918), .B2(KEYINPUT37), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n903), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT38), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n903), .B(KEYINPUT38), .C1(new_n915), .C2(new_n919), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n891), .B1(new_n897), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT106), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n418), .A2(new_n912), .A3(new_n425), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(new_n913), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n912), .B1(new_n651), .B2(new_n657), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n921), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n923), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n923), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n381), .A2(new_n382), .A3(new_n702), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT106), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n939), .B(new_n891), .C1(new_n897), .C2(new_n924), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n926), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n754), .A2(new_n458), .A3(new_n758), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n942), .A2(new_n663), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n941), .B(new_n943), .Z(new_n944));
  INV_X1    g0744(.A(G330), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n879), .B1(new_n893), .B2(new_n894), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n931), .A2(new_n747), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n946), .A2(new_n747), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n922), .A2(new_n923), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n947), .A2(KEYINPUT40), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n458), .A2(new_n747), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n945), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n944), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n209), .B2(new_n761), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n944), .A2(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n890), .B1(new_n957), .B2(new_n958), .ZN(G367));
  OAI21_X1  g0759(.A(new_n672), .B1(new_n635), .B2(new_n702), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n671), .A2(new_n701), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n677), .A2(new_n701), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n520), .A3(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT42), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n645), .B1(new_n960), .B2(new_n678), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n964), .A2(KEYINPUT42), .B1(new_n702), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n595), .B1(new_n565), .B2(new_n702), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n683), .A2(new_n565), .A3(new_n702), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n965), .A2(new_n967), .B1(KEYINPUT43), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n712), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n962), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n973), .B(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n719), .B(KEYINPUT41), .Z(new_n977));
  NAND3_X1  g0777(.A1(new_n962), .A2(new_n713), .A3(new_n714), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT45), .Z(new_n979));
  INV_X1    g0779(.A(KEYINPUT44), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n716), .B2(new_n962), .ZN(new_n981));
  INV_X1    g0781(.A(new_n962), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(KEYINPUT44), .A3(new_n715), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n974), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n704), .A2(KEYINPUT94), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n704), .A2(KEYINPUT94), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(G330), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n714), .B1(new_n711), .B2(new_n963), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n989), .B(new_n990), .Z(new_n991));
  NAND3_X1  g0791(.A1(new_n979), .A2(new_n712), .A3(new_n984), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n759), .A2(new_n986), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n977), .B1(new_n993), .B2(new_n759), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n976), .B1(new_n763), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n781), .B1(new_n213), .B2(new_n443), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n775), .B2(new_n238), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n789), .A2(KEYINPUT46), .A3(G116), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT107), .Z(new_n999));
  INV_X1    g0799(.A(KEYINPUT46), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n855), .B2(new_n459), .ZN(new_n1001));
  INV_X1    g0801(.A(G317), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n795), .A2(new_n600), .B1(new_n798), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G97), .B2(new_n827), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n343), .B1(new_n793), .B2(new_n858), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G294), .B2(new_n811), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n806), .A2(G311), .B1(new_n822), .B2(G107), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1001), .A2(new_n1004), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n809), .A2(new_n250), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n343), .B1(new_n799), .B2(G137), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n827), .A2(G77), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(new_n866), .C2(new_n793), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1009), .B(new_n1012), .C1(new_n806), .C2(new_n863), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n384), .B2(new_n855), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n853), .A2(G50), .B1(new_n811), .B2(G159), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT108), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n999), .A2(new_n1008), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT47), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n783), .B(new_n997), .C1(new_n1018), .C2(new_n780), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n779), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n970), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n995), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT109), .Z(G387));
  INV_X1    g0823(.A(new_n721), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n773), .A2(new_n1024), .B1(new_n433), .B2(new_n718), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n244), .A2(new_n313), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n267), .A2(new_n202), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT50), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n721), .B(new_n313), .C1(new_n250), .C2(new_n205), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n775), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1025), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n783), .B1(new_n1031), .B2(new_n781), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n855), .A2(new_n205), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n305), .B1(new_n805), .B2(new_n553), .C1(new_n807), .C2(new_n387), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n809), .A2(new_n443), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n812), .B2(new_n403), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G50), .A2(new_n851), .B1(new_n799), .B2(G150), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n250), .B2(new_n795), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT110), .Z(new_n1040));
  AOI22_X1  g0840(.A1(new_n789), .A2(G294), .B1(G283), .B2(new_n822), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n793), .A2(new_n1002), .B1(new_n795), .B2(new_n858), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1043), .A2(KEYINPUT111), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(KEYINPUT111), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G322), .A2(new_n806), .B1(new_n811), .B2(G311), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1041), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT112), .Z(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(KEYINPUT49), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n305), .B1(new_n799), .B2(G326), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n459), .B2(new_n805), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n1050), .B2(KEYINPUT49), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1040), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n780), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1032), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n710), .B2(new_n779), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n991), .B2(new_n763), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n759), .A2(new_n991), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n719), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n759), .A2(new_n991), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(G393));
  NAND2_X1  g0863(.A1(new_n986), .A2(new_n992), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1065), .A2(new_n719), .A3(new_n993), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT116), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1065), .A2(KEYINPUT116), .A3(new_n719), .A4(new_n993), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1064), .A2(new_n762), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n982), .A2(new_n779), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n775), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n781), .B1(new_n553), .B2(new_n213), .C1(new_n1073), .C2(new_n248), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n764), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n851), .A2(G159), .B1(new_n806), .B2(G150), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n855), .A2(new_n250), .B1(new_n798), .B2(new_n862), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(KEYINPUT113), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(KEYINPUT113), .B2(new_n1078), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n267), .A2(new_n853), .B1(new_n811), .B2(G50), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1081), .A2(KEYINPUT114), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(KEYINPUT114), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n305), .B1(new_n805), .B2(new_n410), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G77), .B2(new_n822), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n343), .B1(new_n798), .B2(new_n824), .C1(new_n433), .C2(new_n805), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n789), .B2(G283), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT115), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n807), .A2(new_n1002), .B1(new_n818), .B2(new_n793), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n811), .A2(G303), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G294), .A2(new_n853), .B1(new_n822), .B2(G116), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1080), .A2(new_n1086), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1075), .B1(new_n1095), .B2(new_n780), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1071), .B1(new_n1072), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1070), .A2(new_n1097), .ZN(G390));
  NAND2_X1  g0898(.A1(new_n458), .A2(new_n749), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n942), .A2(new_n663), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n946), .A2(new_n747), .A3(G330), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n701), .B(new_n836), .C1(new_n692), .C2(new_n756), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n895), .B1(new_n1103), .B2(new_n841), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT117), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n937), .B1(new_n923), .B2(new_n930), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1105), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n897), .A2(new_n936), .B1(new_n933), .B2(new_n934), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1102), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n931), .A2(new_n936), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n893), .A2(new_n894), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n757), .A2(new_n702), .A3(new_n837), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n839), .ZN(new_n1115));
  OAI21_X1  g0915(.A(KEYINPUT117), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1104), .A2(new_n1106), .A3(new_n1105), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n897), .A2(new_n936), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n933), .A2(new_n934), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1118), .A2(new_n1121), .A3(new_n1101), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n843), .A2(new_n747), .A3(G330), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1113), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1103), .A2(new_n841), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n1101), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n747), .A2(G330), .A3(new_n880), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n749), .A2(new_n946), .B1(new_n1127), .B2(new_n1113), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n896), .A2(new_n841), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1100), .A2(new_n1111), .A3(new_n1122), .A4(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1130), .A2(new_n942), .A3(new_n663), .A4(new_n1099), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1118), .A2(new_n1121), .A3(new_n1101), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1101), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1131), .A2(new_n1135), .A3(new_n719), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1111), .A2(new_n763), .A3(new_n1122), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT119), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n783), .B1(new_n403), .B2(new_n877), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G116), .A2(new_n851), .B1(new_n799), .B2(G294), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n790), .B(new_n1140), .C1(new_n553), .C2(new_n795), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n305), .B1(new_n827), .B2(G68), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n205), .B2(new_n809), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n807), .A2(new_n600), .B1(new_n812), .B2(new_n433), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n789), .A2(G150), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT53), .Z(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT54), .B(G143), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n793), .A2(new_n873), .B1(new_n795), .B2(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n812), .A2(new_n865), .B1(new_n809), .B2(new_n387), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(G128), .C2(new_n806), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n305), .B1(new_n805), .B2(new_n202), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G125), .B2(new_n799), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1145), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1139), .B1(new_n1056), .B2(new_n1156), .C1(new_n935), .C2(new_n771), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1137), .A2(new_n1138), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1138), .B1(new_n1137), .B2(new_n1157), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1136), .B1(new_n1158), .B2(new_n1159), .ZN(G378));
  NAND2_X1  g0960(.A1(new_n288), .A2(new_n898), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n329), .B2(new_n333), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n333), .B(new_n1161), .C1(new_n326), .C2(new_n327), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1165), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1164), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n1162), .B2(new_n1168), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n951), .B2(new_n945), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n949), .A2(new_n950), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n946), .A2(new_n747), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n948), .B1(new_n1174), .B2(new_n931), .ZN(new_n1175));
  OAI211_X1 g0975(.A(G330), .B(new_n1172), .C1(new_n1173), .C2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1177), .A2(new_n941), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n925), .A2(KEYINPUT106), .B1(new_n935), .B2(new_n937), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n940), .A2(new_n1179), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT57), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n942), .A2(new_n663), .A3(new_n1099), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1183), .B2(new_n1130), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n719), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1131), .A2(new_n1100), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1177), .A2(new_n941), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1179), .A2(new_n1171), .A3(new_n940), .A4(new_n1176), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT57), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1185), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n305), .A2(G41), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(G33), .A2(G41), .ZN(new_n1193));
  OR3_X1    g0993(.A1(new_n1192), .A2(G50), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1192), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n805), .A2(new_n384), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1195), .A2(new_n1009), .A3(new_n1196), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n553), .B2(new_n812), .C1(new_n459), .C2(new_n807), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G107), .A2(new_n851), .B1(new_n799), .B2(G283), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n443), .B2(new_n795), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1033), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1194), .B1(new_n1201), .B2(KEYINPUT58), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT120), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G128), .A2(new_n851), .B1(new_n853), .B2(G137), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n811), .A2(G132), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n806), .A2(G125), .B1(new_n822), .B2(G150), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n855), .B2(new_n1148), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  INV_X1    g1009(.A(G124), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1193), .B1(new_n798), .B2(new_n1210), .C1(new_n387), .C2(new_n805), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1208), .B2(KEYINPUT59), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1209), .A2(new_n1212), .B1(new_n1201), .B2(KEYINPUT58), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1056), .B1(new_n1203), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n877), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n764), .B1(G50), .B2(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(new_n1170), .C2(new_n770), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT121), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n763), .B2(new_n1189), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1191), .A2(new_n1219), .ZN(G375));
  INV_X1    g1020(.A(new_n1129), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1127), .A2(new_n1113), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1101), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1125), .A2(new_n1101), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1221), .A2(new_n1223), .B1(new_n1224), .B2(new_n1124), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1182), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT122), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n977), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT122), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1182), .A2(new_n1229), .A3(new_n1225), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1132), .A4(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT123), .B1(new_n1225), .B2(new_n762), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n764), .B1(G68), .B2(new_n1215), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G283), .A2(new_n851), .B1(new_n853), .B2(G107), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n858), .B2(new_n798), .C1(new_n855), .C2(new_n553), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G294), .A2(new_n806), .B1(new_n811), .B2(G116), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1236), .A2(new_n343), .A3(new_n1011), .A4(new_n1035), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G150), .A2(new_n853), .B1(new_n799), .B2(G128), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n865), .B2(new_n793), .C1(new_n855), .C2(new_n387), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n806), .A2(G132), .B1(new_n822), .B2(G50), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1196), .A2(new_n343), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n812), .C2(new_n1148), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1235), .A2(new_n1237), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1233), .B1(new_n1243), .B2(new_n780), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n895), .B2(new_n771), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1232), .A2(new_n1245), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1225), .A2(KEYINPUT123), .A3(new_n762), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1231), .A2(new_n1248), .ZN(G381));
  NOR2_X1   g1049(.A1(G387), .A2(G375), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1137), .A2(new_n1157), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT119), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1137), .A2(new_n1138), .A3(new_n1157), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1111), .A2(new_n1122), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n720), .B1(new_n1254), .B2(new_n1132), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1252), .A2(new_n1253), .B1(new_n1131), .B2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n833), .B(new_n1059), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1250), .A2(new_n1256), .A3(new_n1258), .ZN(G407));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n700), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G407), .B(G213), .C1(G375), .C2(new_n1260), .ZN(G409));
  INV_X1    g1061(.A(KEYINPUT127), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G378), .B(new_n1219), .C1(new_n1185), .C2(new_n1190), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1186), .A2(new_n1228), .A3(new_n1189), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1217), .B1(new_n1189), .B2(new_n763), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1256), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1132), .A2(KEYINPUT60), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1227), .A2(new_n1230), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1182), .A2(KEYINPUT60), .A3(new_n1225), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT124), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT124), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1182), .A2(new_n1273), .A3(KEYINPUT60), .A4(new_n1225), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n719), .A3(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G384), .B(new_n1248), .C1(new_n1270), .C2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1227), .A2(new_n1230), .A3(new_n1269), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n720), .B1(new_n1271), .B2(KEYINPUT124), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1274), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G384), .B1(new_n1280), .B2(new_n1248), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(G213), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(G343), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1268), .A2(new_n1282), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1022), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G393), .A2(G396), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT109), .B1(new_n1290), .B2(new_n1257), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(G390), .A2(new_n1291), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1070), .A2(new_n1097), .B1(new_n1290), .B2(new_n1257), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1289), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1290), .A2(new_n1257), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G390), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1296), .B(new_n1022), .C1(G390), .C2(new_n1291), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1294), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1284), .B1(new_n1263), .B2(new_n1267), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1277), .A2(new_n1281), .A3(new_n1287), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1288), .B(new_n1299), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT125), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1280), .A2(new_n1248), .ZN(new_n1307));
  INV_X1    g1107(.A(G384), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT125), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1276), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1284), .A2(G2897), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1306), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1306), .B2(new_n1311), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1300), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1262), .B1(new_n1305), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1314), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1306), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1300), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1294), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1287), .B2(new_n1286), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT126), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1320), .A2(new_n1322), .A3(new_n1326), .A4(KEYINPUT127), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1316), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1329));
  OR2_X1    g1129(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1298), .A3(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1329), .B1(new_n1332), .B2(new_n1315), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1328), .A2(new_n1333), .ZN(G405));
  NAND2_X1  g1134(.A1(G375), .A2(new_n1256), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1263), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1336), .B(new_n1282), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1337), .B(new_n1329), .ZN(G402));
endmodule


