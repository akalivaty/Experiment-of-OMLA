//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND3_X1   g036(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n461), .B1(new_n477), .B2(new_n478), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n461), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n480), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT67), .Z(G162));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n462), .B2(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n476), .A2(new_n465), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n487), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n489), .A2(KEYINPUT4), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n461), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n494), .A2(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n510), .A2(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n506), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n510), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n513), .A2(new_n512), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n509), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n524), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n505), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n510), .A2(new_n532), .B1(new_n516), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n505), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n510), .A2(new_n538), .B1(new_n516), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  INV_X1    g121(.A(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n507), .B2(new_n508), .ZN(new_n548));
  INV_X1    g123(.A(G53), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(KEYINPUT68), .B2(KEYINPUT9), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n551), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT69), .B(G65), .Z(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(new_n525), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n501), .A2(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n558), .A2(G651), .B1(G91), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n555), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  INV_X1    g137(.A(G168), .ZN(G286));
  INV_X1    g138(.A(G74), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n501), .A2(new_n564), .A3(new_n502), .ZN(new_n565));
  AOI22_X1  g140(.A1(G49), .A2(new_n548), .B1(new_n565), .B2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n503), .A2(new_n509), .A3(G87), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT70), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT70), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G288));
  AOI22_X1  g148(.A1(new_n559), .A2(G86), .B1(new_n548), .B2(G48), .ZN(new_n574));
  OAI21_X1  g149(.A(G61), .B1(new_n513), .B2(new_n512), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n505), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n510), .A2(new_n582), .B1(new_n516), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G301), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n516), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(G54), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT71), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n592), .B1(new_n510), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n548), .A2(KEYINPUT71), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n525), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n594), .A2(new_n595), .B1(G651), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n591), .A2(KEYINPUT72), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT72), .B1(new_n591), .B2(new_n599), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n588), .B1(new_n603), .B2(new_n587), .ZN(G284));
  AOI21_X1  g179(.A(new_n588), .B1(new_n603), .B2(new_n587), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G297));
  XNOR2_X1  g183(.A(G297), .B(KEYINPUT73), .ZN(G280));
  NOR2_X1   g184(.A1(new_n602), .A2(G559), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G860), .B2(new_n603), .ZN(G148));
  INV_X1    g186(.A(new_n541), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n587), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n610), .B2(new_n587), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n492), .A2(new_n466), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n479), .A2(G135), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT74), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G2105), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n481), .B2(G123), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n619), .A2(new_n627), .A3(new_n628), .ZN(G156));
  INV_X1    g204(.A(G14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  INV_X1    g206(.A(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n631), .B(G2430), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(new_n634), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n640), .ZN(new_n642));
  NAND4_X1  g217(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT14), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n641), .A2(new_n647), .A3(new_n643), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n630), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n641), .A2(new_n647), .A3(new_n643), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n647), .B1(new_n641), .B2(new_n643), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n652), .ZN(new_n657));
  AOI21_X1  g232(.A(KEYINPUT76), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT76), .ZN(new_n659));
  NOR4_X1   g234(.A1(new_n654), .A2(new_n655), .A3(new_n659), .A4(new_n652), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n653), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT77), .Z(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  XOR2_X1   g242(.A(new_n665), .B(KEYINPUT17), .Z(new_n668));
  INV_X1    g243(.A(new_n664), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n663), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n671), .A2(new_n663), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT78), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n669), .B2(new_n668), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(KEYINPUT78), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n667), .B(new_n670), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(KEYINPUT79), .B(KEYINPUT19), .Z(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n682), .B(new_n683), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n687), .B(new_n688), .S(new_n681), .Z(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT80), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n690), .B1(new_n686), .B2(new_n689), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n694), .B1(new_n692), .B2(new_n695), .ZN(new_n698));
  AND3_X1   g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n697), .B1(new_n696), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n481), .A2(G119), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT81), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n707));
  INV_X1    g282(.A(G107), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G2105), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n479), .B2(G131), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT82), .Z(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n704), .B1(new_n713), .B2(new_n703), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT83), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT83), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n715), .A2(new_n718), .A3(new_n716), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G22), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G166), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1971), .ZN(new_n725));
  MUX2_X1   g300(.A(G6), .B(G305), .S(G16), .Z(new_n726));
  XOR2_X1   g301(.A(KEYINPUT32), .B(G1981), .Z(new_n727));
  XOR2_X1   g302(.A(new_n726), .B(new_n727), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n722), .A2(G23), .ZN(new_n729));
  INV_X1    g304(.A(new_n568), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n722), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT33), .B(G1976), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n731), .B(new_n732), .Z(new_n733));
  NOR3_X1   g308(.A1(new_n725), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT34), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n722), .A2(G24), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n585), .B2(new_n722), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1986), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n734), .B2(new_n735), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n720), .A2(new_n721), .A3(new_n736), .A4(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n742));
  OR3_X1    g317(.A1(new_n741), .A2(KEYINPUT84), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT84), .B(KEYINPUT36), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G4), .A2(G16), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n603), .B2(G16), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G1348), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n703), .A2(G33), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n479), .A2(G139), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n751), .B(new_n752), .C1(new_n461), .C2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT86), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n749), .B1(new_n755), .B2(new_n703), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(G2072), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(G2072), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n703), .B1(new_n759), .B2(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n759), .B2(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G160), .B2(G29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G2084), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT87), .Z(new_n764));
  NAND3_X1  g339(.A1(new_n757), .A2(new_n758), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n703), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n703), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT29), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n765), .B1(G2090), .B2(new_n768), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n748), .B(new_n769), .C1(G2090), .C2(new_n768), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n771));
  AND3_X1   g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n773), .A2(new_n774), .B1(G105), .B2(new_n466), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n479), .A2(G141), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n481), .A2(G129), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n775), .A2(KEYINPUT89), .A3(new_n776), .A4(new_n777), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G32), .B(new_n782), .S(G29), .Z(new_n783));
  XOR2_X1   g358(.A(KEYINPUT27), .B(G1996), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G168), .A2(new_n722), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n722), .B2(G21), .ZN(new_n787));
  INV_X1    g362(.A(G1966), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT90), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n722), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT23), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n607), .B2(new_n722), .ZN(new_n793));
  INV_X1    g368(.A(G1956), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n703), .A2(G26), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT28), .Z(new_n797));
  OAI21_X1  g372(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n798));
  INV_X1    g373(.A(G116), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(G2105), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n481), .B2(G128), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n479), .A2(G140), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT85), .B(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n790), .A2(new_n795), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n541), .A2(G16), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G16), .B2(G19), .ZN(new_n809));
  INV_X1    g384(.A(G1341), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  NOR2_X1   g387(.A1(G171), .A2(new_n722), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G5), .B2(new_n722), .ZN(new_n814));
  OAI221_X1 g389(.A(new_n811), .B1(new_n812), .B2(new_n814), .C1(new_n788), .C2(new_n787), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n812), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n809), .A2(new_n810), .ZN(new_n817));
  INV_X1    g392(.A(G28), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT30), .ZN(new_n819));
  AOI21_X1  g394(.A(G29), .B1(new_n818), .B2(KEYINPUT30), .ZN(new_n820));
  OR2_X1    g395(.A1(KEYINPUT31), .A2(G11), .ZN(new_n821));
  NAND2_X1  g396(.A1(KEYINPUT31), .A2(G11), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n819), .A2(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n626), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G29), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n816), .A2(new_n817), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n762), .A2(G2084), .ZN(new_n828));
  NOR2_X1   g403(.A1(G27), .A2(G29), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G164), .B2(G29), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(G2078), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n827), .B(new_n831), .C1(G2078), .C2(new_n830), .ZN(new_n832));
  NOR4_X1   g407(.A1(new_n770), .A2(new_n785), .A3(new_n807), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n743), .A2(new_n745), .A3(new_n833), .ZN(G150));
  INV_X1    g409(.A(G150), .ZN(G311));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  INV_X1    g411(.A(G67), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n525), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n505), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT93), .B(G93), .Z(new_n842));
  AOI22_X1  g417(.A1(new_n559), .A2(new_n842), .B1(new_n548), .B2(G55), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n603), .A2(G559), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n844), .A2(new_n612), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n841), .A2(new_n541), .A3(new_n843), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n849), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  INV_X1    g430(.A(G860), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n854), .B2(KEYINPUT39), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n846), .B1(new_n855), .B2(new_n857), .ZN(G145));
  OR2_X1    g433(.A1(G164), .A2(new_n803), .ZN(new_n859));
  NAND2_X1  g434(.A1(G164), .A2(new_n803), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n782), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n780), .A2(new_n859), .A3(new_n781), .A4(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n755), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT94), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n862), .A2(new_n866), .A3(new_n754), .A4(new_n863), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n869));
  INV_X1    g444(.A(new_n617), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n711), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n479), .A2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n481), .A2(G130), .ZN(new_n873));
  OR2_X1    g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n874), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n706), .A2(new_n617), .A3(new_n710), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n871), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n877), .B1(new_n871), .B2(new_n878), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n869), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n706), .A2(new_n617), .A3(new_n710), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n617), .B1(new_n706), .B2(new_n710), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n876), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n879), .A3(KEYINPUT95), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n862), .A2(new_n754), .A3(new_n863), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT94), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n868), .A2(new_n887), .A3(KEYINPUT96), .A4(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n865), .A3(new_n867), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n885), .A2(new_n879), .A3(KEYINPUT95), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT95), .B1(new_n885), .B2(new_n879), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n891), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(new_n895), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G160), .ZN(new_n900));
  XNOR2_X1  g475(.A(G162), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n824), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n880), .A2(new_n881), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n892), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n897), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g483(.A1(new_n850), .A2(new_n851), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n610), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n591), .A2(new_n599), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(G299), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n591), .A2(new_n560), .A3(new_n599), .A4(new_n555), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR3_X1    g489(.A1(new_n910), .A2(KEYINPUT97), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n912), .A2(new_n913), .ZN(new_n918));
  XOR2_X1   g493(.A(KEYINPUT98), .B(KEYINPUT41), .Z(new_n919));
  OAI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT97), .B1(new_n910), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n910), .A2(new_n914), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n915), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT42), .ZN(new_n924));
  NAND2_X1  g499(.A1(G290), .A2(new_n568), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n585), .A2(new_n730), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT99), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n928), .ZN(new_n931));
  XOR2_X1   g506(.A(G303), .B(G305), .Z(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OR3_X1    g508(.A1(new_n932), .A2(new_n928), .A3(new_n927), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n915), .B(new_n936), .C1(new_n922), .C2(new_n921), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n924), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n935), .B1(new_n924), .B2(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n844), .A2(new_n587), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(G295));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n941), .ZN(G331));
  NAND3_X1  g518(.A1(G171), .A2(G168), .A3(KEYINPUT100), .ZN(new_n944));
  NAND2_X1  g519(.A1(G171), .A2(KEYINPUT100), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT100), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n531), .B2(new_n534), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(G286), .A3(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n852), .A2(KEYINPUT102), .A3(new_n944), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n944), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n914), .B1(new_n909), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n948), .A2(new_n850), .A3(new_n851), .A4(new_n944), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n949), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n950), .A2(new_n909), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n952), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n920), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT101), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT101), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n920), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n955), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n962), .B2(new_n935), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(new_n935), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n949), .A2(new_n954), .A3(new_n956), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n914), .A2(new_n919), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n916), .B2(new_n914), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n951), .A2(new_n952), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n965), .B(KEYINPUT103), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n966), .B2(new_n968), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(new_n935), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n963), .A2(new_n964), .A3(new_n971), .A4(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n949), .A2(new_n951), .A3(new_n954), .ZN(new_n976));
  INV_X1    g551(.A(new_n961), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n960), .B1(new_n920), .B2(new_n957), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n935), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G37), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n959), .A2(new_n961), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n935), .B1(new_n982), .B2(new_n976), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT43), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n975), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n986));
  INV_X1    g561(.A(new_n983), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(new_n963), .A3(new_n964), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT104), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n963), .A2(new_n971), .A3(new_n974), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n987), .A2(new_n963), .A3(new_n992), .A4(new_n964), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n986), .B1(KEYINPUT44), .B2(new_n994), .ZN(G397));
  NAND2_X1  g570(.A1(new_n492), .A2(new_n493), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n461), .A2(G138), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n477), .B2(new_n478), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT4), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n496), .A2(new_n497), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n481), .B2(G126), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT105), .B(G40), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n468), .A2(new_n473), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1007), .B1(new_n782), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n1008), .B2(new_n782), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n494), .B2(new_n499), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G125), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n490), .B2(new_n491), .ZN(new_n1016));
  INV_X1    g591(.A(new_n472), .ZN(new_n1017));
  OAI21_X1  g592(.A(G2105), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1005), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n464), .A3(new_n467), .A4(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n803), .A2(G2067), .ZN(new_n1022));
  INV_X1    g597(.A(G2067), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n801), .A2(new_n1023), .A3(new_n802), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1010), .B1(KEYINPUT106), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(KEYINPUT106), .B2(new_n1026), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n711), .B(new_n718), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(new_n1007), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1986), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n585), .B(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1030), .B1(new_n1021), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G303), .A2(G8), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT55), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1012), .A2(KEYINPUT107), .A3(new_n1013), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT45), .B(new_n1011), .C1(new_n494), .C2(new_n499), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1006), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT107), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1040), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1020), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(KEYINPUT108), .A4(new_n1037), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT109), .B(G1971), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1012), .A2(KEYINPUT50), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(new_n1011), .C1(new_n494), .C2(new_n499), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1006), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n1051));
  AOI21_X1  g626(.A(G2090), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT110), .B(G8), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1035), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n548), .A2(G49), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n565), .A2(G651), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1057), .A2(new_n567), .A3(new_n1058), .A4(G1976), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n566), .A2(KEYINPUT111), .A3(G1976), .A4(new_n567), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n569), .A2(new_n1065), .A3(new_n571), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1055), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1981), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n574), .A2(new_n1070), .A3(new_n578), .ZN(new_n1071));
  OAI211_X1 g646(.A(G48), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n1072));
  INV_X1    g647(.A(G86), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n516), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n505), .B1(new_n575), .B2(new_n576), .ZN(new_n1075));
  OAI21_X1  g650(.A(G1981), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1071), .A2(KEYINPUT49), .A3(new_n1076), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n1067), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1055), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1012), .B2(new_n1020), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT52), .B1(new_n1083), .B2(new_n1063), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1069), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G8), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1050), .A2(G2090), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1046), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1035), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1038), .A2(new_n1006), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n788), .B1(new_n1004), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G2084), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1047), .A2(new_n1093), .A3(new_n1006), .A4(new_n1049), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1055), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1095), .A2(G168), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1056), .A2(new_n1090), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT63), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1046), .A2(new_n1087), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(G8), .A3(new_n1089), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1103), .A2(KEYINPUT63), .A3(G168), .A4(new_n1082), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1085), .A2(KEYINPUT112), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1069), .A2(new_n1081), .A3(new_n1106), .A4(new_n1084), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1104), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT116), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1101), .A2(G8), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1035), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1113), .A2(new_n1114), .A3(new_n1102), .A4(new_n1108), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1097), .A2(new_n1117), .A3(new_n1098), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1100), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(G168), .A2(new_n1055), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1103), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1121), .B(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1120), .B1(new_n1103), .B2(G8), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(G168), .B2(new_n1055), .ZN(new_n1126));
  OAI22_X1  g701(.A1(new_n1124), .A2(new_n1125), .B1(new_n1095), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1123), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1130));
  AOI21_X1  g705(.A(G2078), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(KEYINPUT53), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1006), .B1(new_n1003), .B2(new_n1048), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1049), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT119), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1047), .A2(new_n1136), .A3(new_n1006), .A4(new_n1049), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(new_n812), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1139), .A2(G2078), .ZN(new_n1140));
  OR3_X1    g715(.A1(new_n1004), .A2(new_n1091), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(G171), .B1(new_n1132), .B2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1129), .A2(new_n1130), .A3(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1056), .A2(new_n1090), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1081), .A2(new_n1065), .A3(new_n572), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1071), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1067), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1102), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT113), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT113), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1152), .B(new_n1148), .C1(new_n1102), .C2(new_n1149), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1144), .A2(new_n1145), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1119), .A2(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1156), .B(G301), .C1(KEYINPUT53), .C2(new_n1131), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1139), .B1(new_n1160), .B2(G2078), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1161), .A2(KEYINPUT123), .A3(G301), .A4(new_n1156), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1138), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1135), .A2(KEYINPUT122), .A3(new_n812), .A4(new_n1137), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(G40), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n900), .A2(new_n1169), .A3(new_n1140), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1170), .A2(new_n1014), .A3(new_n1038), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1168), .B(new_n1171), .C1(KEYINPUT53), .C2(new_n1131), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1164), .B1(new_n1172), .B2(G171), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1163), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1143), .B1(new_n1172), .B2(G171), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1164), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1177), .A2(new_n1056), .A3(new_n1090), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1174), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT57), .ZN(new_n1180));
  XNOR2_X1  g755(.A(G299), .B(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT56), .B(G2072), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1042), .A2(new_n1043), .A3(new_n1037), .A4(new_n1182), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n794), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT117), .B1(new_n1050), .B2(new_n794), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1181), .B(new_n1183), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1050), .A2(new_n794), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT117), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n794), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1181), .B1(new_n1191), .B2(new_n1183), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1012), .A2(new_n1020), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT118), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1023), .ZN(new_n1195));
  INV_X1    g770(.A(G1348), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1135), .A2(new_n1196), .A3(new_n1137), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n602), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1186), .B1(new_n1192), .B2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(KEYINPUT58), .B(G1341), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1042), .A2(new_n1043), .A3(new_n1037), .ZN(new_n1201));
  OAI22_X1  g776(.A1(new_n1194), .A2(new_n1200), .B1(new_n1201), .B2(G1996), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(new_n541), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT59), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1202), .A2(new_n1205), .A3(new_n541), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1186), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1208), .B1(new_n1192), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1181), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1213), .A2(KEYINPUT61), .A3(new_n1186), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1207), .A2(new_n1210), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT120), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g792(.A(new_n1195), .B(new_n1197), .C1(new_n603), .C2(KEYINPUT60), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n603), .A2(KEYINPUT60), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1218), .B(new_n1219), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1207), .A2(new_n1210), .A3(KEYINPUT120), .A4(new_n1214), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1217), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1179), .B1(new_n1199), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1033), .B1(new_n1155), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n1225));
  AND2_X1   g800(.A1(new_n1030), .A2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g801(.A1(new_n1030), .A2(new_n1225), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1021), .A2(new_n1031), .A3(new_n585), .ZN(new_n1228));
  XOR2_X1   g803(.A(new_n1228), .B(KEYINPUT48), .Z(new_n1229));
  NOR3_X1   g804(.A1(new_n1226), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1021), .A2(new_n1008), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT46), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  XOR2_X1   g808(.A(new_n1233), .B(KEYINPUT124), .Z(new_n1234));
  NAND2_X1  g809(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1021), .B1(new_n782), .B2(new_n1025), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  XOR2_X1   g812(.A(new_n1237), .B(KEYINPUT47), .Z(new_n1238));
  NAND3_X1  g813(.A1(new_n1028), .A2(new_n718), .A3(new_n713), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1007), .B1(new_n1239), .B2(new_n1024), .ZN(new_n1240));
  NOR3_X1   g815(.A1(new_n1230), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1224), .A2(new_n1241), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g817(.A(KEYINPUT126), .ZN(new_n1244));
  NOR2_X1   g818(.A1(G227), .A2(new_n459), .ZN(new_n1245));
  AND3_X1   g819(.A1(new_n661), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g820(.A(new_n1244), .B1(new_n661), .B2(new_n1245), .ZN(new_n1247));
  OAI21_X1  g821(.A(new_n701), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g822(.A(new_n1248), .B1(new_n903), .B2(new_n906), .ZN(new_n1249));
  INV_X1    g823(.A(KEYINPUT127), .ZN(new_n1250));
  AND3_X1   g824(.A1(new_n1249), .A2(new_n985), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g825(.A(new_n1250), .B1(new_n1249), .B2(new_n985), .ZN(new_n1252));
  NOR2_X1   g826(.A1(new_n1251), .A2(new_n1252), .ZN(G308));
  NAND2_X1  g827(.A1(new_n1249), .A2(new_n985), .ZN(G225));
endmodule


