//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n621, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n466), .A2(G137), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n471), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n470), .A2(new_n472), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n477), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n469), .B(new_n476), .C1(new_n478), .C2(new_n466), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT68), .Z(G160));
  NAND3_X1  g055(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n466), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n482), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT70), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n472), .A2(new_n475), .A3(new_n494), .A4(new_n473), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n477), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n500));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n466), .A2(G114), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(G102), .A2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(G114), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G2105), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT71), .A4(G2104), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n500), .A2(new_n502), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n499), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(KEYINPUT73), .B1(G75), .B2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n514), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(G543), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(new_n515), .A3(new_n526), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(G50), .A2(new_n528), .B1(new_n530), .B2(G88), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n531), .B1(new_n519), .B2(KEYINPUT74), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n520), .A2(new_n532), .ZN(G166));
  NAND4_X1  g108(.A1(new_n525), .A2(G51), .A3(G543), .A4(new_n526), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n534), .B(new_n536), .C1(new_n529), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n515), .A2(KEYINPUT75), .ZN(new_n539));
  OR2_X1    g114(.A1(KEYINPUT5), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  NAND2_X1  g116(.A1(KEYINPUT5), .A2(G543), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n539), .A2(G63), .A3(G651), .A4(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n538), .B1(new_n546), .B2(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(new_n539), .A2(new_n543), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G64), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n514), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n554), .A2(new_n527), .B1(new_n529), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(G171));
  AOI22_X1  g132(.A1(G43), .A2(new_n528), .B1(new_n530), .B2(G81), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n549), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(new_n528), .A2(G53), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n515), .A2(G65), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT77), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n514), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(G91), .B2(new_n530), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n571), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  NAND2_X1  g153(.A1(new_n546), .A2(new_n547), .ZN(new_n579));
  INV_X1    g154(.A(new_n538), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G286));
  OR2_X1    g156(.A1(new_n520), .A2(new_n532), .ZN(G303));
  NAND4_X1  g157(.A1(new_n525), .A2(G87), .A3(new_n515), .A4(new_n526), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n525), .A2(G49), .A3(G543), .A4(new_n526), .ZN(new_n584));
  AOI21_X1  g159(.A(G74), .B1(new_n539), .B2(new_n543), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n514), .ZN(G288));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n515), .B2(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n587), .B1(new_n589), .B2(new_n514), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n540), .B2(new_n542), .ZN(new_n592));
  OAI211_X1 g167(.A(KEYINPUT78), .B(G651), .C1(new_n592), .C2(new_n588), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n525), .A2(G86), .A3(new_n515), .A4(new_n526), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n525), .A2(G48), .A3(G543), .A4(new_n526), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n594), .A2(new_n597), .ZN(G305));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n599), .A2(new_n527), .B1(new_n529), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n601), .A2(KEYINPUT79), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n601), .A2(KEYINPUT79), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n550), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n602), .A2(new_n603), .B1(new_n514), .B2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n530), .A2(KEYINPUT10), .A3(G92), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n529), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n527), .A2(new_n612), .B1(new_n613), .B2(new_n514), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(G868), .B2(new_n615), .ZN(G284));
  OAI21_X1  g191(.A(new_n606), .B1(G868), .B2(new_n615), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(KEYINPUT80), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n618), .A2(KEYINPUT80), .ZN(new_n620));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(G299), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n619), .B1(new_n620), .B2(new_n622), .ZN(G297));
  AOI21_X1  g198(.A(new_n619), .B1(new_n620), .B2(new_n622), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n615), .B1(new_n625), .B2(G860), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT81), .Z(G148));
  NAND2_X1  g202(.A1(new_n563), .A2(new_n621), .ZN(new_n628));
  INV_X1    g203(.A(new_n615), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n630), .B2(new_n621), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n468), .A2(new_n477), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  INV_X1    g212(.A(G111), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n637), .A2(KEYINPUT82), .B1(new_n638), .B2(G2105), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(KEYINPUT82), .B2(new_n637), .ZN(new_n640));
  INV_X1    g215(.A(G135), .ZN(new_n641));
  INV_X1    g216(.A(G123), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n482), .A2(G2105), .ZN(new_n643));
  OAI221_X1 g218(.A(new_n640), .B1(new_n483), .B2(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n636), .A2(new_n645), .A3(new_n646), .ZN(G156));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT84), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2451), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT86), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2430), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n652), .B(new_n659), .Z(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2454), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT87), .Z(new_n669));
  NOR2_X1   g244(.A1(G2072), .A2(G2078), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n442), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(KEYINPUT17), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n672), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n667), .B(new_n668), .C1(new_n442), .C2(new_n670), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT18), .Z(new_n676));
  NAND3_X1  g251(.A1(new_n669), .A2(new_n673), .A3(new_n667), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  NAND2_X1  g273(.A1(G166), .A2(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G16), .B2(G22), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  MUX2_X1   g278(.A(G6), .B(G305), .S(G16), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(G288), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT33), .B(G1976), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n702), .A2(new_n703), .A3(new_n706), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT34), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G25), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n466), .A2(G107), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n486), .A2(G119), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n484), .A2(G131), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(new_n715), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(KEYINPUT88), .ZN(new_n729));
  MUX2_X1   g304(.A(G24), .B(G290), .S(G16), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1986), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(KEYINPUT89), .B2(KEYINPUT36), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n728), .A2(KEYINPUT88), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n714), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  OR3_X1    g310(.A1(new_n735), .A2(KEYINPUT89), .A3(KEYINPUT36), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(KEYINPUT89), .B2(KEYINPUT36), .ZN(new_n737));
  NOR2_X1   g312(.A1(G171), .A2(new_n707), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G5), .B2(new_n707), .ZN(new_n739));
  INV_X1    g314(.A(G1961), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n715), .A2(G32), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT26), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n468), .A2(G105), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G141), .ZN(new_n749));
  INV_X1    g324(.A(G129), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n748), .B1(new_n483), .B2(new_n749), .C1(new_n750), .C2(new_n643), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n743), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n742), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n707), .A2(G4), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n615), .B2(new_n707), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1348), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n752), .A2(new_n753), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  INV_X1    g338(.A(G139), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n762), .B1(new_n466), .B2(new_n763), .C1(new_n483), .C2(new_n764), .ZN(new_n765));
  MUX2_X1   g340(.A(G33), .B(new_n765), .S(G29), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2072), .ZN(new_n767));
  NAND2_X1  g342(.A1(G160), .A2(G29), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT24), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n715), .B1(new_n769), .B2(G34), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(KEYINPUT93), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(KEYINPUT93), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n769), .A2(G34), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT94), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n768), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n767), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G29), .A2(G35), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G162), .B2(G29), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT29), .B(G2090), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n754), .A2(new_n759), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n739), .A2(new_n740), .ZN(new_n785));
  INV_X1    g360(.A(G2078), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n512), .A2(new_n715), .ZN(new_n787));
  NOR2_X1   g362(.A1(G27), .A2(G29), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT31), .B(G11), .Z(new_n790));
  INV_X1    g365(.A(G28), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(KEYINPUT30), .ZN(new_n792));
  AOI21_X1  g367(.A(G29), .B1(new_n791), .B2(KEYINPUT30), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OR3_X1    g369(.A1(new_n787), .A2(new_n786), .A3(new_n788), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n785), .A2(new_n789), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G1966), .ZN(new_n797));
  NOR2_X1   g372(.A1(G168), .A2(new_n707), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n707), .B2(G21), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n797), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT95), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n707), .A2(G20), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT23), .Z(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G299), .B2(G16), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1956), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G19), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n564), .B2(G16), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT90), .B(G1341), .Z(new_n809));
  AND2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n644), .A2(new_n715), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n800), .A2(new_n802), .A3(new_n806), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n715), .A2(G26), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT28), .Z(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(G116), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G2105), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n484), .B2(G140), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT91), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n486), .B2(G128), .ZN(new_n822));
  INV_X1    g397(.A(G128), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n643), .A2(KEYINPUT91), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n816), .B1(new_n825), .B2(G29), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT92), .B(G2067), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n784), .A2(new_n814), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n736), .A2(new_n737), .A3(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  NAND2_X1  g406(.A1(new_n615), .A2(G559), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT38), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n550), .A2(G67), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n514), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n837), .A2(new_n527), .B1(new_n529), .B2(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n563), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n836), .A2(new_n839), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n564), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n833), .B(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT97), .B(G860), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n842), .A2(new_n848), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  XNOR2_X1  g427(.A(new_n825), .B(G164), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n484), .A2(G142), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n486), .A2(G130), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n466), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n853), .B(new_n858), .Z(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n722), .B(KEYINPUT98), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n634), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n751), .B(new_n765), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n862), .A2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n862), .A2(new_n863), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n859), .A3(new_n864), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n491), .B(G160), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(new_n644), .Z(new_n872));
  AOI21_X1  g447(.A(G37), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n872), .B2(new_n870), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g450(.A1(new_n840), .A2(new_n621), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(G299), .B2(new_n615), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NOR3_X1   g454(.A1(G299), .A2(new_n877), .A3(new_n615), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(G299), .A2(new_n615), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n883), .A2(KEYINPUT100), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(KEYINPUT100), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n841), .A2(new_n843), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n630), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n879), .B2(new_n880), .ZN(new_n891));
  INV_X1    g466(.A(new_n880), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(KEYINPUT101), .A3(new_n878), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n893), .A3(new_n882), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(G299), .B2(new_n615), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n894), .A2(new_n895), .B1(new_n881), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n889), .B1(new_n888), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G166), .B(G305), .ZN(new_n899));
  XNOR2_X1  g474(.A(G290), .B(new_n709), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n899), .B(new_n900), .Z(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(KEYINPUT42), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n898), .B(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n876), .B1(new_n903), .B2(new_n621), .ZN(G295));
  OAI21_X1  g479(.A(new_n876), .B1(new_n903), .B2(new_n621), .ZN(G331));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  OAI21_X1  g481(.A(G286), .B1(G171), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(G301), .A2(KEYINPUT102), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n844), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n844), .A2(new_n908), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  INV_X1    g488(.A(new_n907), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n914), .A3(new_n909), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n915), .A3(new_n883), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n912), .A2(new_n915), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n897), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n901), .ZN(new_n919));
  INV_X1    g494(.A(G37), .ZN(new_n920));
  INV_X1    g495(.A(new_n901), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n921), .B(new_n916), .C1(new_n917), .C2(new_n897), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n912), .A2(new_n915), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n883), .A2(new_n895), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n926), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n891), .A2(new_n893), .A3(new_n896), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n927), .B2(KEYINPUT104), .ZN(new_n931));
  OAI221_X1 g506(.A(new_n901), .B1(new_n886), .B2(new_n926), .C1(new_n929), .C2(new_n931), .ZN(new_n932));
  AND4_X1   g507(.A1(KEYINPUT43), .A2(new_n932), .A3(new_n920), .A4(new_n922), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n925), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n932), .A2(new_n924), .A3(new_n920), .A4(new_n922), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT103), .B1(new_n923), .B2(KEYINPUT43), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n934), .B1(new_n940), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g516(.A(new_n825), .B(G2067), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(G1996), .B2(new_n751), .ZN(new_n943));
  XOR2_X1   g518(.A(KEYINPUT105), .B(G1384), .Z(new_n944));
  INV_X1    g519(.A(new_n505), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT71), .B1(new_n945), .B2(new_n509), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n504), .A2(new_n505), .A3(new_n503), .ZN(new_n947));
  OAI22_X1  g522(.A1(new_n946), .A2(new_n947), .B1(new_n481), .B2(new_n501), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n495), .A2(KEYINPUT4), .B1(new_n477), .B2(new_n497), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(G113), .A2(G2104), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n474), .A2(G2104), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n473), .ZN(new_n956));
  INV_X1    g531(.A(G125), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(G2105), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(G40), .A3(new_n476), .A4(new_n469), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n953), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n943), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1996), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(new_n751), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT108), .Z(new_n967));
  NOR2_X1   g542(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n723), .A2(new_n725), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n722), .A2(new_n726), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n961), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  OR3_X1    g547(.A1(new_n962), .A2(G1986), .A3(G290), .ZN(new_n973));
  NAND3_X1  g548(.A1(G290), .A2(G1986), .A3(new_n961), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n975), .B(KEYINPUT107), .Z(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT45), .B(new_n944), .C1(new_n948), .C2(new_n949), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n512), .A2(KEYINPUT109), .A3(KEYINPUT45), .A4(new_n944), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n948), .B2(new_n949), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n960), .B1(new_n985), .B2(new_n952), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n982), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n983), .B1(new_n982), .B2(new_n986), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n987), .A2(new_n988), .A3(G1971), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n990), .B(new_n984), .C1(new_n948), .C2(new_n949), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n960), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n993), .B2(KEYINPUT112), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n479), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G1384), .B1(new_n499), .B2(new_n511), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n997), .B2(new_n990), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n994), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(G2090), .ZN(new_n1002));
  OAI21_X1  g577(.A(G8), .B1(new_n989), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(G166), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n993), .A2(new_n991), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(G2090), .ZN(new_n1012));
  OAI211_X1 g587(.A(G8), .B(new_n1008), .C1(new_n989), .C2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(G651), .B1(new_n592), .B2(new_n588), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(new_n595), .A3(new_n596), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G1981), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT111), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n594), .A2(new_n1018), .A3(new_n597), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(new_n1020), .A3(G1981), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1017), .A2(new_n1019), .A3(KEYINPUT49), .A4(new_n1021), .ZN(new_n1025));
  OAI21_X1  g600(.A(G8), .B1(new_n985), .B2(new_n960), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1027), .B(new_n1030), .C1(new_n1029), .C2(G288), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G288), .A2(new_n1029), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT113), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n1033), .A4(new_n1031), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n998), .A2(G2084), .A3(new_n992), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n960), .B1(new_n985), .B2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n984), .B(new_n951), .C1(new_n948), .C2(new_n949), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1966), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(G286), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1010), .A2(new_n1013), .A3(new_n1039), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT63), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(G8), .B1(new_n989), .B2(new_n1012), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1009), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1028), .A2(new_n1034), .A3(new_n1048), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1013), .A3(new_n1046), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1013), .A2(new_n1028), .A3(new_n1034), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1036), .A2(new_n1029), .A3(new_n709), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1026), .B1(new_n1056), .B2(new_n1019), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n998), .A2(new_n992), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G1961), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n786), .B1(new_n987), .B2(new_n988), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n479), .B2(new_n995), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n958), .A2(G2105), .B1(G101), .B2(new_n468), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(KEYINPUT119), .A3(G40), .A4(new_n476), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n951), .B1(new_n512), .B2(new_n944), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT120), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n953), .A2(new_n1073), .A3(new_n1069), .A4(new_n1067), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1064), .A2(G2078), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n982), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT121), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1075), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1065), .A2(new_n1082), .A3(G301), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1042), .A2(new_n1076), .A3(new_n1043), .ZN(new_n1084));
  AOI21_X1  g659(.A(G301), .B1(new_n1065), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1060), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n982), .A2(new_n986), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT110), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n982), .A2(new_n983), .A3(new_n986), .ZN(new_n1089));
  AOI21_X1  g664(.A(G2078), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1090), .A2(KEYINPUT53), .B1(G1961), .B2(new_n1061), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1081), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1080), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(G171), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1065), .A2(G301), .A3(new_n1084), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(KEYINPUT54), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(G168), .B2(new_n1006), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1045), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n996), .B(new_n1043), .C1(new_n997), .C2(KEYINPUT45), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n797), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n993), .A2(new_n777), .A3(new_n991), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1006), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(G286), .A2(KEYINPUT117), .A3(G8), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(G168), .B2(new_n1006), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT51), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT118), .B1(new_n1106), .B2(new_n1100), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1102), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G168), .A2(new_n1006), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1086), .A2(new_n1097), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1039), .A2(new_n1013), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1088), .A2(new_n701), .A3(new_n1089), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(G2090), .B2(new_n1001), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1008), .B1(new_n1121), .B2(G8), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1118), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1010), .A2(KEYINPUT122), .A3(new_n1013), .A4(new_n1039), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1117), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n982), .A2(new_n986), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT114), .ZN(new_n1129));
  INV_X1    g704(.A(G1956), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1129), .B1(new_n1001), .B2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g706(.A(KEYINPUT114), .B(G1956), .C1(new_n994), .C2(new_n1000), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1134));
  OR2_X1    g709(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1135));
  AND3_X1   g710(.A1(G299), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(G299), .B2(new_n1134), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1138), .B(new_n1128), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(KEYINPUT61), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1141), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1140), .A2(KEYINPUT116), .A3(KEYINPUT61), .A4(new_n1141), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n985), .A2(new_n960), .ZN(new_n1150));
  INV_X1    g725(.A(G2067), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1061), .B2(G1348), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1153), .A2(new_n615), .ZN(new_n1154));
  INV_X1    g729(.A(G1348), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1011), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n629), .B1(new_n1156), .B2(new_n1152), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT60), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n629), .A2(KEYINPUT60), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1158), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT58), .B(G1341), .ZN(new_n1161));
  OAI22_X1  g736(.A1(new_n1087), .A2(G1996), .B1(new_n1150), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n564), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT59), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1160), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1144), .A2(new_n1148), .A3(new_n1149), .A4(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1146), .B1(new_n1141), .B2(new_n1157), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1059), .B1(new_n1126), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1113), .A2(new_n1171), .A3(new_n1115), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1172), .A2(new_n1085), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1173), .A2(new_n1123), .A3(KEYINPUT123), .A4(new_n1124), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1116), .A2(KEYINPUT62), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT124), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n977), .B1(new_n1170), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n961), .B1(new_n942), .B2(new_n751), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT125), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n965), .B(KEYINPUT46), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1185), .A2(KEYINPUT47), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(KEYINPUT47), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n973), .B(KEYINPUT48), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n972), .A2(new_n1189), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n825), .A2(G2067), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1192), .B1(new_n968), .B2(new_n970), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1188), .B(new_n1190), .C1(new_n962), .C2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(KEYINPUT126), .B1(new_n1181), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1126), .A2(new_n1169), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1059), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1196), .A2(new_n1180), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n977), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1190), .B1(new_n962), .B2(new_n1193), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1202), .B1(new_n1187), .B2(new_n1186), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1195), .A2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g780(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n1207), .A2(new_n697), .ZN(new_n1208));
  XNOR2_X1  g782(.A(new_n1208), .B(KEYINPUT127), .ZN(new_n1209));
  OAI211_X1 g783(.A(new_n874), .B(new_n1209), .C1(new_n938), .C2(new_n939), .ZN(G225));
  INV_X1    g784(.A(G225), .ZN(G308));
endmodule


