//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT2), .B(G226), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(G264), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n227), .B(new_n230), .ZN(G358));
  XNOR2_X1  g0031(.A(G50), .B(G58), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  NAND3_X1  g0039(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g0041(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(new_n212), .ZN(new_n243));
  NOR2_X1   g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n203), .A2(G20), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n244), .A2(G50), .A3(new_n245), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n246), .B1(G50), .B2(new_n240), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n204), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n250), .A2(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G50), .A2(G58), .ZN(new_n256));
  INV_X1    g0056(.A(G68), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n204), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n243), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n249), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT9), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n203), .A2(G274), .ZN(new_n262));
  XOR2_X1   g0062(.A(KEYINPUT66), .B(G45), .Z(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT67), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G41), .A2(G45), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G1), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n203), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n265), .B1(G226), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  INV_X1    g0075(.A(G77), .ZN(new_n276));
  OAI22_X1  g0076(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n273), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G1698), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n277), .B1(G222), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n266), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n272), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G190), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(G200), .B2(new_n286), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT70), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT10), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n261), .A2(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n290), .B2(new_n291), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n261), .A2(KEYINPUT70), .A3(KEYINPUT10), .A4(new_n289), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n286), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n260), .B(new_n296), .C1(G179), .C2(new_n286), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n271), .A2(G232), .ZN(new_n300));
  INV_X1    g0100(.A(new_n265), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G87), .ZN(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n273), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G226), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n304), .B1(new_n306), .B2(new_n275), .C1(new_n307), .C2(new_n274), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n266), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT72), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n300), .A2(new_n301), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n303), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n295), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT7), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n273), .A2(new_n314), .A3(G20), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT7), .B1(new_n282), .B2(new_n204), .ZN(new_n316));
  OAI21_X1  g0116(.A(G68), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n253), .A2(G159), .ZN(new_n318));
  INV_X1    g0118(.A(G58), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n257), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G58), .A2(G68), .ZN(new_n321));
  OAI21_X1  g0121(.A(G20), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n317), .A2(KEYINPUT16), .A3(new_n318), .A4(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT16), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n314), .B1(new_n273), .B2(G20), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n257), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n318), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n323), .A2(new_n329), .A3(new_n243), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n250), .B1(new_n203), .B2(G20), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(new_n244), .B1(new_n241), .B2(new_n250), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n303), .A2(new_n309), .A3(new_n334), .A4(new_n311), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n313), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT18), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n312), .A2(new_n295), .B1(new_n330), .B2(new_n332), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT18), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n339), .A3(new_n335), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n333), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n312), .A2(G200), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n303), .A2(new_n309), .A3(G190), .A4(new_n311), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT17), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n342), .A2(KEYINPUT17), .A3(new_n343), .A4(new_n344), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n265), .B1(G244), .B2(new_n271), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n273), .A2(G238), .A3(G1698), .ZN(new_n351));
  INV_X1    g0151(.A(G107), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n273), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(G232), .B2(new_n283), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n350), .B1(new_n354), .B2(new_n285), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(G179), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT69), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n250), .A2(new_n254), .B1(new_n204), .B2(new_n276), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n251), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n243), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n244), .A2(G77), .A3(new_n245), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(G77), .C2(new_n240), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT69), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n355), .B2(new_n295), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n366), .A2(new_n356), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n363), .B1(new_n355), .B2(G200), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n287), .B2(new_n355), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n299), .A2(new_n341), .A3(new_n349), .A4(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT14), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT13), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n273), .A2(G232), .A3(G1698), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G97), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n375), .B(new_n376), .C1(new_n306), .C2(new_n307), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n266), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT71), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(new_n380), .A3(new_n266), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n265), .B1(G238), .B2(new_n271), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n374), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n377), .A2(new_n380), .A3(new_n266), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n380), .B1(new_n377), .B2(new_n266), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n374), .B(new_n383), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n373), .B(G169), .C1(new_n384), .C2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT13), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(G179), .A3(new_n387), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n387), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n373), .B1(new_n394), .B2(G169), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n253), .A2(G50), .B1(G20), .B2(new_n257), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n276), .B2(new_n251), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT11), .B1(new_n397), .B2(new_n243), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n241), .A2(new_n257), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT12), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(KEYINPUT11), .A3(new_n243), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n244), .A2(G68), .A3(new_n245), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n393), .A2(new_n395), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n394), .A2(G200), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n403), .A2(new_n398), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n405), .B(new_n406), .C1(new_n287), .C2(new_n394), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n372), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n279), .A2(new_n281), .A3(G250), .A4(new_n305), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT86), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT86), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n273), .A2(new_n413), .A3(G250), .A4(new_n305), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT87), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n279), .A2(new_n281), .A3(G257), .A4(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G294), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n416), .B1(new_n415), .B2(new_n419), .ZN(new_n422));
  OAI211_X1 g0222(.A(KEYINPUT88), .B(new_n266), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT75), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n203), .A2(G45), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT74), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT74), .ZN(new_n428));
  INV_X1    g0228(.A(G45), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G1), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT5), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G41), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n424), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT74), .B1(new_n425), .B2(new_n426), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n430), .A2(new_n428), .A3(new_n432), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(KEYINPUT75), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n285), .A2(G274), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(G264), .A3(new_n285), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n423), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n415), .A2(new_n419), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT87), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n420), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT88), .B1(new_n450), .B2(new_n266), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT89), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n266), .B1(new_n421), .B2(new_n422), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT88), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT89), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(new_n423), .A4(new_n446), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n287), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n446), .A2(new_n453), .ZN(new_n459));
  INV_X1    g0259(.A(G200), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n204), .A2(G107), .ZN(new_n463));
  INV_X1    g0263(.A(G13), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(KEYINPUT85), .A3(KEYINPUT25), .ZN(new_n467));
  OR2_X1    g0267(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n463), .A2(new_n465), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n203), .A2(G33), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n240), .A2(new_n471), .A3(new_n212), .A4(new_n242), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n467), .B(new_n470), .C1(new_n352), .C2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n273), .A2(new_n204), .A3(G87), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT22), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G116), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n463), .A2(KEYINPUT23), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n463), .A2(KEYINPUT23), .ZN(new_n478));
  OAI221_X1 g0278(.A(new_n475), .B1(G20), .B2(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n479), .B(KEYINPUT24), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n473), .B1(new_n480), .B2(new_n243), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n462), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n243), .ZN(new_n483));
  INV_X1    g0283(.A(new_n473), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n295), .B1(new_n452), .B2(new_n457), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n446), .A2(new_n453), .A3(G179), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n273), .A2(G264), .A3(G1698), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n273), .A2(G257), .A3(new_n305), .ZN(new_n491));
  INV_X1    g0291(.A(G303), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n490), .B(new_n491), .C1(new_n492), .C2(new_n273), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n266), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n443), .A2(G270), .A3(new_n285), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n442), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  INV_X1    g0297(.A(G97), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n204), .C1(G33), .C2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n499), .B(new_n243), .C1(new_n204), .C2(G116), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT20), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n240), .A2(G116), .ZN(new_n503));
  INV_X1    g0303(.A(new_n472), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n496), .A2(new_n506), .A3(G169), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT83), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n507), .B(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n506), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n442), .A2(G179), .A3(new_n494), .A4(new_n495), .ZN(new_n512));
  OR3_X1    g0312(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT82), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT82), .B1(new_n511), .B2(new_n512), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n506), .B1(new_n496), .B2(G200), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n517), .A2(KEYINPUT84), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(KEYINPUT84), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n496), .A2(new_n287), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n482), .A2(new_n489), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n443), .A2(G257), .A3(new_n285), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT76), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n443), .A2(KEYINPUT76), .A3(G257), .A4(new_n285), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n442), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT77), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  INV_X1    g0332(.A(G244), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n306), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G250), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n497), .B1(new_n274), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n532), .B1(new_n306), .B2(new_n533), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n285), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G179), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n528), .A2(KEYINPUT77), .A3(new_n442), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n531), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n243), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n253), .A2(G77), .ZN(new_n544));
  XOR2_X1   g0344(.A(new_n544), .B(KEYINPUT73), .Z(new_n545));
  NAND3_X1  g0345(.A1(new_n352), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  XOR2_X1   g0346(.A(G97), .B(G107), .Z(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(KEYINPUT6), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n548), .B2(G20), .ZN(new_n549));
  OAI21_X1  g0349(.A(G107), .B1(new_n315), .B2(new_n316), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n241), .A2(new_n498), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n472), .B2(new_n498), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n440), .B1(new_n434), .B2(new_n437), .ZN(new_n556));
  AOI211_X1 g0356(.A(new_n530), .B(new_n556), .C1(new_n526), .C2(new_n527), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT77), .B1(new_n528), .B2(new_n442), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n557), .A2(new_n558), .A3(new_n539), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n542), .B(new_n555), .C1(new_n559), .C2(G169), .ZN(new_n560));
  INV_X1    g0360(.A(new_n539), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n531), .A2(G190), .A3(new_n541), .A4(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n554), .B(new_n562), .C1(new_n559), .C2(new_n460), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n359), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n240), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n279), .A2(new_n281), .A3(new_n204), .A4(G68), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n204), .B1(new_n376), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  INV_X1    g0370(.A(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n204), .A2(G33), .A3(G97), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT79), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n574), .A2(new_n575), .A3(new_n568), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n575), .B1(new_n574), .B2(new_n568), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n567), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n543), .B1(new_n578), .B2(KEYINPUT80), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n568), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n574), .A2(new_n575), .A3(new_n568), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT80), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(new_n567), .A4(new_n573), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n566), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n279), .A2(new_n281), .A3(G238), .A4(new_n305), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n279), .A2(new_n281), .A3(G244), .A4(G1698), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n476), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n266), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n535), .A2(KEYINPUT78), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n430), .B1(new_n591), .B2(G274), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n426), .A2(KEYINPUT78), .A3(G250), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n266), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n590), .A2(new_n595), .A3(new_n287), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n594), .B1(new_n266), .B2(new_n589), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(G200), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n504), .A2(G87), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n586), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n472), .A2(new_n359), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT81), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n590), .A2(new_n595), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G169), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n597), .A2(G179), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n586), .A2(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n564), .A2(new_n608), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n410), .A2(new_n523), .A3(new_n609), .ZN(G372));
  INV_X1    g0410(.A(KEYINPUT26), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT90), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n600), .B2(new_n607), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n578), .A2(KEYINPUT80), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(new_n585), .A3(new_n243), .ZN(new_n615));
  INV_X1    g0415(.A(new_n566), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n603), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n605), .A2(new_n606), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n586), .A2(new_n598), .A3(new_n599), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(KEYINPUT90), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n613), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n611), .B1(new_n560), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT91), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n560), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(KEYINPUT26), .A3(new_n608), .ZN(new_n627));
  OAI211_X1 g0427(.A(KEYINPUT91), .B(new_n611), .C1(new_n560), .C2(new_n622), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n619), .A2(KEYINPUT90), .A3(new_n620), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT90), .B1(new_n619), .B2(new_n620), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n560), .A2(new_n563), .A3(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n447), .A2(new_n451), .A3(KEYINPUT89), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n285), .B1(new_n449), .B2(new_n420), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n445), .B1(new_n635), .B2(KEYINPUT88), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n456), .B1(new_n636), .B2(new_n455), .ZN(new_n637));
  OAI21_X1  g0437(.A(G169), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n481), .B1(new_n638), .B2(new_n487), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n633), .B(new_n482), .C1(new_n639), .C2(new_n516), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n629), .A2(new_n640), .A3(new_n619), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n409), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n349), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n407), .A2(new_n367), .A3(new_n364), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(new_n404), .ZN(new_n645));
  INV_X1    g0445(.A(new_n341), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n293), .B(new_n294), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n642), .A2(new_n297), .A3(new_n647), .ZN(G369));
  NAND2_X1  g0448(.A1(new_n465), .A2(new_n204), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n511), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n516), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n516), .A2(new_n521), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n656), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n482), .B(new_n489), .C1(new_n481), .C2(new_n655), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n489), .B2(new_n655), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n482), .A2(new_n489), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n654), .B1(new_n510), .B2(new_n515), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n654), .B(KEYINPUT92), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n639), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n207), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n203), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n572), .A2(G116), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n674), .A2(new_n675), .B1(new_n211), .B2(new_n673), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n676), .B(KEYINPUT28), .Z(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT26), .B1(new_n560), .B2(new_n622), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n542), .A2(new_n555), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n531), .A2(new_n541), .A3(new_n561), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n295), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n679), .A2(new_n681), .A3(new_n611), .A4(new_n608), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n607), .B(KEYINPUT95), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT96), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT96), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n678), .A2(new_n686), .A3(new_n682), .A4(new_n683), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n685), .A2(new_n640), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(KEYINPUT29), .A3(new_n655), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n641), .A2(new_n668), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(KEYINPUT29), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n667), .A2(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n512), .A2(KEYINPUT93), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n443), .A2(G270), .A3(new_n285), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n556), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT93), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(G179), .A4(new_n494), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n597), .A2(new_n444), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n694), .A2(new_n698), .A3(new_n453), .A4(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(new_n702), .A3(new_n559), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT30), .B1(new_n680), .B2(new_n700), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n459), .A2(new_n334), .A3(new_n496), .A4(new_n604), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n559), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n693), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n707), .B1(new_n703), .B2(new_n704), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n655), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n564), .A2(new_n608), .A3(new_n668), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n710), .B(new_n713), .C1(new_n523), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT94), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(KEYINPUT94), .A3(G330), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n692), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n677), .B1(new_n721), .B2(G1), .ZN(G364));
  NOR2_X1   g0522(.A1(new_n464), .A2(G20), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT97), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G45), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n674), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n660), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G330), .B2(new_n659), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n207), .A2(new_n273), .ZN(new_n730));
  INV_X1    g0530(.A(G355), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n730), .A2(new_n731), .B1(G116), .B2(new_n207), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n235), .A2(new_n429), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n207), .A2(new_n282), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n211), .B2(new_n263), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n732), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n212), .B1(G20), .B2(new_n295), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n727), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n204), .A2(new_n287), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(new_n334), .A3(G200), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT98), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G303), .ZN(new_n751));
  NAND3_X1  g0551(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n753), .A2(KEYINPUT99), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(KEYINPUT99), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(KEYINPUT33), .B(G317), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n204), .B1(new_n759), .B2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n204), .A2(G190), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(new_n334), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(G283), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n282), .B1(new_n760), .B2(new_n761), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n752), .A2(new_n287), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(G326), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n334), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n744), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G322), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n762), .A2(new_n759), .ZN(new_n771));
  INV_X1    g0571(.A(G329), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n762), .A2(new_n768), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n773), .B1(G311), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n751), .A2(new_n758), .A3(new_n767), .A4(new_n776), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n352), .A2(new_n763), .B1(new_n769), .B2(new_n319), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n282), .B(new_n778), .C1(G77), .C2(new_n775), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n750), .A2(G87), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n771), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT32), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n782), .A2(new_n783), .B1(G50), .B2(new_n766), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n760), .A2(new_n498), .ZN(new_n785));
  INV_X1    g0585(.A(new_n782), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(new_n786), .B2(KEYINPUT32), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n779), .A2(new_n780), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n756), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n257), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n777), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT100), .ZN(new_n792));
  INV_X1    g0592(.A(new_n740), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n791), .B2(KEYINPUT100), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n743), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n739), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n659), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n729), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(G396));
  INV_X1    g0599(.A(new_n720), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n363), .A2(new_n654), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n368), .A2(new_n370), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n368), .B2(new_n801), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n667), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n641), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n690), .B2(new_n803), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n800), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n727), .B1(new_n800), .B2(new_n807), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n804), .A2(new_n737), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n793), .A2(new_n738), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n727), .B1(G77), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n750), .A2(G107), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n282), .B1(new_n763), .B2(new_n571), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n785), .B(new_n815), .C1(G303), .C2(new_n766), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n756), .A2(G283), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n769), .A2(new_n761), .B1(new_n771), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G116), .B2(new_n775), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n814), .A2(new_n816), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n769), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G143), .A2(new_n822), .B1(new_n775), .B2(G159), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  INV_X1    g0624(.A(new_n766), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n824), .B2(new_n825), .C1(new_n789), .C2(new_n252), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(KEYINPUT101), .B(KEYINPUT34), .Z(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n763), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n282), .B1(new_n830), .B2(G68), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n319), .B2(new_n760), .C1(new_n832), .C2(new_n771), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G50), .B2(new_n750), .ZN(new_n834));
  INV_X1    g0634(.A(new_n828), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n826), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n821), .B1(new_n829), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n813), .B1(new_n837), .B2(new_n740), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G384));
  OR2_X1    g0640(.A1(new_n548), .A2(KEYINPUT35), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n548), .A2(KEYINPUT35), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n841), .A2(G116), .A3(new_n213), .A4(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT36), .Z(new_n844));
  OAI211_X1 g0644(.A(new_n211), .B(G77), .C1(new_n319), .C2(new_n257), .ZN(new_n845));
  INV_X1    g0645(.A(G50), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(G68), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n203), .B(G13), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n647), .A2(new_n297), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n692), .B2(new_n409), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n368), .A2(new_n654), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n806), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n347), .A2(new_n337), .A3(new_n340), .A4(new_n348), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n652), .B1(new_n330), .B2(new_n332), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n857), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n345), .A2(new_n336), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n857), .B2(KEYINPUT102), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n861), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n857), .B1(new_n338), .B2(new_n335), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n345), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n855), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n856), .A2(new_n857), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n862), .A4(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n406), .A2(new_n655), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n404), .A2(new_n407), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n404), .B2(new_n407), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n854), .A2(new_n870), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n646), .A2(new_n652), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n404), .A2(new_n654), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n869), .ZN(new_n881));
  INV_X1    g0681(.A(new_n869), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n860), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT37), .B1(new_n864), .B2(new_n345), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT103), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n860), .A2(new_n883), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT103), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n864), .A2(KEYINPUT37), .A3(new_n345), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n886), .A2(new_n868), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n882), .B1(new_n855), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n880), .B(new_n881), .C1(new_n892), .C2(KEYINPUT39), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n877), .A2(new_n878), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n851), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n891), .A2(new_n855), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n869), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n803), .B1(new_n873), .B2(new_n874), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AND4_X1   g0699(.A1(new_n608), .A2(new_n560), .A3(new_n563), .A4(new_n668), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n900), .A2(new_n489), .A3(new_n482), .A4(new_n522), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n702), .B1(new_n701), .B2(new_n559), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n680), .A2(new_n700), .A3(KEYINPUT30), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n708), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n901), .A2(new_n713), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n897), .A2(new_n899), .A3(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n905), .A2(new_n713), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n898), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT40), .B1(new_n867), .B2(new_n869), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n907), .A2(KEYINPUT40), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n906), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n911), .B1(new_n410), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n909), .B2(new_n897), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n909), .A2(new_n910), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n409), .B(new_n906), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(new_n917), .A3(G330), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n895), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n203), .B2(new_n724), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n895), .A2(new_n918), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n849), .B1(new_n920), .B2(new_n921), .ZN(G367));
  NAND2_X1  g0722(.A1(new_n626), .A2(new_n667), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n560), .B(new_n563), .C1(new_n554), .C2(new_n668), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n664), .A2(new_n925), .A3(new_n665), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n639), .A2(new_n563), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n667), .B1(new_n928), .B2(new_n560), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n926), .B2(KEYINPUT42), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT105), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT105), .B1(new_n933), .B2(new_n929), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n586), .A2(new_n599), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n619), .A2(new_n936), .A3(new_n655), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n655), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n937), .B1(new_n622), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT104), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT104), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n935), .A2(new_n944), .A3(new_n940), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n943), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n944), .B1(new_n935), .B2(new_n940), .ZN(new_n948));
  INV_X1    g0748(.A(new_n940), .ZN(new_n949));
  AOI211_X1 g0749(.A(KEYINPUT104), .B(new_n949), .C1(new_n932), .C2(new_n934), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n947), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n925), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n663), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n946), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT106), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n725), .A2(G1), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n721), .ZN(new_n960));
  INV_X1    g0760(.A(new_n663), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n666), .A2(new_n669), .A3(new_n925), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n666), .A2(KEYINPUT45), .A3(new_n669), .A4(new_n925), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT44), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n670), .B2(new_n925), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n666), .A2(new_n669), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(KEYINPUT44), .A3(new_n952), .ZN(new_n969));
  AOI221_X4 g0769(.A(new_n961), .B1(new_n964), .B2(new_n965), .C1(new_n967), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n964), .A2(new_n965), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n663), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n666), .B1(new_n662), .B2(new_n665), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n660), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n960), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n673), .B(KEYINPUT41), .Z(new_n978));
  OAI21_X1  g0778(.A(new_n959), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n946), .A2(new_n951), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n953), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n946), .A2(new_n951), .A3(KEYINPUT106), .A4(new_n954), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n957), .A2(new_n979), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n741), .B1(new_n207), .B2(new_n359), .C1(new_n230), .C2(new_n734), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n727), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n750), .A2(G58), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n756), .A2(G159), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n760), .A2(new_n257), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n273), .B1(new_n769), .B2(new_n252), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G143), .C2(new_n766), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n763), .A2(new_n276), .B1(new_n771), .B2(new_n824), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G50), .B2(new_n775), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n986), .A2(new_n987), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n750), .A2(KEYINPUT46), .A3(G116), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT46), .ZN(new_n995));
  INV_X1    g0795(.A(G116), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n995), .B1(new_n749), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n994), .B(new_n997), .C1(new_n761), .C2(new_n789), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n825), .A2(new_n818), .ZN(new_n999));
  INV_X1    g0799(.A(new_n771), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n273), .B(new_n999), .C1(G317), .C2(new_n1000), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n763), .A2(new_n498), .B1(new_n774), .B2(new_n764), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G303), .B2(new_n822), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1001), .B(new_n1003), .C1(new_n352), .C2(new_n760), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n993), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT47), .Z(new_n1006));
  OAI221_X1 g0806(.A(new_n985), .B1(new_n939), .B2(new_n796), .C1(new_n793), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n983), .A2(new_n1007), .ZN(G387));
  NAND2_X1  g0808(.A1(new_n721), .A2(new_n976), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n673), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n721), .A2(new_n976), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n227), .A2(new_n263), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1013), .A2(new_n734), .B1(new_n675), .B2(new_n730), .ZN(new_n1014));
  AOI21_X1  g0814(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n250), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1016), .A2(KEYINPUT50), .A3(new_n846), .ZN(new_n1017));
  AOI21_X1  g0817(.A(KEYINPUT50), .B1(new_n1016), .B2(new_n846), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n675), .B(new_n1015), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1014), .A2(new_n1019), .B1(new_n352), .B2(new_n672), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n727), .B1(new_n1020), .B2(new_n742), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n756), .A2(new_n1016), .B1(G68), .B2(new_n775), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT107), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n749), .A2(new_n276), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G50), .A2(new_n822), .B1(new_n1000), .B2(G150), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1025), .B(new_n273), .C1(new_n498), .C2(new_n763), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n825), .A2(new_n781), .B1(new_n760), .B2(new_n359), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT108), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G317), .A2(new_n822), .B1(new_n775), .B2(G303), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n770), .B2(new_n825), .C1(new_n789), .C2(new_n818), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT109), .Z(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT48), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(KEYINPUT48), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n760), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n750), .A2(G294), .B1(G283), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT49), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT110), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n763), .A2(new_n996), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n273), .B(new_n1042), .C1(G326), .C2(new_n1000), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1029), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1021), .B1(new_n1045), .B2(new_n740), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT111), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n662), .A2(new_n796), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1048), .A2(new_n1049), .B1(new_n958), .B2(new_n976), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1012), .A2(new_n1050), .ZN(G393));
  NAND2_X1  g0851(.A1(new_n971), .A2(new_n972), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n961), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT112), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n971), .A2(new_n663), .A3(new_n972), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n970), .B1(new_n973), .B2(KEYINPUT112), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n1009), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n974), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1058), .B(new_n673), .C1(new_n1009), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n952), .A2(new_n739), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n741), .B1(new_n498), .B2(new_n207), .C1(new_n238), .C2(new_n734), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n727), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n282), .B1(new_n763), .B2(new_n352), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n774), .A2(new_n761), .B1(new_n771), .B2(new_n770), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G116), .C2(new_n1035), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n764), .B2(new_n749), .C1(new_n492), .C2(new_n789), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n822), .A2(G311), .B1(G317), .B2(new_n766), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT52), .ZN(new_n1070));
  INV_X1    g0870(.A(G143), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n774), .A2(new_n250), .B1(new_n771), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n273), .B1(new_n763), .B2(new_n571), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n760), .A2(new_n276), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n257), .B2(new_n749), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n825), .A2(new_n252), .B1(new_n769), .B2(new_n781), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1078));
  XNOR2_X1  g0878(.A(new_n1077), .B(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n789), .B2(new_n846), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1068), .A2(new_n1070), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1064), .B1(new_n1081), .B2(new_n740), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1061), .A2(new_n958), .B1(new_n1062), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1060), .A2(new_n1083), .ZN(G390));
  NAND3_X1  g0884(.A1(new_n688), .A2(new_n655), .A3(new_n803), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT114), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n1085), .A2(new_n1086), .A3(new_n853), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n1085), .B2(new_n853), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(G330), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n904), .A2(new_n654), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n709), .B1(new_n1091), .B2(new_n711), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n717), .B(new_n1090), .C1(new_n1092), .C2(new_n901), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT94), .B1(new_n715), .B2(G330), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n899), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n906), .A2(G330), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n875), .B1(new_n1096), .B2(new_n804), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(KEYINPUT116), .B1(new_n1089), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1090), .B1(new_n908), .B2(new_n901), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n876), .B1(new_n1100), .B2(new_n803), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n720), .B2(new_n899), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1085), .A2(new_n853), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(KEYINPUT114), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1085), .A2(new_n1086), .A3(new_n853), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT116), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1102), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n803), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n875), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1096), .A2(new_n898), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1099), .A2(new_n1108), .B1(new_n854), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n409), .A2(new_n1100), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n851), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1104), .A2(new_n876), .A3(new_n1105), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n892), .A2(new_n880), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n852), .B1(new_n641), .B2(new_n805), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n879), .B1(new_n1120), .B2(new_n875), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT115), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n869), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT39), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n897), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT115), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1127), .B(new_n879), .C1(new_n1120), .C2(new_n875), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1122), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1119), .A2(new_n1095), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1112), .B1(new_n1119), .B2(new_n1129), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1114), .A2(new_n1116), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1113), .A2(new_n854), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1089), .A2(new_n1098), .A3(KEYINPUT116), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1107), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1119), .A2(new_n1129), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1111), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1119), .A2(new_n1095), .A3(new_n1129), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1116), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1132), .A2(new_n1141), .A3(new_n673), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1126), .A2(new_n737), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n727), .B1(new_n1016), .B2(new_n812), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n282), .B1(new_n763), .B2(new_n257), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1074), .B(new_n1145), .C1(G283), .C2(new_n766), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n756), .A2(G107), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n769), .A2(new_n996), .B1(new_n774), .B2(new_n498), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G294), .B2(new_n1000), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n780), .A2(new_n1146), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n750), .A2(G150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT53), .ZN(new_n1152));
  INV_X1    g0952(.A(G128), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n825), .A2(new_n1153), .B1(new_n760), .B2(new_n781), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n273), .B1(new_n769), .B2(new_n832), .ZN(new_n1155));
  INV_X1    g0955(.A(G125), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n763), .A2(new_n846), .B1(new_n771), .B2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT117), .Z(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1158), .B1(new_n1161), .B2(new_n774), .C1(new_n824), .C2(new_n789), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1150), .B1(new_n1152), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1144), .B1(new_n1163), .B2(new_n740), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT118), .Z(new_n1165));
  NAND2_X1  g0965(.A1(new_n1143), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1125), .B1(new_n1121), .B2(KEYINPUT115), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1117), .A2(new_n1118), .B1(new_n1167), .B2(new_n1128), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1139), .B1(new_n1168), .B2(new_n1112), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1166), .B1(new_n1169), .B2(new_n959), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1142), .A2(new_n1171), .ZN(G378));
  NOR2_X1   g0972(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1116), .B1(new_n1173), .B2(new_n1136), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1175));
  NAND2_X1  g0975(.A1(new_n298), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n652), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n260), .A2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT119), .Z(new_n1179));
  INV_X1    g0979(.A(new_n1175), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n293), .A2(new_n294), .A3(new_n297), .A4(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1176), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1179), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n911), .B2(new_n1090), .ZN(new_n1186));
  OAI211_X1 g0986(.A(G330), .B(new_n1184), .C1(new_n916), .C2(new_n915), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1186), .A2(new_n894), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n894), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT57), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n673), .B1(new_n1174), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1186), .A2(new_n894), .A3(new_n1187), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(KEYINPUT120), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(KEYINPUT120), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1140), .B1(new_n1169), .B2(new_n1114), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1192), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n273), .A2(G41), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G50), .B(new_n1200), .C1(new_n278), .C2(new_n264), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n763), .A2(new_n319), .B1(new_n771), .B2(new_n764), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1202), .B(new_n1024), .C1(new_n565), .C2(new_n775), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1200), .B1(new_n352), .B2(new_n769), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n988), .B(new_n1204), .C1(G116), .C2(new_n766), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(new_n498), .C2(new_n789), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT58), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1201), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n760), .A2(new_n252), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n769), .A2(new_n1153), .B1(new_n774), .B2(new_n824), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G125), .C2(new_n766), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n749), .B2(new_n1161), .C1(new_n789), .C2(new_n832), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n278), .B(new_n264), .C1(new_n763), .C2(new_n781), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G124), .B2(new_n1000), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1208), .B1(new_n1207), .B2(new_n1206), .C1(new_n1213), .C2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n740), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n727), .C1(G50), .C2(new_n812), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1185), .B2(new_n737), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1196), .B2(new_n958), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1199), .A2(new_n1222), .ZN(G375));
  NAND2_X1  g1023(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n978), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n875), .A2(new_n737), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n727), .B1(G68), .B2(new_n812), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n749), .A2(new_n498), .B1(new_n492), .B2(new_n771), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT121), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n789), .A2(new_n996), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G283), .A2(new_n822), .B1(new_n775), .B2(G107), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1233), .B(new_n282), .C1(new_n276), .C2(new_n763), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n825), .A2(new_n761), .B1(new_n760), .B2(new_n359), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1231), .A2(new_n1232), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1236), .A2(KEYINPUT122), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(KEYINPUT122), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n750), .A2(G159), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n273), .B1(new_n763), .B2(new_n319), .C1(new_n832), .C2(new_n825), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G50), .B2(new_n1035), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n756), .A2(new_n1160), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n769), .A2(new_n824), .B1(new_n771), .B2(new_n1153), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G150), .B2(new_n775), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .A4(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1237), .A2(new_n1238), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1229), .B1(new_n1246), .B2(new_n740), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1136), .A2(new_n958), .B1(new_n1228), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1227), .A2(new_n1248), .ZN(G381));
  INV_X1    g1049(.A(G390), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1012), .A2(new_n798), .A3(new_n1050), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1252), .A3(new_n839), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1253), .A2(G387), .A3(G381), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n673), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1224), .B2(new_n1169), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1170), .B1(new_n1256), .B2(new_n1141), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1257), .A3(new_n1199), .A4(new_n1222), .ZN(G407));
  NAND3_X1  g1058(.A1(new_n1257), .A2(G213), .A3(new_n653), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G407), .B(G213), .C1(G375), .C2(new_n1259), .ZN(G409));
  NAND3_X1  g1060(.A1(new_n983), .A2(new_n1007), .A3(G390), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT126), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1250), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT126), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n983), .A2(new_n1264), .A3(G390), .A4(new_n1007), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n798), .B1(new_n1012), .B2(new_n1050), .ZN(new_n1268));
  OR3_X1    g1068(.A1(new_n1252), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n1252), .B2(new_n1268), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1266), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT127), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1263), .B(new_n1261), .C1(new_n1252), .C2(new_n1268), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G378), .B(new_n1222), .C1(new_n1192), .C2(new_n1198), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1196), .A2(new_n1197), .A3(new_n1226), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1221), .B1(new_n1190), .B2(new_n958), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1257), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n653), .A2(G213), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1099), .A2(new_n1108), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1285), .A2(KEYINPUT60), .A3(new_n1116), .A4(new_n1133), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n673), .ZN(new_n1287));
  OAI21_X1  g1087(.A(KEYINPUT60), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1225), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1248), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1289), .A2(new_n839), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1225), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1286), .A2(new_n673), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G384), .B1(new_n1294), .B2(new_n1248), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1283), .A2(new_n1284), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT123), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1283), .A2(KEYINPUT123), .A3(new_n1296), .A4(new_n1284), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT62), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n839), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1294), .A2(G384), .A3(new_n1248), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n653), .A2(G213), .A3(G2897), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1303), .A2(new_n1304), .A3(new_n1306), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT124), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1303), .A2(new_n1304), .A3(KEYINPUT124), .A4(new_n1306), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1302), .A2(new_n1308), .A3(new_n1311), .A4(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1297), .A2(KEYINPUT62), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1277), .B1(new_n1301), .B2(new_n1316), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1283), .A2(new_n1284), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT61), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1299), .A2(new_n1321), .A3(new_n1300), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1323));
  OR2_X1    g1123(.A1(new_n1297), .A2(new_n1321), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1320), .A2(new_n1322), .A3(new_n1323), .A4(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1317), .A2(new_n1325), .ZN(G405));
  NAND2_X1  g1126(.A1(G375), .A2(new_n1257), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1278), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1296), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1323), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1327), .A2(new_n1278), .A3(new_n1305), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1329), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1330), .B1(new_n1329), .B2(new_n1331), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(G402));
endmodule


