//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(G478), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT15), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G128), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(KEYINPUT13), .A3(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n196), .B(G134), .C1(KEYINPUT13), .C2(new_n193), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n198), .A3(new_n195), .ZN(new_n199));
  INV_X1    g013(.A(G116), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G122), .ZN(new_n201));
  INV_X1    g015(.A(G122), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G116), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT90), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT90), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n203), .A3(new_n206), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n205), .A2(G107), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(G107), .B1(new_n205), .B2(new_n207), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n197), .B(new_n199), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT9), .B(G234), .ZN(new_n211));
  INV_X1    g025(.A(G217), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n211), .A2(new_n212), .A3(G953), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT14), .B1(new_n202), .B2(G116), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT91), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n201), .A2(KEYINPUT91), .A3(KEYINPUT14), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n203), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT14), .ZN(new_n220));
  INV_X1    g034(.A(new_n201), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n219), .A2(KEYINPUT92), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT92), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n217), .A2(new_n218), .A3(new_n223), .A4(new_n203), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n214), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n193), .A2(new_n195), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G134), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n199), .ZN(new_n228));
  INV_X1    g042(.A(new_n209), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n210), .B(new_n213), .C1(new_n225), .C2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT93), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n219), .A2(KEYINPUT92), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n221), .A2(new_n220), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n224), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G107), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n209), .B1(new_n227), .B2(new_n199), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(KEYINPUT93), .A3(new_n210), .A4(new_n213), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n210), .B1(new_n225), .B2(new_n230), .ZN(new_n241));
  INV_X1    g055(.A(new_n213), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n233), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G902), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT94), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT94), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(new_n248), .A3(new_n245), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n188), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n188), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(G214), .B1(G237), .B2(G902), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(G116), .B(G119), .Z(new_n256));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT2), .B(G113), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT2), .B(G113), .Z(new_n260));
  XNOR2_X1  g074(.A(G116), .B(G119), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT67), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI22_X1  g076(.A1(new_n259), .A2(new_n262), .B1(new_n261), .B2(new_n260), .ZN(new_n263));
  INV_X1    g077(.A(G104), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G107), .ZN(new_n265));
  OR2_X1    g079(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n214), .A2(G104), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n264), .A2(G107), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G101), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n266), .B1(new_n267), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G101), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n269), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n265), .A4(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(KEYINPUT4), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT4), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n280), .B(G101), .C1(new_n268), .C2(new_n272), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n263), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n276), .B1(new_n267), .B2(new_n265), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n268), .A2(new_n272), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(new_n276), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n257), .B1(new_n256), .B2(new_n258), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n289));
  INV_X1    g103(.A(G119), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(G116), .ZN(new_n291));
  OAI211_X1 g105(.A(G113), .B(new_n291), .C1(new_n256), .C2(new_n289), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n285), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n282), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(G110), .B(G122), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n282), .A2(new_n293), .A3(new_n295), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(KEYINPUT6), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT0), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT64), .B1(new_n300), .B2(new_n194), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT64), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT0), .A3(G128), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n194), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G146), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G143), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT65), .B(G143), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(G146), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n190), .A2(new_n192), .A3(G146), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(G143), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n312), .A2(KEYINPUT0), .A3(G128), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n194), .B1(new_n313), .B2(KEYINPUT1), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n312), .A2(new_n313), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G224), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(G953), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n324), .B(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n295), .B1(new_n282), .B2(new_n293), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT6), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n328), .A2(KEYINPUT81), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT81), .B1(new_n328), .B2(new_n329), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n299), .B(new_n327), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n295), .B(KEYINPUT8), .ZN(new_n333));
  INV_X1    g147(.A(new_n283), .ZN(new_n334));
  AND4_X1   g148(.A1(new_n288), .A2(new_n278), .A3(new_n334), .A4(new_n292), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n288), .A2(new_n292), .B1(new_n278), .B2(new_n334), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n333), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT83), .B1(new_n325), .B2(G953), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT7), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n326), .B2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n316), .A2(new_n323), .A3(new_n338), .A4(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n337), .A2(new_n298), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n316), .A2(KEYINPUT82), .A3(new_n323), .ZN(new_n344));
  OAI221_X1 g158(.A(new_n344), .B1(KEYINPUT82), .B2(new_n323), .C1(new_n339), .C2(new_n326), .ZN(new_n345));
  AOI21_X1  g159(.A(G902), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n332), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G210), .B1(G237), .B2(G902), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n332), .A2(new_n348), .A3(new_n346), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n255), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G475), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  INV_X1    g168(.A(G953), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G214), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n190), .A3(new_n192), .ZN(new_n357));
  INV_X1    g171(.A(G131), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n354), .A2(new_n355), .A3(G143), .A4(G214), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n357), .B2(new_n359), .ZN(new_n361));
  OR3_X1    g175(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT17), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n190), .A2(new_n192), .ZN(new_n363));
  INV_X1    g177(.A(G214), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n364), .A2(G237), .A3(G953), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n359), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT17), .A3(G131), .ZN(new_n367));
  INV_X1    g181(.A(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G125), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n320), .A2(G140), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT16), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n320), .A2(G140), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT16), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n306), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n371), .A2(new_n374), .A3(G146), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n367), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AND4_X1   g192(.A1(G143), .A2(new_n354), .A3(new_n355), .A4(G214), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n309), .B2(new_n356), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT18), .A2(G131), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT84), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT84), .ZN(new_n383));
  INV_X1    g197(.A(new_n381), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n366), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n369), .A2(new_n370), .A3(new_n306), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n368), .A2(G125), .ZN(new_n388));
  OAI21_X1  g202(.A(G146), .B1(new_n372), .B2(new_n388), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n380), .A2(new_n381), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n362), .A2(new_n378), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(G113), .B(G122), .Z(new_n392));
  XOR2_X1   g206(.A(KEYINPUT86), .B(G104), .Z(new_n393));
  XOR2_X1   g207(.A(new_n392), .B(new_n393), .Z(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n391), .B(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n353), .B1(new_n396), .B2(new_n245), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT19), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT19), .B1(new_n369), .B2(new_n370), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n306), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT85), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT19), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n372), .B2(new_n388), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT19), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n306), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n371), .A2(G146), .A3(new_n374), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n366), .A2(G131), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n386), .A2(new_n390), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT87), .B1(new_n413), .B2(new_n395), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n362), .A2(new_n378), .ZN(new_n415));
  INV_X1    g229(.A(new_n385), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n383), .B1(new_n366), .B2(new_n384), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n390), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n395), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n377), .B1(new_n360), .B2(new_n361), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n407), .B2(new_n401), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n389), .A2(new_n387), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n366), .B2(new_n384), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n382), .B2(new_n385), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n420), .B(new_n394), .C1(new_n422), .C2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n414), .A2(new_n419), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G475), .A2(G902), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT88), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n410), .A2(new_n411), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n406), .B1(new_n405), .B2(new_n306), .ZN(new_n432));
  AOI211_X1 g246(.A(KEYINPUT85), .B(G146), .C1(new_n403), .C2(new_n404), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n377), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n395), .B1(new_n434), .B2(new_n418), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n420), .A2(new_n435), .B1(new_n391), .B2(new_n395), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT89), .B1(new_n436), .B2(new_n414), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n430), .B1(new_n437), .B2(KEYINPUT20), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n427), .A2(KEYINPUT89), .A3(new_n439), .A4(new_n429), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n397), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n355), .A2(G952), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(G234), .B2(G237), .ZN(new_n443));
  NAND2_X1  g257(.A1(G234), .A2(G237), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(G902), .A3(G953), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(G898), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AND4_X1   g263(.A1(new_n253), .A2(new_n352), .A3(new_n441), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(G217), .A2(G902), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n212), .B2(G234), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n452), .B(KEYINPUT71), .Z(new_n453));
  NAND3_X1  g267(.A1(new_n355), .A2(G221), .A3(G234), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT74), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT22), .B(G137), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT23), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n290), .B2(G128), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n290), .A2(G128), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G119), .B(G128), .ZN(new_n464));
  INV_X1    g278(.A(G110), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT24), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT24), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G110), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n463), .A2(G110), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(G146), .B1(new_n371), .B2(new_n374), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n409), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT72), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n470), .B(KEYINPUT72), .C1(new_n409), .C2(new_n471), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT73), .ZN(new_n477));
  OAI22_X1  g291(.A1(new_n463), .A2(G110), .B1(new_n464), .B2(new_n469), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n377), .A3(new_n387), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n477), .B1(new_n476), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n458), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n376), .A2(new_n377), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT72), .B1(new_n483), .B2(new_n470), .ZN(new_n484));
  INV_X1    g298(.A(new_n475), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n479), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n457), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT25), .B1(new_n488), .B2(new_n245), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT25), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n490), .B(G902), .C1(new_n482), .C2(new_n487), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n453), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n453), .A2(G902), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n493), .B(KEYINPUT75), .Z(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G472), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n245), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT11), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n198), .B2(G137), .ZN(new_n500));
  INV_X1    g314(.A(G137), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(KEYINPUT11), .A3(G134), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n198), .A2(G137), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(KEYINPUT66), .A2(G131), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n500), .A2(new_n502), .A3(new_n505), .A4(new_n503), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n311), .A3(new_n314), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n500), .A2(new_n502), .A3(new_n358), .A4(new_n503), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n198), .A2(G137), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n501), .A2(G134), .ZN(new_n513));
  OAI21_X1  g327(.A(G131), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n191), .A2(G143), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n306), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n317), .B1(new_n518), .B2(new_n308), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n312), .A2(new_n313), .A3(new_n321), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n510), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n510), .B2(new_n521), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n263), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n286), .A2(new_n287), .B1(new_n256), .B2(new_n258), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n510), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n354), .A2(new_n355), .A3(G210), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT27), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT26), .B(G101), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n525), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n525), .A2(KEYINPUT31), .A3(new_n527), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n510), .A2(new_n521), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n263), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n527), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT28), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(KEYINPUT68), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT68), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n510), .A2(new_n521), .A3(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n541), .A2(new_n526), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n540), .B1(new_n544), .B2(KEYINPUT28), .ZN(new_n545));
  INV_X1    g359(.A(new_n531), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n498), .B1(new_n536), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n263), .B1(new_n537), .B2(KEYINPUT68), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT28), .B1(new_n549), .B2(new_n543), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n527), .A2(KEYINPUT70), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT70), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n510), .A2(new_n521), .A3(new_n553), .A4(new_n526), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n538), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT28), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n551), .A2(new_n556), .A3(KEYINPUT29), .A4(new_n531), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT29), .ZN(new_n558));
  INV_X1    g372(.A(new_n527), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n537), .A2(KEYINPUT30), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n510), .A2(new_n521), .A3(new_n522), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n559), .B1(new_n562), .B2(new_n263), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n558), .B1(new_n563), .B2(new_n531), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT28), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(new_n538), .B2(new_n527), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n550), .A2(new_n566), .A3(new_n546), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n557), .B(new_n245), .C1(new_n564), .C2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(KEYINPUT32), .A2(new_n548), .B1(new_n568), .B2(G472), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT69), .B(KEYINPUT32), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n534), .A2(new_n535), .B1(new_n545), .B2(new_n546), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n571), .B2(new_n498), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n496), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(G221), .B1(new_n211), .B2(G902), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n278), .A2(new_n334), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n312), .A2(new_n313), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT1), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n363), .B2(new_n306), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n577), .B1(new_n579), .B2(new_n194), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n576), .B1(new_n322), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT78), .B1(new_n581), .B2(KEYINPUT10), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT1), .B1(new_n309), .B2(G146), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n583), .A2(G128), .B1(new_n313), .B2(new_n312), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n285), .B1(new_n520), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT78), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n281), .A2(new_n311), .A3(new_n314), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n587), .B1(new_n319), .B2(new_n322), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n589), .A2(new_n279), .B1(new_n590), .B2(new_n285), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n582), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n509), .ZN(new_n593));
  INV_X1    g407(.A(new_n509), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n582), .A2(new_n588), .A3(new_n591), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(G110), .B(G140), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n355), .A2(G227), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT79), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n307), .B1(new_n363), .B2(new_n306), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n322), .B1(new_n602), .B2(new_n317), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n285), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n576), .A2(KEYINPUT79), .A3(new_n319), .A4(new_n322), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n585), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n509), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT12), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n606), .A2(KEYINPUT12), .A3(new_n509), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n599), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n595), .A2(KEYINPUT80), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT80), .B1(new_n595), .B2(new_n612), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n600), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G469), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n245), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n245), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n606), .A2(KEYINPUT12), .A3(new_n509), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT12), .B1(new_n606), .B2(new_n509), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n595), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n599), .B(KEYINPUT76), .Z(new_n623));
  AND2_X1   g437(.A1(new_n595), .A2(new_n612), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n622), .A2(new_n623), .B1(new_n624), .B2(new_n593), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n619), .B1(new_n625), .B2(G469), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n575), .B1(new_n618), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n450), .A2(new_n573), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  OAI21_X1  g443(.A(G472), .B1(new_n571), .B2(G902), .ZN(new_n630));
  INV_X1    g444(.A(new_n548), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n492), .A2(new_n495), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n627), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n352), .A2(new_n449), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n241), .B2(new_n242), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n244), .A2(new_n638), .B1(new_n231), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n187), .A2(G902), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n640), .A2(new_n641), .B1(new_n187), .B2(new_n246), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT95), .B1(new_n441), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n396), .A2(new_n245), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G475), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT89), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n426), .A2(new_n419), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n435), .A2(new_n420), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n649), .A2(new_n439), .B1(new_n427), .B2(new_n429), .ZN(new_n650));
  AND4_X1   g464(.A1(KEYINPUT89), .A2(new_n427), .A3(new_n439), .A4(new_n429), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n645), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT95), .ZN(new_n653));
  INV_X1    g467(.A(new_n642), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n643), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n635), .A2(new_n637), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT34), .B(G104), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  XNOR2_X1  g473(.A(new_n448), .B(KEYINPUT96), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n332), .A2(new_n348), .A3(new_n346), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n348), .B1(new_n332), .B2(new_n346), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n254), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n427), .A2(new_n439), .A3(new_n429), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n439), .B1(new_n427), .B2(new_n429), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n645), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n188), .ZN(new_n668));
  INV_X1    g482(.A(new_n249), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n248), .B1(new_n244), .B2(new_n245), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n667), .B1(new_n671), .B2(new_n251), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT97), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n664), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n430), .A2(KEYINPUT20), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n427), .A2(new_n439), .A3(new_n429), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n397), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n250), .B2(new_n252), .ZN(new_n678));
  OAI21_X1  g492(.A(KEYINPUT97), .B1(new_n678), .B2(new_n663), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n635), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT35), .B(G107), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  INV_X1    g497(.A(new_n494), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n486), .A2(KEYINPUT73), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n687), .B1(KEYINPUT36), .B2(new_n458), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n458), .A2(KEYINPUT36), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n684), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n487), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n687), .B2(new_n458), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n490), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n488), .A2(KEYINPUT25), .A3(new_n245), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n691), .B1(new_n696), .B2(new_n453), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n632), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n450), .A2(new_n627), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  NAND2_X1  g515(.A1(new_n548), .A2(KEYINPUT32), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n568), .A2(G472), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n703), .A3(new_n572), .ZN(new_n704));
  INV_X1    g518(.A(new_n691), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n492), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n627), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n443), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n445), .A2(G900), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n667), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n671), .A2(new_n251), .ZN(new_n713));
  AND4_X1   g527(.A1(KEYINPUT98), .A2(new_n712), .A3(new_n352), .A4(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n707), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT98), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n712), .A2(new_n713), .ZN(new_n717));
  INV_X1    g531(.A(new_n352), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT99), .B(G128), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G30));
  XNOR2_X1  g536(.A(new_n710), .B(KEYINPUT39), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n627), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(KEYINPUT40), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n350), .A2(new_n351), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT38), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n563), .A2(new_n546), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n245), .B1(new_n555), .B2(new_n531), .ZN(new_n729));
  OAI21_X1  g543(.A(G472), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n702), .A2(new_n572), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n727), .A2(new_n254), .A3(new_n697), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n713), .A2(new_n652), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n725), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(KEYINPUT40), .B2(new_n724), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n363), .ZN(G45));
  AND4_X1   g550(.A1(new_n704), .A2(new_n627), .A3(new_n352), .A4(new_n706), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT100), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n438), .A2(new_n440), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n642), .B1(new_n739), .B2(new_n645), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n738), .B1(new_n740), .B2(new_n710), .ZN(new_n741));
  NOR4_X1   g555(.A1(new_n441), .A2(KEYINPUT100), .A3(new_n642), .A4(new_n711), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G146), .ZN(G48));
  AND3_X1   g559(.A1(new_n616), .A2(new_n617), .A3(new_n245), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n617), .B1(new_n616), .B2(new_n245), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n746), .A2(new_n747), .A3(new_n575), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n573), .A2(new_n656), .A3(new_n748), .A4(new_n637), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT41), .B(G113), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT101), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n749), .B(new_n751), .ZN(G15));
  INV_X1    g566(.A(KEYINPUT102), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n673), .B1(new_n664), .B2(new_n672), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n678), .A2(new_n663), .A3(KEYINPUT97), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n573), .A2(new_n748), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n680), .A2(KEYINPUT102), .A3(new_n573), .A4(new_n748), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  AOI21_X1  g575(.A(new_n697), .B1(new_n569), .B2(new_n572), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n713), .A2(new_n652), .A3(new_n448), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n748), .A3(new_n352), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G119), .ZN(G21));
  NOR2_X1   g579(.A1(new_n718), .A2(new_n733), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n551), .A2(new_n556), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n546), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n536), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n498), .B(KEYINPUT103), .Z(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n492), .A2(new_n630), .A3(new_n771), .A4(new_n495), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n766), .A2(new_n748), .A3(new_n773), .A4(new_n660), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  NAND2_X1  g589(.A1(new_n616), .A2(new_n245), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(G469), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n574), .A3(new_n618), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n718), .ZN(new_n779));
  AOI21_X1  g593(.A(G902), .B1(new_n536), .B2(new_n547), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n546), .A2(new_n767), .B1(new_n534), .B2(new_n535), .ZN(new_n781));
  INV_X1    g595(.A(new_n770), .ZN(new_n782));
  OAI22_X1  g596(.A1(new_n780), .A2(new_n497), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n697), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n743), .A2(KEYINPUT104), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT104), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n652), .A2(new_n654), .A3(new_n710), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT100), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n652), .A2(new_n654), .A3(new_n738), .A4(new_n710), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n746), .A2(new_n747), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n574), .A3(new_n352), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n786), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n785), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G125), .ZN(G27));
  NAND2_X1  g609(.A1(new_n622), .A2(new_n623), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT105), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n624), .A2(new_n593), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n622), .A2(KEYINPUT105), .A3(new_n623), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(G469), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n619), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n618), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n661), .A2(new_n662), .A3(new_n575), .A4(new_n255), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n634), .A2(new_n803), .A3(new_n704), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n743), .A2(new_n805), .A3(KEYINPUT106), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT42), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT106), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n788), .A2(new_n789), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n634), .A2(new_n803), .A3(new_n704), .A4(new_n804), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n806), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n569), .B1(KEYINPUT32), .B2(new_n548), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n634), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n807), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n743), .A3(new_n803), .A4(new_n804), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g631(.A(KEYINPUT107), .B(G131), .Z(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(G33));
  OR2_X1    g633(.A1(new_n810), .A2(new_n717), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G134), .ZN(G36));
  NOR2_X1   g635(.A1(new_n726), .A2(new_n255), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT43), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n652), .B2(KEYINPUT109), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n441), .A2(new_n654), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n826), .A2(new_n633), .A3(new_n697), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n822), .B1(new_n827), .B2(KEYINPUT44), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(KEYINPUT44), .B2(new_n827), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n625), .A2(KEYINPUT45), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n617), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n798), .A2(KEYINPUT45), .A3(new_n799), .A4(new_n800), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n619), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n746), .B1(new_n833), .B2(KEYINPUT46), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(KEYINPUT108), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n833), .A2(KEYINPUT46), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n834), .B2(KEYINPUT108), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n575), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n829), .A2(new_n723), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(G137), .ZN(G39));
  NOR2_X1   g655(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n839), .B1(new_n844), .B2(new_n842), .ZN(new_n845));
  INV_X1    g659(.A(new_n822), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n809), .A2(new_n634), .A3(new_n704), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n843), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(G140), .ZN(G42));
  NOR4_X1   g663(.A1(new_n496), .A2(new_n825), .A3(new_n575), .A4(new_n255), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT49), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n850), .B1(new_n851), .B2(new_n791), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT111), .Z(new_n853));
  AOI211_X1 g667(.A(new_n731), .B(new_n727), .C1(new_n851), .C2(new_n791), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n826), .A2(new_n708), .ZN(new_n856));
  INV_X1    g670(.A(new_n814), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n778), .A2(new_n846), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT48), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n731), .A2(new_n496), .A3(new_n708), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n858), .A2(new_n656), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n856), .A2(new_n773), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n779), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n442), .B(KEYINPUT116), .Z(new_n866));
  NAND4_X1  g680(.A1(new_n860), .A2(new_n862), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n863), .A2(KEYINPUT115), .A3(new_n846), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT115), .B1(new_n863), .B2(new_n846), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n845), .B1(new_n839), .B2(new_n842), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n791), .A2(new_n575), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n727), .A2(new_n778), .A3(new_n254), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n864), .A2(KEYINPUT50), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n876));
  INV_X1    g690(.A(new_n874), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n876), .B1(new_n863), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n856), .A2(new_n784), .A3(new_n858), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n858), .A2(new_n441), .A3(new_n642), .A4(new_n861), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT51), .B1(new_n873), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n843), .A2(new_n845), .B1(new_n575), .B2(new_n791), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(new_n870), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n867), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(KEYINPUT117), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n890), .B(new_n867), .C1(new_n883), .C2(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n817), .A2(new_n820), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT112), .B1(new_n253), .B2(new_n652), .ZN(new_n893));
  INV_X1    g707(.A(new_n740), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT112), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n713), .A2(new_n441), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n635), .A2(new_n897), .A3(new_n664), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n627), .B(new_n450), .C1(new_n573), .C2(new_n698), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n749), .A2(new_n774), .A3(new_n764), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n803), .A2(new_n574), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n712), .A2(new_n253), .ZN(new_n903));
  OAI22_X1  g717(.A1(new_n790), .A2(new_n902), .B1(new_n707), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n822), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n760), .A2(new_n900), .A3(new_n901), .A4(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n892), .A2(new_n906), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n715), .A2(new_n719), .B1(new_n737), .B2(new_n743), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n706), .A2(new_n575), .A3(new_n711), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n766), .A2(new_n909), .A3(new_n731), .A4(new_n803), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n794), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT52), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n794), .A2(new_n908), .A3(KEYINPUT52), .A4(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n907), .A2(new_n915), .A3(KEYINPUT53), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT114), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n907), .A2(new_n915), .A3(KEYINPUT114), .A4(KEYINPUT53), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT113), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n914), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n913), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n911), .A2(new_n921), .A3(new_n912), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT53), .B1(new_n925), .B2(new_n907), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT54), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(KEYINPUT53), .A3(new_n907), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT54), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n907), .A2(new_n915), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT53), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n889), .A2(new_n891), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(G952), .A2(G953), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n855), .B1(new_n935), .B2(new_n936), .ZN(G75));
  NOR2_X1   g751(.A1(new_n355), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n245), .B1(new_n928), .B2(new_n932), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT56), .B1(new_n940), .B2(G210), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n299), .B1(new_n330), .B2(new_n331), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n327), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n939), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n941), .A2(new_n944), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT118), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n941), .A2(KEYINPUT118), .A3(new_n944), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G51));
  NAND2_X1  g764(.A1(new_n928), .A2(new_n932), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT54), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n933), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n619), .B(KEYINPUT57), .Z(new_n955));
  OAI21_X1  g769(.A(new_n616), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n940), .A2(new_n832), .A3(new_n831), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n938), .B1(new_n956), .B2(new_n957), .ZN(G54));
  NAND3_X1  g772(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n959));
  INV_X1    g773(.A(new_n427), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n939), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT119), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n938), .B1(new_n959), .B2(new_n960), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT119), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n965), .B(new_n966), .C1(new_n960), .C2(new_n959), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(G60));
  XNOR2_X1  g782(.A(new_n640), .B(KEYINPUT120), .ZN(new_n969));
  NAND2_X1  g783(.A1(G478), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT59), .Z(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n934), .B2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n969), .A2(new_n972), .ZN(new_n974));
  INV_X1    g788(.A(new_n933), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n929), .B1(new_n928), .B2(new_n932), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n939), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT121), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n938), .B1(new_n953), .B2(new_n974), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT121), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n971), .B1(new_n927), .B2(new_n933), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n980), .B(new_n981), .C1(new_n982), .C2(new_n969), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n979), .A2(new_n983), .ZN(G63));
  INV_X1    g798(.A(new_n951), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n688), .A2(new_n690), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n451), .B(KEYINPUT122), .Z(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT60), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n693), .B1(new_n985), .B2(new_n988), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n989), .A2(new_n939), .A3(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n989), .A2(KEYINPUT61), .A3(new_n939), .A4(new_n990), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(G66));
  NAND3_X1  g809(.A1(new_n760), .A2(new_n900), .A3(new_n901), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT123), .Z(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n355), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n447), .B2(new_n325), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n942), .B1(G898), .B2(new_n355), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(G69));
  AOI21_X1  g816(.A(new_n355), .B1(G227), .B2(G900), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT125), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n562), .B(new_n405), .Z(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(G900), .B2(G953), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n848), .A2(new_n840), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n839), .A2(new_n723), .A3(new_n766), .A4(new_n857), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n794), .A2(new_n908), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1010), .B1(KEYINPUT126), .B2(new_n892), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1007), .B(new_n1011), .C1(KEYINPUT126), .C2(new_n892), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1006), .B1(new_n1012), .B2(G953), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT124), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1004), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1009), .A2(new_n735), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT62), .Z(new_n1017));
  INV_X1    g831(.A(new_n724), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1018), .A2(new_n897), .A3(new_n573), .A4(new_n822), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1007), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1005), .B1(new_n1021), .B2(G953), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n1013), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1015), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1022), .B(new_n1013), .C1(new_n1014), .C2(new_n1004), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n1024), .A2(new_n1025), .ZN(G72));
  XNOR2_X1  g840(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1027));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1029), .B1(new_n1012), .B2(new_n997), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1030), .A2(new_n546), .A3(new_n563), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1029), .B1(new_n1020), .B2(new_n997), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n938), .B1(new_n1032), .B2(new_n728), .ZN(new_n1033));
  INV_X1    g847(.A(new_n532), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n563), .A2(new_n531), .ZN(new_n1035));
  OAI221_X1 g849(.A(new_n1029), .B1(new_n1034), .B2(new_n1035), .C1(new_n920), .C2(new_n926), .ZN(new_n1036));
  AND3_X1   g850(.A1(new_n1031), .A2(new_n1033), .A3(new_n1036), .ZN(G57));
endmodule


