

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580;

  NOR2_X1 U320 ( .A1(n536), .A2(n399), .ZN(n400) );
  XOR2_X1 U321 ( .A(n460), .B(KEYINPUT68), .Z(n524) );
  XOR2_X1 U322 ( .A(G29GAT), .B(G36GAT), .Z(n288) );
  NOR2_X1 U323 ( .A1(n564), .A2(n554), .ZN(n395) );
  XNOR2_X1 U324 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U325 ( .A(n317), .B(n316), .ZN(n320) );
  XNOR2_X1 U326 ( .A(n409), .B(n327), .ZN(n328) );
  XNOR2_X1 U327 ( .A(n368), .B(n438), .ZN(n369) );
  XNOR2_X1 U328 ( .A(n329), .B(n328), .ZN(n447) );
  XNOR2_X1 U329 ( .A(n370), .B(n369), .ZN(n375) );
  XNOR2_X1 U330 ( .A(n377), .B(n376), .ZN(n378) );
  INV_X1 U331 ( .A(G183GAT), .ZN(n444) );
  XNOR2_X1 U332 ( .A(n379), .B(n378), .ZN(n525) );
  NOR2_X1 U333 ( .A1(n507), .A2(n496), .ZN(n504) );
  XOR2_X1 U334 ( .A(KEYINPUT38), .B(n467), .Z(n493) );
  XNOR2_X1 U335 ( .A(n444), .B(KEYINPUT124), .ZN(n445) );
  XNOR2_X1 U336 ( .A(n468), .B(G43GAT), .ZN(n469) );
  XNOR2_X1 U337 ( .A(n446), .B(n445), .ZN(G1350GAT) );
  XNOR2_X1 U338 ( .A(n470), .B(n469), .ZN(G1330GAT) );
  XOR2_X1 U339 ( .A(G211GAT), .B(G78GAT), .Z(n290) );
  XNOR2_X1 U340 ( .A(G22GAT), .B(G155GAT), .ZN(n289) );
  XNOR2_X1 U341 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U342 ( .A(G71GAT), .B(G127GAT), .Z(n292) );
  XNOR2_X1 U343 ( .A(G15GAT), .B(G183GAT), .ZN(n291) );
  XNOR2_X1 U344 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U345 ( .A(n294), .B(n293), .Z(n299) );
  XOR2_X1 U346 ( .A(G8GAT), .B(G1GAT), .Z(n377) );
  XOR2_X1 U347 ( .A(G57GAT), .B(KEYINPUT13), .Z(n392) );
  XOR2_X1 U348 ( .A(n392), .B(KEYINPUT78), .Z(n296) );
  NAND2_X1 U349 ( .A1(G231GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n377), .B(n297), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n307) );
  XOR2_X1 U353 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n301) );
  XNOR2_X1 U354 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U356 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n303) );
  XNOR2_X1 U357 ( .A(KEYINPUT77), .B(KEYINPUT12), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U359 ( .A(n305), .B(n304), .Z(n306) );
  XOR2_X1 U360 ( .A(n307), .B(n306), .Z(n548) );
  XOR2_X1 U361 ( .A(KEYINPUT3), .B(KEYINPUT89), .Z(n309) );
  XNOR2_X1 U362 ( .A(KEYINPUT88), .B(G155GAT), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U364 ( .A(KEYINPUT2), .B(n310), .Z(n347) );
  XOR2_X1 U365 ( .A(KEYINPUT85), .B(KEYINPUT24), .Z(n312) );
  XOR2_X1 U366 ( .A(G141GAT), .B(G22GAT), .Z(n364) );
  XOR2_X1 U367 ( .A(G50GAT), .B(G162GAT), .Z(n348) );
  XNOR2_X1 U368 ( .A(n364), .B(n348), .ZN(n311) );
  XOR2_X1 U369 ( .A(n312), .B(n311), .Z(n313) );
  XNOR2_X1 U370 ( .A(n347), .B(n313), .ZN(n317) );
  NAND2_X1 U371 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  INV_X1 U372 ( .A(KEYINPUT92), .ZN(n314) );
  XNOR2_X1 U373 ( .A(G106GAT), .B(G78GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n318), .B(G148GAT), .ZN(n385) );
  XNOR2_X1 U375 ( .A(n385), .B(KEYINPUT22), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n329) );
  XOR2_X1 U377 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n322) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(G211GAT), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U380 ( .A(G218GAT), .B(KEYINPUT21), .Z(n323) );
  XOR2_X1 U381 ( .A(n324), .B(n323), .Z(n409) );
  XOR2_X1 U382 ( .A(G204GAT), .B(KEYINPUT23), .Z(n326) );
  XNOR2_X1 U383 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U385 ( .A(G57GAT), .B(G120GAT), .Z(n331) );
  XNOR2_X1 U386 ( .A(G1GAT), .B(G113GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U388 ( .A(G85GAT), .B(G148GAT), .Z(n333) );
  XNOR2_X1 U389 ( .A(G141GAT), .B(G134GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n345) );
  XOR2_X1 U392 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n337) );
  XNOR2_X1 U393 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U395 ( .A(KEYINPUT4), .B(G162GAT), .Z(n339) );
  XOR2_X1 U396 ( .A(KEYINPUT0), .B(G127GAT), .Z(n433) );
  XNOR2_X1 U397 ( .A(G29GAT), .B(n433), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U399 ( .A(n341), .B(n340), .Z(n343) );
  NAND2_X1 U400 ( .A1(G225GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n509) );
  XOR2_X1 U404 ( .A(G85GAT), .B(G92GAT), .Z(n381) );
  XOR2_X1 U405 ( .A(n348), .B(n381), .Z(n350) );
  NAND2_X1 U406 ( .A1(G232GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U408 ( .A(KEYINPUT11), .B(G106GAT), .Z(n352) );
  XNOR2_X1 U409 ( .A(G190GAT), .B(G99GAT), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U411 ( .A(n354), .B(n353), .Z(n359) );
  XOR2_X1 U412 ( .A(G43GAT), .B(G134GAT), .Z(n437) );
  XOR2_X1 U413 ( .A(KEYINPUT64), .B(KEYINPUT67), .Z(n356) );
  XNOR2_X1 U414 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n437), .B(n357), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U418 ( .A(n360), .B(KEYINPUT9), .Z(n363) );
  XNOR2_X1 U419 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n288), .B(n361), .ZN(n365) );
  XNOR2_X1 U421 ( .A(n365), .B(KEYINPUT66), .ZN(n362) );
  XOR2_X1 U422 ( .A(n363), .B(n362), .Z(n558) );
  INV_X1 U423 ( .A(n558), .ZN(n536) );
  INV_X1 U424 ( .A(n548), .ZN(n573) );
  XNOR2_X1 U425 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n396) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n370) );
  XOR2_X1 U427 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n367) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n366) );
  XOR2_X1 U429 ( .A(n367), .B(n366), .Z(n368) );
  XOR2_X1 U430 ( .A(G113GAT), .B(G15GAT), .Z(n438) );
  XOR2_X1 U431 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n372) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(G197GAT), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n373), .B(KEYINPUT69), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n379) );
  XNOR2_X1 U436 ( .A(G50GAT), .B(G43GAT), .ZN(n376) );
  INV_X1 U437 ( .A(n525), .ZN(n564) );
  XNOR2_X1 U438 ( .A(G99GAT), .B(G71GAT), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n380), .B(G120GAT), .ZN(n430) );
  XNOR2_X1 U440 ( .A(n381), .B(n430), .ZN(n383) );
  AND2_X1 U441 ( .A1(G230GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n384), .B(KEYINPUT32), .ZN(n387) );
  XOR2_X1 U444 ( .A(n385), .B(KEYINPUT31), .Z(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U446 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n389) );
  XNOR2_X1 U447 ( .A(G176GAT), .B(KEYINPUT72), .ZN(n388) );
  XOR2_X1 U448 ( .A(n389), .B(n388), .Z(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n394) );
  XOR2_X1 U450 ( .A(G204GAT), .B(G64GAT), .Z(n413) );
  XNOR2_X1 U451 ( .A(n392), .B(n413), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n569) );
  XNOR2_X1 U453 ( .A(n569), .B(KEYINPUT41), .ZN(n554) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  NOR2_X1 U455 ( .A1(n573), .A2(n397), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n398), .B(KEYINPUT113), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(KEYINPUT47), .ZN(n406) );
  XOR2_X1 U458 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n402) );
  XOR2_X1 U459 ( .A(KEYINPUT36), .B(n558), .Z(n575) );
  NAND2_X1 U460 ( .A1(n573), .A2(n575), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n403) );
  NOR2_X1 U462 ( .A1(n403), .A2(n569), .ZN(n404) );
  NAND2_X1 U463 ( .A1(n404), .A2(n564), .ZN(n405) );
  NAND2_X1 U464 ( .A1(n406), .A2(n405), .ZN(n408) );
  XOR2_X1 U465 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n520) );
  INV_X1 U467 ( .A(n409), .ZN(n417) );
  XOR2_X1 U468 ( .A(KEYINPUT94), .B(G92GAT), .Z(n411) );
  XNOR2_X1 U469 ( .A(G8GAT), .B(G36GAT), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U471 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U474 ( .A(n417), .B(n416), .Z(n425) );
  XOR2_X1 U475 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n419) );
  XNOR2_X1 U476 ( .A(KEYINPUT82), .B(KEYINPUT17), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U478 ( .A(n420), .B(G176GAT), .Z(n422) );
  XNOR2_X1 U479 ( .A(G190GAT), .B(KEYINPUT81), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n424) );
  XOR2_X1 U481 ( .A(G169GAT), .B(G183GAT), .Z(n423) );
  XOR2_X1 U482 ( .A(n424), .B(n423), .Z(n442) );
  XOR2_X1 U483 ( .A(n425), .B(n442), .Z(n450) );
  NOR2_X1 U484 ( .A1(n520), .A2(n450), .ZN(n427) );
  INV_X1 U485 ( .A(KEYINPUT54), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  NOR2_X1 U487 ( .A1(n509), .A2(n428), .ZN(n563) );
  NAND2_X1 U488 ( .A1(n447), .A2(n563), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n429), .B(KEYINPUT55), .ZN(n443) );
  XOR2_X1 U490 ( .A(KEYINPUT80), .B(n430), .Z(n432) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n436) );
  XNOR2_X1 U493 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U495 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n521) );
  NAND2_X1 U499 ( .A1(n443), .A2(n521), .ZN(n559) );
  NOR2_X1 U500 ( .A1(n548), .A2(n559), .ZN(n446) );
  XOR2_X1 U501 ( .A(KEYINPUT27), .B(n450), .Z(n458) );
  NOR2_X1 U502 ( .A1(n447), .A2(n521), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n448), .B(KEYINPUT26), .ZN(n562) );
  AND2_X1 U504 ( .A1(n458), .A2(n562), .ZN(n449) );
  XOR2_X1 U505 ( .A(KEYINPUT95), .B(n449), .Z(n454) );
  INV_X1 U506 ( .A(n450), .ZN(n512) );
  NAND2_X1 U507 ( .A1(n512), .A2(n521), .ZN(n451) );
  NAND2_X1 U508 ( .A1(n447), .A2(n451), .ZN(n452) );
  XNOR2_X1 U509 ( .A(KEYINPUT25), .B(n452), .ZN(n453) );
  NOR2_X1 U510 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n455), .B(KEYINPUT96), .ZN(n456) );
  NOR2_X1 U512 ( .A1(n456), .A2(n509), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n457), .B(KEYINPUT97), .ZN(n464) );
  NAND2_X1 U514 ( .A1(n509), .A2(n458), .ZN(n519) );
  XNOR2_X1 U515 ( .A(KEYINPUT84), .B(n521), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n519), .A2(n459), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n447), .B(KEYINPUT28), .ZN(n460) );
  INV_X1 U518 ( .A(n524), .ZN(n461) );
  NAND2_X1 U519 ( .A1(n462), .A2(n461), .ZN(n463) );
  NAND2_X1 U520 ( .A1(n464), .A2(n463), .ZN(n473) );
  AND2_X1 U521 ( .A1(n548), .A2(n575), .ZN(n465) );
  AND2_X1 U522 ( .A1(n473), .A2(n465), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n466), .B(KEYINPUT37), .ZN(n508) );
  OR2_X1 U524 ( .A1(n564), .A2(n569), .ZN(n475) );
  OR2_X1 U525 ( .A1(n508), .A2(n475), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n493), .A2(n521), .ZN(n470) );
  XOR2_X1 U527 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n468) );
  NAND2_X1 U528 ( .A1(n573), .A2(n558), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT16), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(KEYINPUT79), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n496) );
  NOR2_X1 U532 ( .A1(n475), .A2(n496), .ZN(n486) );
  NAND2_X1 U533 ( .A1(n509), .A2(n486), .ZN(n479) );
  XOR2_X1 U534 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n477) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U538 ( .A(KEYINPUT98), .B(n480), .ZN(G1324GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n482) );
  NAND2_X1 U540 ( .A1(n486), .A2(n512), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U544 ( .A1(n486), .A2(n521), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U546 ( .A1(n524), .A2(n486), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n487), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U548 ( .A1(n493), .A2(n509), .ZN(n490) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n493), .A2(n512), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  XNOR2_X1 U555 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n495) );
  NAND2_X1 U556 ( .A1(n524), .A2(n493), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1331GAT) );
  INV_X1 U558 ( .A(n554), .ZN(n528) );
  NAND2_X1 U559 ( .A1(n564), .A2(n528), .ZN(n507) );
  NAND2_X1 U560 ( .A1(n509), .A2(n504), .ZN(n500) );
  XOR2_X1 U561 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n498) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(G1332GAT) );
  NAND2_X1 U565 ( .A1(n504), .A2(n512), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U567 ( .A(G71GAT), .B(KEYINPUT109), .Z(n503) );
  NAND2_X1 U568 ( .A1(n504), .A2(n521), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n503), .B(n502), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(G78GAT), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U571 ( .A1(n504), .A2(n524), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(G1335GAT) );
  NOR2_X1 U573 ( .A1(n508), .A2(n507), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n509), .A2(n516), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(KEYINPUT110), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U577 ( .A1(n516), .A2(n512), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U579 ( .A(G99GAT), .B(KEYINPUT111), .Z(n515) );
  NAND2_X1 U580 ( .A1(n516), .A2(n521), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(G1338GAT) );
  NAND2_X1 U582 ( .A1(n524), .A2(n516), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(KEYINPUT44), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n518), .ZN(G1339GAT) );
  XNOR2_X1 U585 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n527) );
  NOR2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n542) );
  NAND2_X1 U587 ( .A1(n542), .A2(n521), .ZN(n522) );
  XOR2_X1 U588 ( .A(KEYINPUT115), .B(n522), .Z(n523) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n537), .A2(n525), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT117), .Z(n530) );
  NAND2_X1 U593 ( .A1(n537), .A2(n528), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n534) );
  NAND2_X1 U598 ( .A1(n537), .A2(n573), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT121), .Z(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n542), .A2(n562), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n564), .A2(n550), .ZN(n543) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n547) );
  NOR2_X1 U612 ( .A1(n554), .A2(n550), .ZN(n546) );
  XOR2_X1 U613 ( .A(n547), .B(n546), .Z(G1345GAT) );
  NOR2_X1 U614 ( .A1(n548), .A2(n550), .ZN(n549) );
  XOR2_X1 U615 ( .A(G155GAT), .B(n549), .Z(G1346GAT) );
  NOR2_X1 U616 ( .A1(n558), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G162GAT), .B(KEYINPUT123), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1347GAT) );
  NOR2_X1 U619 ( .A1(n564), .A2(n559), .ZN(n553) );
  XOR2_X1 U620 ( .A(G169GAT), .B(n553), .Z(G1348GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n559), .ZN(n556) );
  XNOR2_X1 U622 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(n557), .ZN(G1349GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(G190GAT), .B(n560), .Z(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT58), .B(n561), .ZN(G1351GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n568) );
  NOR2_X1 U629 ( .A1(n564), .A2(n568), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n571) );
  INV_X1 U634 ( .A(n568), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n576), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n576), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT127), .B(KEYINPUT126), .Z(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1355GAT) );
endmodule

