//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  OAI221_X1 g0009(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n202), .C2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT66), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n210), .A2(new_n211), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n205), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  AND3_X1   g0018(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n219));
  AOI21_X1  g0019(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OR3_X1    g0026(.A1(new_n205), .A2(KEYINPUT64), .A3(G13), .ZN(new_n227));
  OAI21_X1  g0027(.A(KEYINPUT64), .B1(new_n205), .B2(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n218), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n217), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  INV_X1    g0043(.A(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT68), .B(G50), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NOR2_X1   g0051(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n252));
  INV_X1    g0052(.A(G97), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT81), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT81), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G97), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(G20), .B1(G33), .B2(G283), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n252), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT65), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G116), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G20), .ZN(new_n269));
  AND3_X1   g0069(.A1(new_n267), .A2(KEYINPUT85), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT85), .B1(new_n267), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n261), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT86), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT20), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n261), .B1(new_n273), .B2(new_n274), .C1(new_n270), .C2(new_n271), .ZN(new_n277));
  INV_X1    g0077(.A(new_n267), .ZN(new_n278));
  INV_X1    g0078(.A(G1), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G13), .A3(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G116), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n268), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n276), .A2(new_n277), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  OAI211_X1 g0088(.A(G264), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  OAI211_X1 g0090(.A(G257), .B(new_n290), .C1(new_n287), .C2(new_n288), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT3), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n258), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G303), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n289), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(new_n219), .B2(new_n220), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT5), .B(G41), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n297), .A2(G1), .A3(G13), .ZN(new_n302));
  INV_X1    g0102(.A(G45), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G1), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n301), .A2(G274), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n262), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n301), .A2(new_n304), .B1(new_n306), .B2(new_n297), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT84), .B1(new_n307), .B2(G270), .ZN(new_n308));
  AND2_X1   g0108(.A1(KEYINPUT5), .A2(G41), .ZN(new_n309));
  NOR2_X1   g0109(.A1(KEYINPUT5), .A2(G41), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n304), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AND4_X1   g0111(.A1(KEYINPUT84), .A2(new_n311), .A3(G270), .A4(new_n302), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n300), .B(new_n305), .C1(new_n308), .C2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  INV_X1    g0116(.A(new_n305), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT84), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n311), .A2(new_n302), .ZN(new_n319));
  INV_X1    g0119(.A(G270), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n307), .A2(KEYINPUT84), .A3(G270), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n317), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n316), .B1(new_n323), .B2(new_n300), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n286), .A2(new_n315), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n313), .A2(KEYINPUT21), .A3(G169), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(G179), .A3(new_n300), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n272), .A2(new_n275), .B1(new_n283), .B2(new_n284), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n326), .A2(new_n327), .B1(new_n328), .B2(new_n277), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n323), .B2(new_n300), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT21), .B1(new_n286), .B2(new_n331), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n325), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n287), .A2(new_n288), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G77), .ZN(new_n335));
  OAI211_X1 g0135(.A(G222), .B(new_n290), .C1(new_n287), .C2(new_n288), .ZN(new_n336));
  OAI211_X1 g0136(.A(G223), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT70), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n335), .A2(KEYINPUT70), .A3(new_n336), .A4(new_n337), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n299), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(G33), .A2(G41), .ZN(new_n343));
  OAI21_X1  g0143(.A(G274), .B1(new_n343), .B2(new_n262), .ZN(new_n344));
  INV_X1    g0144(.A(G41), .ZN(new_n345));
  AOI21_X1  g0145(.A(G1), .B1(new_n345), .B2(new_n303), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT69), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n279), .B1(G41), .B2(G45), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT69), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n344), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n302), .A2(new_n349), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(G226), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n342), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(G20), .A2(G33), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G150), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT8), .B(G58), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n222), .A2(G33), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n201), .A2(new_n222), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n267), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n264), .A2(new_n280), .A3(new_n265), .A4(new_n266), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n279), .A2(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(G50), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n280), .ZN(new_n370));
  INV_X1    g0170(.A(G50), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n365), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n358), .B(new_n373), .C1(G169), .C2(new_n356), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n355), .A2(G200), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n342), .A2(G190), .A3(new_n354), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT9), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n365), .A2(new_n369), .A3(KEYINPUT9), .A4(new_n372), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n376), .A2(new_n377), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT10), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n316), .B1(new_n342), .B2(new_n354), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT10), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(new_n377), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n375), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n359), .A2(G50), .B1(G20), .B2(new_n207), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n202), .B2(new_n362), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n267), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT11), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n367), .A2(G68), .A3(new_n368), .ZN(new_n394));
  OR2_X1    g0194(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n395));
  NAND2_X1  g0195(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n395), .B(new_n396), .C1(new_n280), .C2(G68), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n370), .A2(new_n207), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT79), .B(new_n397), .C1(new_n398), .C2(KEYINPUT12), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n394), .B(new_n399), .C1(KEYINPUT79), .C2(new_n397), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G274), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n306), .B2(new_n297), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n346), .A2(new_n347), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n349), .A2(KEYINPUT69), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n353), .A2(G238), .ZN(new_n407));
  NOR2_X1   g0207(.A1(G226), .A2(G1698), .ZN(new_n408));
  INV_X1    g0208(.A(G232), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n293), .A2(new_n294), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n410), .A2(new_n411), .B1(G33), .B2(G97), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n406), .B(new_n407), .C1(new_n412), .C2(new_n298), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(KEYINPUT13), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n352), .A2(new_n208), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n351), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n409), .A2(G1698), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n418), .B1(G226), .B2(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G97), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n299), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n415), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n401), .B1(new_n424), .B2(new_n316), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT77), .ZN(new_n427));
  AOI211_X1 g0227(.A(KEYINPUT76), .B(new_n415), .C1(new_n417), .C2(new_n422), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT76), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n413), .B2(KEYINPUT13), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n406), .A2(new_n407), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n412), .A2(new_n298), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n314), .B1(new_n434), .B2(new_n415), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n427), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n413), .A2(KEYINPUT13), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT76), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n423), .A2(new_n429), .ZN(new_n439));
  AND4_X1   g0239(.A1(new_n427), .A2(new_n435), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n426), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(G169), .B1(new_n414), .B2(new_n423), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT14), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n414), .A2(new_n357), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(new_n439), .A3(new_n438), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(G169), .C1(new_n414), .C2(new_n423), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n401), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n388), .A2(new_n441), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G87), .ZN(new_n452));
  INV_X1    g0252(.A(G223), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n290), .ZN(new_n454));
  INV_X1    g0254(.A(G226), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G1698), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n454), .B(new_n456), .C1(new_n287), .C2(new_n288), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n298), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n302), .A2(G232), .A3(new_n349), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n458), .A2(new_n351), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n357), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(G169), .B2(new_n460), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n293), .A2(new_n222), .A3(new_n294), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT7), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n293), .A2(KEYINPUT7), .A3(new_n222), .A4(new_n294), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n207), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n244), .A2(new_n207), .ZN(new_n468));
  NOR2_X1   g0268(.A1(G58), .A2(G68), .ZN(new_n469));
  OAI21_X1  g0269(.A(G20), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n359), .A2(G159), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT80), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT16), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT16), .ZN(new_n475));
  OAI211_X1 g0275(.A(KEYINPUT80), .B(new_n475), .C1(new_n467), .C2(new_n472), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n267), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n361), .B1(new_n279), .B2(G20), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(new_n367), .B1(new_n370), .B2(new_n361), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n462), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT18), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n479), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n278), .B1(new_n473), .B2(KEYINPUT16), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n476), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT18), .B1(new_n485), .B2(new_n462), .ZN(new_n486));
  NOR4_X1   g0286(.A1(new_n458), .A2(new_n351), .A3(new_n314), .A4(new_n459), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n457), .A2(new_n452), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n459), .B1(new_n488), .B2(new_n299), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n316), .B1(new_n489), .B2(new_n406), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT80), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT7), .B1(new_n334), .B2(new_n222), .ZN(new_n493));
  INV_X1    g0293(.A(new_n466), .ZN(new_n494));
  OAI21_X1  g0294(.A(G68), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n472), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n267), .B1(new_n497), .B2(new_n475), .ZN(new_n498));
  INV_X1    g0298(.A(new_n476), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n491), .B(new_n479), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT17), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n485), .A2(KEYINPUT17), .A3(new_n491), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n482), .A2(new_n486), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  XOR2_X1   g0305(.A(KEYINPUT8), .B(G58), .Z(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(new_n359), .B1(G20), .B2(G77), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT15), .B(G87), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n362), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n267), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n370), .A2(new_n202), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n511), .B(KEYINPUT72), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n368), .A2(G77), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n366), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n514), .A2(KEYINPUT73), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(KEYINPUT73), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n510), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n406), .B1(new_n209), .B2(new_n352), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n411), .A2(G232), .A3(new_n290), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n411), .A2(G238), .A3(G1698), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n334), .A2(G107), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT71), .A4(new_n521), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n522), .A2(new_n299), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT71), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n518), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n517), .B1(new_n527), .B2(G169), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT74), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n299), .A3(new_n522), .ZN(new_n530));
  INV_X1    g0330(.A(new_n518), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n529), .B1(new_n532), .B2(G179), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n527), .A2(KEYINPUT74), .A3(new_n357), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n528), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT75), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n517), .B1(G190), .B2(new_n527), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n532), .A2(G200), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n540), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT75), .B1(new_n542), .B2(new_n535), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n505), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n451), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n311), .A2(G257), .A3(new_n302), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n305), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT82), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G250), .A2(G1698), .ZN(new_n549));
  NAND2_X1  g0349(.A1(KEYINPUT4), .A2(G244), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(G1698), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n411), .A2(new_n551), .B1(G33), .B2(G283), .ZN(new_n552));
  OAI211_X1 g0352(.A(G244), .B(new_n290), .C1(new_n287), .C2(new_n288), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT4), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n299), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT82), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n546), .A2(new_n558), .A3(new_n305), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n548), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n330), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n546), .A2(new_n558), .A3(new_n305), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n558), .B1(new_n546), .B2(new_n305), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(G179), .B1(new_n556), .B2(new_n299), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G107), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n465), .B2(new_n466), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n253), .B2(KEYINPUT6), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT6), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(G97), .A3(G107), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT6), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n573), .A3(G20), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n359), .A2(G77), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n267), .B1(new_n568), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n280), .A2(G97), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n366), .B1(new_n279), .B2(G33), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n561), .A2(new_n566), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n548), .A2(new_n557), .A3(G190), .A4(new_n559), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(new_n577), .A3(new_n580), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n316), .B1(new_n564), .B2(new_n557), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT83), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n581), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n560), .A2(G200), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT83), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n583), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n582), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G257), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n592));
  OAI211_X1 g0392(.A(G250), .B(new_n290), .C1(new_n287), .C2(new_n288), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G33), .A2(G294), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(new_n299), .B1(new_n307), .B2(G264), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(new_n314), .A3(new_n305), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n305), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n599), .B2(G200), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT22), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n222), .B(G87), .C1(new_n287), .C2(new_n288), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT88), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(G20), .B1(new_n293), .B2(new_n294), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n601), .A2(KEYINPUT87), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n605), .A2(KEYINPUT88), .A3(G87), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(KEYINPUT87), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT23), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n222), .B2(G107), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n567), .A2(KEYINPUT23), .A3(G20), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n258), .A2(new_n268), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n610), .A2(new_n611), .B1(new_n612), .B2(new_n222), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n604), .A2(new_n607), .A3(new_n608), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT24), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n608), .A2(new_n613), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT24), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n604), .A4(new_n607), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n267), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT25), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n280), .B2(G107), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n370), .A2(KEYINPUT25), .A3(new_n567), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n579), .A2(G107), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n600), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n599), .A2(new_n357), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n598), .A2(new_n330), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n278), .B1(new_n615), .B2(new_n618), .ZN(new_n628));
  INV_X1    g0428(.A(new_n624), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT19), .ZN(new_n631));
  XNOR2_X1  g0431(.A(KEYINPUT81), .B(G97), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n362), .ZN(new_n633));
  NOR2_X1   g0433(.A1(G87), .A2(G107), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n254), .A2(new_n256), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n222), .B1(new_n420), .B2(new_n631), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n411), .A2(new_n222), .A3(G68), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n633), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n267), .B1(new_n370), .B2(new_n508), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n579), .A2(G87), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n612), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n208), .A2(new_n290), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n209), .A2(G1698), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n645), .B(new_n646), .C1(new_n287), .C2(new_n288), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n298), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G250), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n279), .B2(G45), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n302), .ZN(new_n651));
  INV_X1    g0451(.A(new_n304), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n344), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(G200), .B1(new_n648), .B2(new_n653), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n403), .A2(new_n304), .B1(new_n302), .B2(new_n650), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n645), .A2(new_n646), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n612), .B1(new_n656), .B2(new_n411), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n655), .B(G190), .C1(new_n657), .C2(new_n298), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n330), .B1(new_n648), .B2(new_n653), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n655), .B(new_n357), .C1(new_n657), .C2(new_n298), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n639), .A2(new_n267), .ZN(new_n663));
  INV_X1    g0463(.A(new_n508), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n579), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n508), .A2(new_n370), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n643), .A2(new_n659), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n625), .A2(new_n630), .A3(new_n668), .ZN(new_n669));
  AND4_X1   g0469(.A1(new_n333), .A2(new_n545), .A3(new_n591), .A4(new_n669), .ZN(G372));
  NAND2_X1  g0470(.A1(new_n286), .A2(new_n331), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT21), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n326), .A2(new_n327), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n286), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n673), .A2(new_n675), .A3(new_n630), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n667), .A2(new_n661), .A3(new_n660), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT89), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n654), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g0479(.A(KEYINPUT89), .B(G200), .C1(new_n648), .C2(new_n653), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n658), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n677), .B1(new_n681), .B2(new_n642), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n628), .A2(new_n629), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(new_n600), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n591), .A2(new_n676), .A3(new_n684), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n564), .A2(new_n565), .B1(new_n577), .B2(new_n580), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n640), .A2(new_n658), .A3(new_n641), .A4(new_n654), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n686), .A2(new_n677), .A3(new_n561), .A4(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT90), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n582), .A2(new_n668), .A3(new_n691), .A4(KEYINPUT26), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n686), .A2(new_n561), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n689), .B1(new_n682), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n685), .A2(new_n695), .A3(new_n677), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n545), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n482), .A2(new_n486), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n441), .A2(new_n535), .B1(new_n449), .B2(new_n448), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n502), .A2(new_n503), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT91), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n381), .A2(KEYINPUT10), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n386), .B1(new_n385), .B2(new_n377), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n382), .A2(new_n387), .A3(KEYINPUT91), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n375), .B1(new_n701), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n697), .A2(new_n708), .ZN(G369));
  NAND2_X1  g0509(.A1(new_n673), .A2(new_n675), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n279), .A2(new_n222), .A3(G13), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G213), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G343), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n286), .A2(new_n716), .ZN(new_n717));
  MUX2_X1   g0517(.A(new_n710), .B(new_n333), .S(new_n717), .Z(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT92), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  INV_X1    g0520(.A(new_n716), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n625), .B(new_n630), .C1(new_n683), .C2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n630), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n716), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT93), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(new_n724), .A3(KEYINPUT93), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n720), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n710), .A2(new_n721), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n728), .A2(new_n733), .B1(new_n723), .B2(new_n721), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(G399));
  INV_X1    g0535(.A(new_n229), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G41), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n635), .A2(G116), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n737), .A2(new_n279), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n225), .B2(new_n737), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT28), .Z(new_n742));
  INV_X1    g0542(.A(KEYINPUT29), .ZN(new_n743));
  INV_X1    g0543(.A(new_n682), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(KEYINPUT26), .A3(new_n582), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n688), .A2(KEYINPUT94), .A3(new_n689), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT94), .B1(new_n688), .B2(new_n689), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n685), .B(new_n677), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n743), .B1(new_n749), .B2(new_n721), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n696), .A2(new_n743), .A3(new_n721), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n669), .A2(new_n333), .A3(new_n591), .A4(new_n721), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n648), .A2(new_n653), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n564), .A2(new_n557), .A3(new_n755), .A4(new_n596), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n754), .B1(new_n756), .B2(new_n327), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n755), .A2(new_n596), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n560), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n313), .A2(new_n357), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n759), .A2(KEYINPUT30), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n755), .A2(G179), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n560), .A2(new_n762), .A3(new_n313), .A4(new_n598), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n757), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT31), .B1(new_n764), .B2(new_n716), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n764), .A2(KEYINPUT31), .A3(new_n716), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n753), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G330), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n752), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n742), .B1(new_n771), .B2(G1), .ZN(G364));
  NOR2_X1   g0572(.A1(new_n222), .A2(G179), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(new_n314), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT97), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G283), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n222), .A2(new_n357), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(G190), .A3(new_n316), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n334), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n773), .A2(new_n785), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n784), .B(new_n788), .C1(G329), .C2(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n314), .A2(G179), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n222), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n781), .A2(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n314), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT99), .B(G326), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G294), .A2(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n795), .A2(G190), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT33), .B(G317), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n799), .A2(new_n800), .B1(new_n802), .B2(G303), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n780), .A2(new_n791), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n411), .B1(new_n786), .B2(new_n202), .C1(new_n244), .C2(new_n782), .ZN(new_n805));
  INV_X1    g0605(.A(G159), .ZN(new_n806));
  OAI21_X1  g0606(.A(KEYINPUT32), .B1(new_n789), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n796), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n371), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n802), .A2(G87), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n789), .A2(KEYINPUT32), .A3(new_n806), .ZN(new_n812));
  OR4_X1    g0612(.A1(new_n805), .A2(new_n809), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n799), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n814), .A2(new_n207), .B1(new_n253), .B2(new_n793), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT98), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n779), .A2(G107), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(KEYINPUT98), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n804), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n221), .B1(G20), .B2(new_n330), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G13), .A2(G33), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n229), .A2(new_n411), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT96), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G355), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(G116), .B2(new_n229), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n736), .A2(new_n411), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(G45), .B2(new_n224), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n247), .B2(G45), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n826), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G13), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n835), .A2(new_n303), .A3(G20), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT95), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(KEYINPUT95), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n837), .A2(G1), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n737), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n822), .A2(new_n834), .A3(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT100), .Z(new_n843));
  INV_X1    g0643(.A(new_n825), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n718), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n841), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n720), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n719), .A2(G330), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT101), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G396));
  NAND2_X1  g0651(.A1(new_n535), .A2(new_n721), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n538), .A2(new_n539), .B1(new_n517), .B2(new_n716), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n535), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n696), .B2(new_n721), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n542), .A2(new_n535), .A3(new_n716), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n696), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n770), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT103), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n858), .A2(new_n770), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n841), .B1(new_n861), .B2(KEYINPUT104), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n860), .B(new_n862), .C1(KEYINPUT104), .C2(new_n861), .ZN(new_n863));
  INV_X1    g0663(.A(new_n782), .ZN(new_n864));
  INV_X1    g0664(.A(new_n786), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n864), .A2(G143), .B1(new_n865), .B2(G159), .ZN(new_n866));
  INV_X1    g0666(.A(G137), .ZN(new_n867));
  INV_X1    g0667(.A(G150), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n866), .B1(new_n808), .B2(new_n867), .C1(new_n868), .C2(new_n814), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT34), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n779), .A2(G68), .ZN(new_n873));
  INV_X1    g0673(.A(G132), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n411), .B1(new_n789), .B2(new_n874), .C1(new_n793), .C2(new_n244), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(G50), .B2(new_n802), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n779), .A2(G87), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n787), .B2(new_n789), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT102), .Z(new_n880));
  INV_X1    g0680(.A(G283), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n814), .A2(new_n881), .B1(new_n253), .B2(new_n793), .ZN(new_n882));
  INV_X1    g0682(.A(G303), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n808), .A2(new_n883), .B1(new_n801), .B2(new_n567), .ZN(new_n884));
  INV_X1    g0684(.A(G294), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n334), .B1(new_n786), .B2(new_n268), .C1(new_n885), .C2(new_n782), .ZN(new_n886));
  OR3_X1    g0686(.A1(new_n882), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n877), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n821), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n821), .A2(new_n823), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n846), .B1(new_n890), .B2(new_n202), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n889), .B(new_n891), .C1(new_n855), .C2(new_n824), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n863), .A2(new_n892), .ZN(G384));
  NAND2_X1  g0693(.A1(new_n572), .A2(new_n573), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT35), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n223), .B(G116), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT36), .Z(new_n898));
  OAI21_X1  g0698(.A(G77), .B1(new_n244), .B2(new_n207), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n899), .A2(new_n224), .B1(G50), .B2(new_n207), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(G1), .A3(new_n835), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT105), .Z(new_n903));
  XNOR2_X1  g0703(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT108), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n768), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n764), .A2(KEYINPUT31), .A3(new_n716), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n765), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT108), .A3(new_n753), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n449), .A2(new_n716), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n450), .A2(new_n441), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT77), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n431), .A2(new_n427), .A3(new_n435), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n425), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n449), .B(new_n716), .C1(new_n916), .C2(new_n448), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n854), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n907), .A2(new_n910), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n500), .B1(new_n485), .B2(new_n462), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n485), .A2(new_n714), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n477), .A2(new_n479), .ZN(new_n923));
  INV_X1    g0723(.A(new_n714), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(KEYINPUT106), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT106), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n485), .B2(new_n714), .ZN(new_n927));
  INV_X1    g0727(.A(new_n462), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n925), .A2(new_n927), .A3(new_n929), .A4(new_n500), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n922), .B1(new_n930), .B2(KEYINPUT37), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n504), .A2(new_n921), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n931), .A2(KEYINPUT38), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT38), .B1(new_n931), .B2(new_n932), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n905), .B1(new_n919), .B2(new_n935), .ZN(new_n936));
  AND4_X1   g0736(.A1(KEYINPUT108), .A2(new_n753), .A3(new_n766), .A4(new_n767), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT108), .B1(new_n909), .B2(new_n753), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT38), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n930), .A2(KEYINPUT37), .ZN(new_n941));
  INV_X1    g0741(.A(new_n920), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT37), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n942), .A2(new_n943), .A3(new_n927), .A4(new_n925), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n925), .A2(new_n927), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n941), .A2(new_n944), .B1(new_n504), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n940), .B1(new_n946), .B2(KEYINPUT38), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n939), .A2(KEYINPUT40), .A3(new_n947), .A4(new_n918), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n936), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n939), .A2(new_n545), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(G330), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n698), .A2(new_n924), .ZN(new_n954));
  INV_X1    g0754(.A(new_n935), .ZN(new_n955));
  INV_X1    g0755(.A(new_n852), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n696), .B2(new_n857), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n917), .A2(new_n912), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n954), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT39), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n941), .A2(new_n944), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n504), .A2(new_n945), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT38), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n962), .B1(new_n965), .B2(new_n933), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n448), .A2(new_n449), .A3(new_n721), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n931), .A2(new_n932), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT38), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(KEYINPUT39), .A3(new_n940), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n966), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n961), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n545), .B1(new_n750), .B2(new_n751), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n708), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n974), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n953), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(G1), .B1(new_n835), .B2(G20), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n953), .A2(new_n977), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n903), .B1(new_n980), .B2(new_n981), .ZN(G367));
  AND2_X1   g0782(.A1(new_n831), .A2(new_n236), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n826), .B1(new_n229), .B2(new_n508), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n841), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n411), .B1(new_n789), .B2(new_n867), .C1(new_n782), .C2(new_n868), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n794), .A2(G68), .ZN(new_n987));
  INV_X1    g0787(.A(G143), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n808), .B2(new_n988), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n986), .B(new_n989), .C1(G58), .C2(new_n802), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n814), .A2(new_n806), .B1(new_n786), .B2(new_n371), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT113), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n779), .A2(G77), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n992), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n990), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n864), .A2(G303), .B1(new_n865), .B2(G283), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n802), .A2(KEYINPUT46), .A3(G116), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n801), .B2(new_n268), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n411), .B1(new_n790), .B2(G317), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G294), .A2(new_n799), .B1(new_n796), .B2(G311), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n567), .B2(new_n793), .C1(new_n632), .C2(new_n778), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n996), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT115), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1005), .B(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n985), .B1(new_n1008), .B2(new_n821), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n642), .A2(new_n716), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n744), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n677), .B2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1009), .B1(new_n844), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n728), .B(new_n733), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT111), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n719), .A2(new_n1015), .A3(G330), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1015), .B1(new_n719), .B2(G330), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1014), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT112), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(new_n1022), .A3(new_n771), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n591), .B1(new_n587), .B2(new_n721), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n582), .A2(new_n716), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n734), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT45), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT45), .B1(new_n734), .B2(new_n1026), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n734), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1026), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT44), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT44), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n734), .A2(new_n1034), .A3(new_n1026), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n1029), .A2(new_n1030), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT110), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n731), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1019), .A2(new_n1020), .A3(new_n771), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(KEYINPUT112), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1036), .A2(new_n1037), .A3(new_n730), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1023), .A2(new_n1039), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n771), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n737), .B(KEYINPUT41), .Z(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n840), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1026), .B(KEYINPUT109), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n723), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n716), .B1(new_n1050), .B2(new_n693), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n728), .A2(new_n733), .A3(new_n1026), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT42), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1048), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n730), .A2(new_n1049), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1013), .B1(new_n1047), .B2(new_n1058), .ZN(G387));
  NAND2_X1  g0859(.A1(new_n1023), .A2(new_n1041), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n737), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1021), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n771), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n729), .A2(new_n825), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n821), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n864), .A2(G317), .B1(new_n865), .B2(G303), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n808), .B2(new_n783), .C1(new_n787), .C2(new_n814), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n794), .A2(G283), .B1(new_n802), .B2(G294), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1075), .A2(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(KEYINPUT49), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n778), .A2(new_n268), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n411), .B(new_n1078), .C1(new_n790), .C2(new_n797), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n814), .A2(new_n361), .B1(new_n801), .B2(new_n202), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n664), .B2(new_n794), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n796), .A2(G159), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT116), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n411), .B1(new_n786), .B2(new_n207), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n782), .A2(new_n371), .B1(new_n789), .B2(new_n868), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(KEYINPUT116), .C2(new_n1083), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n779), .A2(G97), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1082), .A2(new_n1084), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1067), .B1(new_n1080), .B2(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n828), .A2(new_n739), .B1(new_n567), .B2(new_n736), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n241), .A2(new_n303), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n506), .A2(new_n371), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT50), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n738), .B(new_n303), .C1(new_n207), .C2(new_n202), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n831), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1091), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n846), .B(new_n1090), .C1(new_n826), .C2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1021), .A2(new_n840), .B1(new_n1066), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1065), .A2(new_n1099), .ZN(G393));
  AND2_X1   g0900(.A1(new_n1023), .A2(new_n1041), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1036), .B(new_n731), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1043), .B(new_n737), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1049), .A2(new_n844), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n411), .B1(new_n789), .B2(new_n988), .C1(new_n361), .C2(new_n786), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n814), .A2(new_n371), .B1(new_n202), .B2(new_n793), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G68), .C2(new_n802), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n808), .A2(new_n868), .B1(new_n806), .B2(new_n782), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT51), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n878), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G317), .A2(new_n796), .B1(new_n864), .B2(G311), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT52), .Z(new_n1114));
  OAI21_X1  g0914(.A(new_n334), .B1(new_n786), .B2(new_n885), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G322), .B2(new_n790), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n814), .A2(new_n883), .B1(new_n801), .B2(new_n881), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G116), .B2(new_n794), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1114), .A2(new_n817), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1067), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n831), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n826), .B1(new_n229), .B2(new_n632), .C1(new_n1121), .C2(new_n250), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT117), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n846), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1123), .B2(new_n1122), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1104), .A2(new_n1120), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1102), .B2(new_n840), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1103), .A2(new_n1127), .ZN(G390));
  NAND2_X1  g0928(.A1(new_n966), .A2(new_n972), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT118), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1130), .B(new_n967), .C1(new_n957), .C2(new_n959), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n967), .B1(new_n957), .B2(new_n959), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT118), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1129), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n947), .A2(new_n967), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n853), .A2(new_n535), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n749), .A2(new_n721), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n959), .B1(new_n1138), .B2(new_n852), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n768), .A2(new_n958), .A3(G330), .A4(new_n855), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1134), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n966), .A2(new_n972), .B1(new_n1132), .B2(KEYINPUT118), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n1131), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n907), .A2(G330), .A3(new_n910), .A4(new_n918), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n545), .A2(new_n907), .A3(G330), .A4(new_n910), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n975), .A2(new_n1148), .A3(new_n708), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n959), .B1(new_n769), .B2(new_n854), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1146), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n957), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n907), .A2(G330), .A3(new_n855), .A4(new_n910), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n959), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1141), .A2(new_n852), .A3(new_n1138), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1149), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1147), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1142), .B(new_n1158), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n737), .A3(new_n1161), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1147), .A2(new_n839), .ZN(new_n1163));
  INV_X1    g0963(.A(G128), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n1164), .A2(new_n808), .B1(new_n814), .B2(new_n867), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G159), .B2(new_n794), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT54), .B(G143), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n782), .A2(new_n874), .B1(new_n786), .B2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n334), .B(new_n1168), .C1(G125), .C2(new_n790), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n801), .A2(new_n868), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT53), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n779), .A2(G50), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1166), .A2(new_n1169), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n782), .A2(new_n268), .B1(new_n786), .B2(new_n632), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n411), .B(new_n1174), .C1(G294), .C2(new_n790), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n811), .B1(G77), .B2(new_n794), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G107), .A2(new_n799), .B1(new_n796), .B2(G283), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1175), .A2(new_n873), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1067), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n846), .B(new_n1179), .C1(new_n361), .C2(new_n890), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1129), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n824), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1162), .A2(new_n1163), .A3(new_n1182), .ZN(G378));
  INV_X1    g0983(.A(KEYINPUT120), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n705), .A2(new_n374), .A3(new_n706), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n373), .A2(new_n924), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n705), .A2(new_n374), .A3(new_n706), .A4(new_n1186), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1184), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1190), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(KEYINPUT120), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1193), .A2(new_n1198), .A3(new_n823), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n890), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n841), .B1(G50), .B2(new_n1200), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n782), .A2(new_n567), .B1(new_n789), .B2(new_n881), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n987), .B1(new_n808), .B2(new_n268), .C1(new_n253), .C2(new_n814), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n664), .C2(new_n865), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n345), .B(new_n334), .C1(new_n801), .C2(new_n202), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT119), .Z(new_n1206));
  NAND2_X1  g1006(.A1(new_n779), .A2(G58), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT58), .ZN(new_n1209));
  AOI21_X1  g1009(.A(G50), .B1(new_n258), .B2(new_n345), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n411), .B2(G41), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n796), .A2(G125), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n814), .B2(new_n874), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n864), .A2(G128), .B1(new_n865), .B2(G137), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n801), .B2(new_n1167), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(G150), .C2(new_n794), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G33), .B(G41), .C1(new_n790), .C2(G124), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT59), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1219), .B1(new_n806), .B2(new_n778), .C1(new_n1216), .C2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1209), .B(new_n1211), .C1(new_n1218), .C2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1201), .B1(new_n1222), .B2(new_n821), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1199), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n936), .A2(G330), .A3(new_n948), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1193), .A2(new_n1198), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1229), .A2(G330), .A3(new_n936), .A4(new_n948), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n974), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n974), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1225), .B1(new_n1235), .B2(new_n840), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1149), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1232), .A2(new_n1234), .B1(new_n1161), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n737), .B1(new_n1239), .B2(KEYINPUT57), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT121), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1232), .A2(new_n1242), .A3(new_n1234), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT57), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1161), .B2(new_n1238), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1233), .A2(new_n1228), .A3(new_n1230), .A4(KEYINPUT121), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1237), .B1(new_n1241), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(G375));
  NAND3_X1  g1049(.A1(new_n1153), .A2(new_n1157), .A3(new_n1149), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1159), .A2(new_n1046), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n839), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n959), .A2(new_n823), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n841), .B1(G68), .B2(new_n1200), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n782), .A2(new_n881), .B1(new_n789), .B2(new_n883), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n411), .B(new_n1255), .C1(G107), .C2(new_n865), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n664), .A2(new_n794), .B1(new_n796), .B2(G294), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n799), .A2(G116), .B1(new_n802), .B2(G97), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1256), .A2(new_n994), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n411), .B1(new_n786), .B2(new_n868), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G137), .B2(new_n864), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n794), .A2(G50), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1167), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G132), .A2(new_n796), .B1(new_n799), .B2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1207), .A2(new_n1261), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n801), .A2(new_n806), .B1(new_n789), .B2(new_n1164), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT122), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1259), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1254), .B1(new_n1268), .B2(new_n821), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1252), .B1(new_n1253), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1251), .A2(new_n1270), .ZN(G381));
  NAND3_X1  g1071(.A1(new_n1065), .A2(new_n850), .A3(new_n1099), .ZN(new_n1272));
  OR3_X1    g1072(.A1(new_n1272), .A2(G384), .A3(G381), .ZN(new_n1273));
  NOR4_X1   g1073(.A1(new_n1273), .A2(G387), .A3(G390), .A4(G378), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1248), .B(KEYINPUT123), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1276), .B(KEYINPUT124), .Z(G407));
  INV_X1    g1077(.A(G213), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(G343), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(G378), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1278), .B1(new_n1275), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G407), .A2(new_n1282), .ZN(G409));
  NAND2_X1  g1083(.A1(G393), .A2(G396), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1272), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT126), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1284), .A2(new_n1287), .A3(new_n1272), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(G387), .A2(new_n1103), .A3(new_n1127), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G390), .B(new_n1013), .C1(new_n1047), .C2(new_n1058), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1289), .A2(KEYINPUT127), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1289), .A2(new_n1295), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT60), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1250), .B1(new_n1158), .B2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1153), .A2(new_n1157), .A3(new_n1149), .A4(KEYINPUT60), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n737), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1270), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(new_n892), .A3(new_n863), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(G384), .A2(new_n1270), .A3(new_n1302), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1279), .A2(G2897), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1306), .B(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1225), .B1(new_n1239), .B2(new_n1046), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1243), .A2(new_n840), .A3(new_n1246), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G378), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1243), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G378), .B(new_n1236), .C1(new_n1240), .C2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1247), .B(new_n737), .C1(KEYINPUT57), .C2(new_n1239), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1316), .A2(KEYINPUT125), .A3(G378), .A4(new_n1236), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1311), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1308), .B1(new_n1318), .B2(new_n1279), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1318), .A2(new_n1279), .A3(new_n1306), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1298), .B(new_n1319), .C1(new_n1320), .C2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1315), .A2(new_n1317), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1311), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1280), .ZN(new_n1326));
  NOR3_X1   g1126(.A1(new_n1326), .A2(KEYINPUT62), .A3(new_n1306), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1297), .B1(new_n1322), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1326), .B2(new_n1306), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT61), .B1(new_n1326), .B2(new_n1308), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1289), .A2(new_n1295), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1292), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1320), .A2(KEYINPUT63), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1330), .A2(new_n1331), .A3(new_n1335), .A4(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1328), .A2(new_n1337), .ZN(G405));
  OAI21_X1  g1138(.A(new_n1323), .B1(G378), .B2(new_n1248), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1306), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1297), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1343), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1335), .B1(new_n1345), .B2(new_n1341), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1344), .A2(new_n1346), .ZN(G402));
endmodule


