

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762;

  INV_X1 U379 ( .A(G953), .ZN(n754) );
  NOR2_X2 U380 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X2 U381 ( .A(n746), .B(n373), .ZN(n725) );
  XNOR2_X2 U382 ( .A(n407), .B(G122), .ZN(n511) );
  XOR2_X2 U383 ( .A(KEYINPUT38), .B(n611), .Z(n702) );
  INV_X1 U384 ( .A(n664), .ZN(n667) );
  NAND2_X1 U385 ( .A1(n667), .A2(n670), .ZN(n601) );
  NOR2_X1 U386 ( .A1(n588), .A2(n587), .ZN(n589) );
  INV_X1 U387 ( .A(n577), .ZN(n691) );
  NAND2_X1 U388 ( .A1(n534), .A2(n684), .ZN(n372) );
  INV_X1 U389 ( .A(G104), .ZN(n407) );
  NOR2_X1 U390 ( .A1(n635), .A2(n732), .ZN(n637) );
  NOR2_X1 U391 ( .A1(n631), .A2(n732), .ZN(n632) );
  AND2_X1 U392 ( .A1(n680), .A2(n405), .ZN(n404) );
  XNOR2_X1 U393 ( .A(n584), .B(KEYINPUT39), .ZN(n385) );
  XNOR2_X1 U394 ( .A(n581), .B(KEYINPUT42), .ZN(n762) );
  NOR2_X1 U395 ( .A1(n600), .A2(n700), .ZN(n581) );
  XNOR2_X1 U396 ( .A(n477), .B(KEYINPUT33), .ZN(n682) );
  AND2_X1 U397 ( .A1(n417), .A2(n359), .ZN(n415) );
  AND2_X1 U398 ( .A1(n574), .A2(n357), .ZN(n576) );
  OR2_X1 U399 ( .A1(n642), .A2(G902), .ZN(n427) );
  XNOR2_X1 U400 ( .A(n466), .B(n465), .ZN(n574) );
  AND2_X1 U401 ( .A1(n424), .A2(n423), .ZN(n422) );
  OR2_X1 U402 ( .A1(n633), .A2(G902), .ZN(n531) );
  XNOR2_X1 U403 ( .A(n481), .B(G131), .ZN(n376) );
  XNOR2_X1 U404 ( .A(n386), .B(KEYINPUT71), .ZN(n504) );
  XNOR2_X1 U405 ( .A(n437), .B(G146), .ZN(n481) );
  XNOR2_X1 U406 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n437) );
  XNOR2_X1 U407 ( .A(G902), .B(KEYINPUT15), .ZN(n616) );
  NOR2_X2 U408 ( .A1(n722), .A2(G953), .ZN(n723) );
  AND2_X2 U409 ( .A1(n551), .A2(n760), .ZN(n567) );
  OR2_X2 U410 ( .A1(n760), .A2(KEYINPUT81), .ZN(n361) );
  XNOR2_X2 U411 ( .A(n382), .B(n533), .ZN(n760) );
  XNOR2_X2 U412 ( .A(n367), .B(KEYINPUT72), .ZN(n681) );
  NAND2_X1 U413 ( .A1(n399), .A2(n370), .ZN(n398) );
  INV_X1 U414 ( .A(n762), .ZN(n370) );
  NAND2_X1 U415 ( .A1(n402), .A2(n607), .ZN(n401) );
  XNOR2_X1 U416 ( .A(n673), .B(KEYINPUT80), .ZN(n402) );
  NAND2_X1 U417 ( .A1(n701), .A2(KEYINPUT19), .ZN(n416) );
  NAND2_X1 U418 ( .A1(n388), .A2(n387), .ZN(n386) );
  INV_X1 U419 ( .A(G953), .ZN(n388) );
  INV_X1 U420 ( .A(G134), .ZN(n436) );
  NAND2_X1 U421 ( .A1(n421), .A2(n616), .ZN(n420) );
  INV_X1 U422 ( .A(n492), .ZN(n421) );
  NAND2_X1 U423 ( .A1(n490), .A2(n492), .ZN(n423) );
  XNOR2_X1 U424 ( .A(G101), .B(KEYINPUT3), .ZN(n471) );
  INV_X1 U425 ( .A(G119), .ZN(n469) );
  NAND2_X1 U426 ( .A1(n361), .A2(n355), .ZN(n369) );
  INV_X1 U427 ( .A(G146), .ZN(n512) );
  XNOR2_X1 U428 ( .A(n395), .B(n394), .ZN(n615) );
  INV_X1 U429 ( .A(KEYINPUT48), .ZN(n394) );
  XNOR2_X1 U430 ( .A(n398), .B(n397), .ZN(n396) );
  XNOR2_X1 U431 ( .A(n393), .B(n392), .ZN(n391) );
  XNOR2_X1 U432 ( .A(KEYINPUT99), .B(KEYINPUT30), .ZN(n392) );
  NAND2_X1 U433 ( .A1(n691), .A2(n701), .ZN(n393) );
  NAND2_X1 U434 ( .A1(n414), .A2(n413), .ZN(n412) );
  INV_X1 U435 ( .A(G469), .ZN(n442) );
  INV_X1 U436 ( .A(KEYINPUT6), .ZN(n426) );
  XNOR2_X1 U437 ( .A(n746), .B(n474), .ZN(n642) );
  XOR2_X1 U438 ( .A(KEYINPUT5), .B(G137), .Z(n467) );
  AND2_X1 U439 ( .A1(n615), .A2(n614), .ZN(n381) );
  INV_X1 U440 ( .A(G140), .ZN(n439) );
  XNOR2_X1 U441 ( .A(G104), .B(G101), .ZN(n440) );
  XNOR2_X1 U442 ( .A(KEYINPUT18), .B(G125), .ZN(n479) );
  NAND2_X1 U443 ( .A1(n428), .A2(n685), .ZN(n431) );
  NAND2_X1 U444 ( .A1(n591), .A2(KEYINPUT36), .ZN(n428) );
  XNOR2_X1 U445 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U446 ( .A(n488), .B(n487), .ZN(n741) );
  XOR2_X1 U447 ( .A(KEYINPUT90), .B(KEYINPUT11), .Z(n507) );
  INV_X1 U448 ( .A(KEYINPUT46), .ZN(n397) );
  INV_X1 U449 ( .A(G902), .ZN(n491) );
  XNOR2_X1 U450 ( .A(n555), .B(KEYINPUT1), .ZN(n534) );
  XNOR2_X1 U451 ( .A(G125), .B(KEYINPUT10), .ZN(n457) );
  NAND2_X1 U452 ( .A1(G234), .A2(G237), .ZN(n495) );
  XNOR2_X1 U453 ( .A(G146), .B(G128), .ZN(n451) );
  XNOR2_X1 U454 ( .A(G122), .B(G116), .ZN(n522) );
  XOR2_X1 U455 ( .A(KEYINPUT9), .B(G107), .Z(n523) );
  XNOR2_X1 U456 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U457 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U458 ( .A1(n378), .A2(n377), .ZN(n625) );
  NAND2_X1 U459 ( .A1(n490), .A2(KEYINPUT2), .ZN(n377) );
  NAND2_X1 U460 ( .A1(n735), .A2(n379), .ZN(n378) );
  AND2_X1 U461 ( .A1(n381), .A2(n490), .ZN(n379) );
  XNOR2_X1 U462 ( .A(n679), .B(n406), .ZN(n405) );
  NOR2_X1 U463 ( .A1(n381), .A2(KEYINPUT2), .ZN(n679) );
  XNOR2_X1 U464 ( .A(n371), .B(n365), .ZN(n700) );
  NOR2_X1 U465 ( .A1(n704), .A2(n705), .ZN(n371) );
  XNOR2_X1 U466 ( .A(n582), .B(n390), .ZN(n389) );
  INV_X1 U467 ( .A(KEYINPUT98), .ZN(n390) );
  AND2_X1 U468 ( .A1(n412), .A2(n410), .ZN(n409) );
  NOR2_X1 U469 ( .A1(G902), .A2(n731), .ZN(n466) );
  AND2_X2 U470 ( .A1(n681), .A2(n625), .ZN(n729) );
  XNOR2_X1 U471 ( .A(n375), .B(n374), .ZN(n373) );
  XNOR2_X1 U472 ( .A(n485), .B(n362), .ZN(n374) );
  XNOR2_X1 U473 ( .A(n441), .B(n458), .ZN(n375) );
  XNOR2_X1 U474 ( .A(n741), .B(n489), .ZN(n628) );
  NOR2_X1 U475 ( .A1(n754), .A2(G952), .ZN(n732) );
  NOR2_X1 U476 ( .A1(n685), .A2(n609), .ZN(n610) );
  XNOR2_X1 U477 ( .A(n586), .B(n585), .ZN(n759) );
  NAND2_X1 U478 ( .A1(n385), .A2(n664), .ZN(n586) );
  OR2_X1 U479 ( .A1(n432), .A2(n591), .ZN(n429) );
  AND2_X1 U480 ( .A1(n548), .A2(n639), .ZN(n355) );
  AND2_X1 U481 ( .A1(n433), .A2(KEYINPUT36), .ZN(n356) );
  OR2_X1 U482 ( .A1(n573), .A2(n572), .ZN(n357) );
  AND2_X1 U483 ( .A1(n614), .A2(KEYINPUT2), .ZN(n358) );
  OR2_X1 U484 ( .A1(n422), .A2(n416), .ZN(n359) );
  AND2_X1 U485 ( .A1(n391), .A2(n357), .ZN(n360) );
  AND2_X1 U486 ( .A1(G227), .A2(n754), .ZN(n362) );
  AND2_X1 U487 ( .A1(n577), .A2(n574), .ZN(n363) );
  AND2_X1 U488 ( .A1(n611), .A2(n435), .ZN(n364) );
  INV_X1 U489 ( .A(G237), .ZN(n387) );
  XNOR2_X1 U490 ( .A(KEYINPUT102), .B(KEYINPUT41), .ZN(n365) );
  INV_X1 U491 ( .A(KEYINPUT36), .ZN(n435) );
  OR2_X1 U492 ( .A1(KEYINPUT81), .A2(KEYINPUT44), .ZN(n366) );
  NAND2_X1 U493 ( .A1(n380), .A2(n735), .ZN(n367) );
  NAND2_X1 U494 ( .A1(n556), .A2(n538), .ZN(n541) );
  XNOR2_X2 U495 ( .A(n502), .B(n501), .ZN(n556) );
  NAND2_X1 U496 ( .A1(n368), .A2(n363), .ZN(n639) );
  XNOR2_X1 U497 ( .A(n564), .B(KEYINPUT94), .ZN(n368) );
  NOR2_X2 U498 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U499 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U500 ( .A1(n369), .A2(n366), .ZN(n569) );
  AND2_X2 U501 ( .A1(n547), .A2(n592), .ZN(n564) );
  NAND2_X1 U502 ( .A1(n549), .A2(n639), .ZN(n408) );
  NAND2_X1 U503 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U504 ( .A1(n401), .A2(n598), .ZN(n400) );
  NOR2_X1 U505 ( .A1(n356), .A2(n431), .ZN(n430) );
  NAND2_X1 U506 ( .A1(n434), .A2(n664), .ZN(n608) );
  XNOR2_X1 U507 ( .A(n552), .B(KEYINPUT95), .ZN(n476) );
  XNOR2_X2 U508 ( .A(n372), .B(KEYINPUT70), .ZN(n552) );
  XNOR2_X2 U509 ( .A(n376), .B(n525), .ZN(n746) );
  XNOR2_X2 U510 ( .A(n482), .B(n436), .ZN(n525) );
  XNOR2_X2 U511 ( .A(n425), .B(KEYINPUT65), .ZN(n482) );
  XNOR2_X1 U512 ( .A(n617), .B(KEYINPUT79), .ZN(n380) );
  XNOR2_X2 U513 ( .A(n570), .B(KEYINPUT45), .ZN(n735) );
  NAND2_X1 U514 ( .A1(n383), .A2(n532), .ZN(n382) );
  XNOR2_X1 U515 ( .A(n503), .B(n384), .ZN(n383) );
  INV_X1 U516 ( .A(KEYINPUT34), .ZN(n384) );
  NAND2_X1 U517 ( .A1(n385), .A2(n658), .ZN(n677) );
  NAND2_X1 U518 ( .A1(n504), .A2(G210), .ZN(n468) );
  NAND2_X1 U519 ( .A1(n360), .A2(n389), .ZN(n594) );
  NAND2_X1 U520 ( .A1(n684), .A2(n555), .ZN(n582) );
  NAND2_X1 U521 ( .A1(n400), .A2(n396), .ZN(n395) );
  INV_X1 U522 ( .A(n759), .ZN(n399) );
  NAND2_X1 U523 ( .A1(n403), .A2(n683), .ZN(n720) );
  NAND2_X1 U524 ( .A1(n404), .A2(n681), .ZN(n403) );
  INV_X1 U525 ( .A(KEYINPUT78), .ZN(n406) );
  NAND2_X1 U526 ( .A1(n408), .A2(n550), .ZN(n551) );
  NAND2_X1 U527 ( .A1(n422), .A2(n419), .ZN(n611) );
  NAND2_X1 U528 ( .A1(n415), .A2(n409), .ZN(n599) );
  NAND2_X1 U529 ( .A1(n411), .A2(n494), .ZN(n410) );
  INV_X1 U530 ( .A(n701), .ZN(n411) );
  INV_X1 U531 ( .A(n416), .ZN(n413) );
  INV_X1 U532 ( .A(n419), .ZN(n414) );
  NAND2_X1 U533 ( .A1(n418), .A2(n422), .ZN(n417) );
  AND2_X1 U534 ( .A1(n419), .A2(n494), .ZN(n418) );
  OR2_X1 U535 ( .A1(n628), .A2(n420), .ZN(n419) );
  NAND2_X1 U536 ( .A1(n628), .A2(n492), .ZN(n424) );
  XNOR2_X2 U537 ( .A(G143), .B(G128), .ZN(n425) );
  XNOR2_X1 U538 ( .A(n577), .B(n426), .ZN(n588) );
  XNOR2_X2 U539 ( .A(n427), .B(n475), .ZN(n577) );
  NAND2_X1 U540 ( .A1(n615), .A2(n358), .ZN(n617) );
  NAND2_X1 U541 ( .A1(n664), .A2(n611), .ZN(n433) );
  NAND2_X1 U542 ( .A1(n430), .A2(n429), .ZN(n673) );
  NAND2_X1 U543 ( .A1(n664), .A2(n364), .ZN(n432) );
  INV_X1 U544 ( .A(n591), .ZN(n434) );
  NOR2_X1 U545 ( .A1(n735), .A2(KEYINPUT2), .ZN(n678) );
  INV_X1 U546 ( .A(n677), .ZN(n613) );
  NOR2_X1 U547 ( .A1(n638), .A2(n613), .ZN(n614) );
  XNOR2_X1 U548 ( .A(n450), .B(n449), .ZN(n453) );
  XNOR2_X1 U549 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U550 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U551 ( .A(n442), .B(KEYINPUT68), .ZN(n443) );
  XNOR2_X1 U552 ( .A(n453), .B(n452), .ZN(n456) );
  XNOR2_X1 U553 ( .A(n484), .B(n483), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n462), .B(KEYINPUT86), .ZN(n464) );
  XNOR2_X1 U555 ( .A(n464), .B(n463), .ZN(n465) );
  AND2_X1 U556 ( .A1(n729), .A2(G472), .ZN(n644) );
  XNOR2_X1 U557 ( .A(n521), .B(n520), .ZN(n560) );
  XNOR2_X1 U558 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U559 ( .A(KEYINPUT101), .B(KEYINPUT40), .ZN(n585) );
  XOR2_X1 U560 ( .A(G137), .B(KEYINPUT67), .Z(n458) );
  INV_X1 U561 ( .A(G110), .ZN(n438) );
  XNOR2_X1 U562 ( .A(n438), .B(G107), .ZN(n485) );
  NOR2_X2 U563 ( .A1(G902), .A2(n725), .ZN(n444) );
  XNOR2_X2 U564 ( .A(n444), .B(n443), .ZN(n555) );
  NAND2_X1 U565 ( .A1(G234), .A2(n616), .ZN(n445) );
  XNOR2_X1 U566 ( .A(KEYINPUT20), .B(n445), .ZN(n461) );
  AND2_X1 U567 ( .A1(n461), .A2(G221), .ZN(n448) );
  INV_X1 U568 ( .A(KEYINPUT87), .ZN(n446) );
  XNOR2_X1 U569 ( .A(n446), .B(KEYINPUT21), .ZN(n447) );
  XNOR2_X1 U570 ( .A(n448), .B(n447), .ZN(n575) );
  INV_X1 U571 ( .A(n575), .ZN(n688) );
  XOR2_X1 U572 ( .A(G119), .B(G110), .Z(n450) );
  XOR2_X1 U573 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n449) );
  XNOR2_X1 U574 ( .A(n451), .B(KEYINPUT85), .ZN(n452) );
  NAND2_X1 U575 ( .A1(G234), .A2(n754), .ZN(n454) );
  XOR2_X1 U576 ( .A(KEYINPUT8), .B(n454), .Z(n526) );
  NAND2_X1 U577 ( .A1(n526), .A2(G221), .ZN(n455) );
  XNOR2_X1 U578 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X1 U579 ( .A(n457), .B(G140), .ZN(n505) );
  INV_X1 U580 ( .A(n458), .ZN(n459) );
  XNOR2_X1 U581 ( .A(n505), .B(n459), .ZN(n745) );
  XNOR2_X1 U582 ( .A(n460), .B(n745), .ZN(n731) );
  NAND2_X1 U583 ( .A1(n461), .A2(G217), .ZN(n462) );
  XNOR2_X1 U584 ( .A(KEYINPUT25), .B(KEYINPUT73), .ZN(n463) );
  NOR2_X1 U585 ( .A1(n688), .A2(n574), .ZN(n684) );
  XNOR2_X1 U586 ( .A(n468), .B(n467), .ZN(n473) );
  XNOR2_X1 U587 ( .A(G116), .B(G113), .ZN(n470) );
  XNOR2_X1 U588 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U589 ( .A(n472), .B(n471), .ZN(n487) );
  XNOR2_X1 U590 ( .A(n473), .B(n487), .ZN(n474) );
  INV_X1 U591 ( .A(G472), .ZN(n475) );
  INV_X1 U592 ( .A(n588), .ZN(n562) );
  NAND2_X1 U593 ( .A1(n476), .A2(n562), .ZN(n477) );
  NAND2_X1 U594 ( .A1(n754), .A2(G224), .ZN(n478) );
  XNOR2_X1 U595 ( .A(n478), .B(KEYINPUT17), .ZN(n480) );
  XNOR2_X1 U596 ( .A(n480), .B(n479), .ZN(n484) );
  XNOR2_X1 U597 ( .A(n511), .B(KEYINPUT16), .ZN(n486) );
  XNOR2_X1 U598 ( .A(n486), .B(n485), .ZN(n488) );
  INV_X1 U599 ( .A(n616), .ZN(n490) );
  NAND2_X1 U600 ( .A1(n491), .A2(n387), .ZN(n493) );
  AND2_X1 U601 ( .A1(n493), .A2(G210), .ZN(n492) );
  NAND2_X1 U602 ( .A1(n493), .A2(G214), .ZN(n701) );
  INV_X1 U603 ( .A(KEYINPUT19), .ZN(n494) );
  XNOR2_X1 U604 ( .A(n495), .B(KEYINPUT14), .ZN(n498) );
  NAND2_X1 U605 ( .A1(G902), .A2(n498), .ZN(n496) );
  XOR2_X1 U606 ( .A(KEYINPUT84), .B(n496), .Z(n497) );
  NAND2_X1 U607 ( .A1(G953), .A2(n497), .ZN(n571) );
  NOR2_X1 U608 ( .A1(n571), .A2(G898), .ZN(n499) );
  NAND2_X1 U609 ( .A1(n498), .A2(G952), .ZN(n717) );
  NOR2_X1 U610 ( .A1(n717), .A2(G953), .ZN(n573) );
  NOR2_X1 U611 ( .A1(n499), .A2(n573), .ZN(n500) );
  OR2_X2 U612 ( .A1(n599), .A2(n500), .ZN(n502) );
  INV_X1 U613 ( .A(KEYINPUT0), .ZN(n501) );
  NAND2_X1 U614 ( .A1(n682), .A2(n556), .ZN(n503) );
  NAND2_X1 U615 ( .A1(n504), .A2(G214), .ZN(n517) );
  XOR2_X1 U616 ( .A(n505), .B(G131), .Z(n510) );
  XNOR2_X1 U617 ( .A(G143), .B(KEYINPUT89), .ZN(n506) );
  XNOR2_X1 U618 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U619 ( .A(n508), .B(KEYINPUT12), .ZN(n509) );
  XNOR2_X1 U620 ( .A(n510), .B(n509), .ZN(n515) );
  XNOR2_X1 U621 ( .A(n511), .B(G113), .ZN(n513) );
  XNOR2_X1 U622 ( .A(n517), .B(n516), .ZN(n619) );
  NOR2_X1 U623 ( .A1(G902), .A2(n619), .ZN(n521) );
  XNOR2_X1 U624 ( .A(KEYINPUT91), .B(KEYINPUT13), .ZN(n519) );
  INV_X1 U625 ( .A(G475), .ZN(n518) );
  XNOR2_X1 U626 ( .A(KEYINPUT92), .B(KEYINPUT7), .ZN(n530) );
  XNOR2_X1 U627 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U628 ( .A(n525), .B(n524), .Z(n528) );
  NAND2_X1 U629 ( .A1(G217), .A2(n526), .ZN(n527) );
  XNOR2_X1 U630 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U631 ( .A(n530), .B(n529), .ZN(n633) );
  XNOR2_X1 U632 ( .A(G478), .B(n531), .ZN(n558) );
  NAND2_X1 U633 ( .A1(n560), .A2(n558), .ZN(n597) );
  INV_X1 U634 ( .A(n597), .ZN(n532) );
  INV_X1 U635 ( .A(KEYINPUT35), .ZN(n533) );
  INV_X1 U636 ( .A(n534), .ZN(n592) );
  INV_X1 U637 ( .A(n592), .ZN(n685) );
  INV_X1 U638 ( .A(KEYINPUT93), .ZN(n535) );
  XNOR2_X1 U639 ( .A(n574), .B(n535), .ZN(n687) );
  NAND2_X1 U640 ( .A1(n685), .A2(n687), .ZN(n536) );
  NOR2_X1 U641 ( .A1(n562), .A2(n536), .ZN(n537) );
  XOR2_X1 U642 ( .A(KEYINPUT74), .B(n537), .Z(n542) );
  NOR2_X1 U643 ( .A1(n560), .A2(n558), .ZN(n580) );
  AND2_X1 U644 ( .A1(n580), .A2(n575), .ZN(n538) );
  INV_X1 U645 ( .A(KEYINPUT69), .ZN(n539) );
  XNOR2_X1 U646 ( .A(n539), .B(KEYINPUT22), .ZN(n540) );
  XNOR2_X1 U647 ( .A(n541), .B(n540), .ZN(n546) );
  NOR2_X1 U648 ( .A1(n542), .A2(n546), .ZN(n544) );
  XNOR2_X1 U649 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n543) );
  XNOR2_X1 U650 ( .A(n544), .B(n543), .ZN(n761) );
  INV_X1 U651 ( .A(KEYINPUT44), .ZN(n545) );
  NOR2_X1 U652 ( .A1(n761), .A2(n545), .ZN(n548) );
  INV_X1 U653 ( .A(n546), .ZN(n547) );
  NOR2_X1 U654 ( .A1(n761), .A2(KEYINPUT44), .ZN(n549) );
  INV_X1 U655 ( .A(KEYINPUT81), .ZN(n550) );
  NOR2_X1 U656 ( .A1(n552), .A2(n577), .ZN(n694) );
  NAND2_X1 U657 ( .A1(n694), .A2(n556), .ZN(n554) );
  XOR2_X1 U658 ( .A(KEYINPUT88), .B(KEYINPUT31), .Z(n553) );
  XNOR2_X1 U659 ( .A(n554), .B(n553), .ZN(n671) );
  NOR2_X1 U660 ( .A1(n582), .A2(n691), .ZN(n557) );
  NAND2_X1 U661 ( .A1(n557), .A2(n556), .ZN(n653) );
  NAND2_X1 U662 ( .A1(n671), .A2(n653), .ZN(n561) );
  INV_X1 U663 ( .A(n558), .ZN(n559) );
  AND2_X1 U664 ( .A1(n560), .A2(n559), .ZN(n664) );
  NOR2_X1 U665 ( .A1(n560), .A2(n559), .ZN(n658) );
  INV_X1 U666 ( .A(n658), .ZN(n670) );
  NAND2_X1 U667 ( .A1(n561), .A2(n601), .ZN(n565) );
  NOR2_X1 U668 ( .A1(n562), .A2(n687), .ZN(n563) );
  NAND2_X1 U669 ( .A1(n564), .A2(n563), .ZN(n648) );
  NAND2_X1 U670 ( .A1(n565), .A2(n648), .ZN(n566) );
  NOR2_X1 U671 ( .A1(G900), .A2(n571), .ZN(n572) );
  NAND2_X1 U672 ( .A1(n576), .A2(n575), .ZN(n587) );
  NOR2_X1 U673 ( .A1(n577), .A2(n587), .ZN(n578) );
  XNOR2_X1 U674 ( .A(n578), .B(KEYINPUT28), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n579), .A2(n555), .ZN(n600) );
  INV_X1 U676 ( .A(n580), .ZN(n704) );
  NAND2_X1 U677 ( .A1(n702), .A2(n701), .ZN(n705) );
  INV_X1 U678 ( .A(n594), .ZN(n583) );
  NAND2_X1 U679 ( .A1(n702), .A2(n583), .ZN(n584) );
  XNOR2_X1 U680 ( .A(n589), .B(KEYINPUT96), .ZN(n590) );
  NAND2_X1 U681 ( .A1(n590), .A2(n701), .ZN(n591) );
  INV_X1 U682 ( .A(n611), .ZN(n593) );
  NOR2_X1 U683 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U684 ( .A(KEYINPUT100), .B(n595), .Z(n596) );
  NOR2_X1 U685 ( .A1(n597), .A2(n596), .ZN(n662) );
  XNOR2_X1 U686 ( .A(KEYINPUT76), .B(n662), .ZN(n598) );
  NOR2_X1 U687 ( .A1(n600), .A2(n599), .ZN(n665) );
  XOR2_X1 U688 ( .A(KEYINPUT47), .B(n665), .Z(n603) );
  INV_X1 U689 ( .A(n601), .ZN(n706) );
  NAND2_X1 U690 ( .A1(n665), .A2(n706), .ZN(n602) );
  NAND2_X1 U691 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n706), .A2(KEYINPUT47), .ZN(n604) );
  XOR2_X1 U693 ( .A(KEYINPUT75), .B(n604), .Z(n605) );
  AND2_X1 U694 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U695 ( .A(KEYINPUT97), .B(n608), .Z(n609) );
  XNOR2_X1 U696 ( .A(n610), .B(KEYINPUT43), .ZN(n612) );
  NOR2_X1 U697 ( .A1(n612), .A2(n611), .ZN(n638) );
  AND2_X1 U698 ( .A1(n625), .A2(G475), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n618), .A2(n681), .ZN(n621) );
  XOR2_X1 U700 ( .A(n619), .B(KEYINPUT59), .Z(n620) );
  XNOR2_X1 U701 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X1 U702 ( .A1(n622), .A2(n732), .ZN(n624) );
  XNOR2_X1 U703 ( .A(KEYINPUT118), .B(KEYINPUT60), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n624), .B(n623), .ZN(G60) );
  NAND2_X1 U705 ( .A1(n729), .A2(G210), .ZN(n630) );
  XOR2_X1 U706 ( .A(KEYINPUT82), .B(KEYINPUT55), .Z(n626) );
  XNOR2_X1 U707 ( .A(n626), .B(KEYINPUT54), .ZN(n627) );
  XNOR2_X1 U708 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U709 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n632), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U711 ( .A1(n729), .A2(G478), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n634), .B(n633), .ZN(n635) );
  INV_X1 U713 ( .A(KEYINPUT119), .ZN(n636) );
  XNOR2_X1 U714 ( .A(n637), .B(n636), .ZN(G63) );
  XOR2_X1 U715 ( .A(G140), .B(n638), .Z(G42) );
  XNOR2_X1 U716 ( .A(n639), .B(G110), .ZN(G12) );
  XNOR2_X1 U717 ( .A(KEYINPUT83), .B(KEYINPUT103), .ZN(n640) );
  XOR2_X1 U718 ( .A(n640), .B(KEYINPUT62), .Z(n641) );
  XNOR2_X1 U719 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X1 U721 ( .A1(n645), .A2(n732), .ZN(n647) );
  XOR2_X1 U722 ( .A(KEYINPUT104), .B(KEYINPUT63), .Z(n646) );
  XNOR2_X1 U723 ( .A(n647), .B(n646), .ZN(G57) );
  XNOR2_X1 U724 ( .A(G101), .B(n648), .ZN(G3) );
  NOR2_X1 U725 ( .A1(n653), .A2(n667), .ZN(n650) );
  XNOR2_X1 U726 ( .A(G104), .B(KEYINPUT105), .ZN(n649) );
  XNOR2_X1 U727 ( .A(n650), .B(n649), .ZN(G6) );
  XOR2_X1 U728 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n652) );
  XNOR2_X1 U729 ( .A(KEYINPUT106), .B(KEYINPUT27), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n652), .B(n651), .ZN(n657) );
  NOR2_X1 U731 ( .A1(n653), .A2(n670), .ZN(n655) );
  XNOR2_X1 U732 ( .A(G107), .B(KEYINPUT26), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U734 ( .A(n657), .B(n656), .ZN(G9) );
  XOR2_X1 U735 ( .A(KEYINPUT109), .B(KEYINPUT29), .Z(n660) );
  NAND2_X1 U736 ( .A1(n665), .A2(n658), .ZN(n659) );
  XNOR2_X1 U737 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X1 U738 ( .A(G128), .B(n661), .Z(G30) );
  XOR2_X1 U739 ( .A(G143), .B(n662), .Z(n663) );
  XNOR2_X1 U740 ( .A(KEYINPUT110), .B(n663), .ZN(G45) );
  NAND2_X1 U741 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n666), .B(G146), .ZN(G48) );
  NOR2_X1 U743 ( .A1(n671), .A2(n667), .ZN(n669) );
  XNOR2_X1 U744 ( .A(G113), .B(KEYINPUT111), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n669), .B(n668), .ZN(G15) );
  NOR2_X1 U746 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U747 ( .A(G116), .B(n672), .Z(G18) );
  INV_X1 U748 ( .A(n673), .ZN(n674) );
  XNOR2_X1 U749 ( .A(n674), .B(KEYINPUT37), .ZN(n675) );
  XNOR2_X1 U750 ( .A(n675), .B(KEYINPUT112), .ZN(n676) );
  XNOR2_X1 U751 ( .A(G125), .B(n676), .ZN(G27) );
  XNOR2_X1 U752 ( .A(G134), .B(n677), .ZN(G36) );
  XNOR2_X1 U753 ( .A(n678), .B(KEYINPUT77), .ZN(n680) );
  INV_X1 U754 ( .A(n682), .ZN(n710) );
  OR2_X1 U755 ( .A1(n710), .A2(n700), .ZN(n683) );
  XOR2_X1 U756 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n716) );
  OR2_X1 U757 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n686), .B(KEYINPUT50), .ZN(n693) );
  NAND2_X1 U759 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U760 ( .A(KEYINPUT49), .B(n689), .ZN(n690) );
  NOR2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n696) );
  INV_X1 U763 ( .A(n694), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U765 ( .A(n697), .B(KEYINPUT51), .Z(n698) );
  XNOR2_X1 U766 ( .A(KEYINPUT113), .B(n698), .ZN(n699) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U773 ( .A(n711), .B(KEYINPUT114), .ZN(n712) );
  NOR2_X1 U774 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U775 ( .A(n714), .B(KEYINPUT52), .ZN(n715) );
  XNOR2_X1 U776 ( .A(n716), .B(n715), .ZN(n718) );
  NOR2_X1 U777 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U778 ( .A(n721), .B(KEYINPUT117), .ZN(n722) );
  XNOR2_X1 U779 ( .A(n723), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U780 ( .A1(n729), .A2(G469), .ZN(n727) );
  XOR2_X1 U781 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n724) );
  XNOR2_X1 U782 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U783 ( .A1(n732), .A2(n728), .ZN(G54) );
  NAND2_X1 U784 ( .A1(n729), .A2(G217), .ZN(n730) );
  XNOR2_X1 U785 ( .A(n731), .B(n730), .ZN(n733) );
  XNOR2_X1 U786 ( .A(n734), .B(KEYINPUT120), .ZN(G66) );
  NAND2_X1 U787 ( .A1(n735), .A2(n754), .ZN(n739) );
  NAND2_X1 U788 ( .A1(G953), .A2(G224), .ZN(n736) );
  XNOR2_X1 U789 ( .A(KEYINPUT61), .B(n736), .ZN(n737) );
  NAND2_X1 U790 ( .A1(n737), .A2(G898), .ZN(n738) );
  NAND2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n744) );
  OR2_X1 U792 ( .A1(G898), .A2(n754), .ZN(n740) );
  NAND2_X1 U793 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U794 ( .A(n742), .B(KEYINPUT121), .ZN(n743) );
  XNOR2_X1 U795 ( .A(n744), .B(n743), .ZN(G69) );
  XNOR2_X1 U796 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U797 ( .A(n747), .B(KEYINPUT122), .ZN(n752) );
  XNOR2_X1 U798 ( .A(n752), .B(G227), .ZN(n748) );
  XNOR2_X1 U799 ( .A(n748), .B(KEYINPUT124), .ZN(n749) );
  NAND2_X1 U800 ( .A1(n749), .A2(G900), .ZN(n750) );
  NAND2_X1 U801 ( .A1(G953), .A2(n750), .ZN(n751) );
  XOR2_X1 U802 ( .A(KEYINPUT125), .B(n751), .Z(n757) );
  XNOR2_X1 U803 ( .A(n752), .B(n381), .ZN(n753) );
  XNOR2_X1 U804 ( .A(n753), .B(KEYINPUT123), .ZN(n755) );
  NAND2_X1 U805 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U806 ( .A1(n757), .A2(n756), .ZN(G72) );
  XOR2_X1 U807 ( .A(G131), .B(KEYINPUT126), .Z(n758) );
  XNOR2_X1 U808 ( .A(n759), .B(n758), .ZN(G33) );
  XNOR2_X1 U809 ( .A(n760), .B(G122), .ZN(G24) );
  XOR2_X1 U810 ( .A(G119), .B(n761), .Z(G21) );
  XOR2_X1 U811 ( .A(G137), .B(n762), .Z(G39) );
endmodule

