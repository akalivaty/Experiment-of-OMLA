//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  AND3_X1   g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G50gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G43gat), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT15), .B1(new_n213), .B2(G50gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n208), .B(new_n209), .C1(new_n212), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n213), .A2(G50gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n214), .B1(KEYINPUT87), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(KEYINPUT87), .B2(new_n221), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(new_n215), .A3(new_n208), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT88), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n220), .A2(KEYINPUT88), .A3(new_n224), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT16), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G1gat), .B2(new_n231), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(G8gat), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n225), .A2(KEYINPUT17), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n230), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n236), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n227), .A3(new_n229), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G169gat), .B(G197gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT12), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n227), .A2(new_n229), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n236), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n241), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n239), .B(KEYINPUT13), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n238), .A2(KEYINPUT18), .A3(new_n239), .A4(new_n241), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n244), .A2(new_n250), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n242), .A2(new_n243), .B1(new_n253), .B2(new_n254), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n250), .B1(new_n259), .B2(new_n256), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262));
  INV_X1    g061(.A(G134gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G127gat), .ZN(new_n264));
  INV_X1    g063(.A(G127gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G134gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G120gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G113gat), .ZN(new_n270));
  INV_X1    g069(.A(G113gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G113gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n274), .A3(G120gat), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n268), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(G120gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n278), .A2(new_n267), .B1(new_n264), .B2(new_n266), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n262), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n266), .ZN(new_n281));
  XNOR2_X1  g080(.A(G113gat), .B(G120gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(KEYINPUT1), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n271), .A2(G120gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT67), .B(G113gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n285), .B2(G120gat), .ZN(new_n286));
  OAI211_X1 g085(.A(KEYINPUT68), .B(new_n283), .C1(new_n286), .C2(new_n268), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  INV_X1    g088(.A(G190gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT66), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(G183gat), .B2(G190gat), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT24), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(G183gat), .A3(G190gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G169gat), .ZN(new_n301));
  INV_X1    g100(.A(G176gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT23), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT25), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n289), .A2(KEYINPUT27), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G183gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n311), .A3(new_n290), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n312), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(new_n301), .A3(new_n302), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(new_n306), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n309), .A2(new_n311), .A3(new_n318), .A4(new_n290), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n321), .B(new_n306), .C1(new_n322), .C2(KEYINPUT23), .ZN(new_n323));
  OR2_X1    g122(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n304), .A2(G169gat), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n289), .A2(new_n290), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n299), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n313), .A2(new_n320), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n288), .A2(new_n308), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n312), .A2(KEYINPUT28), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n333), .A2(new_n295), .A3(new_n319), .A4(new_n317), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n305), .A2(new_n306), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n327), .A2(new_n324), .A3(new_n325), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n330), .A2(new_n335), .A3(new_n321), .A4(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n307), .B1(new_n294), .B2(new_n299), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n334), .B(new_n337), .C1(new_n321), .C2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(new_n280), .A3(new_n287), .ZN(new_n340));
  NAND2_X1  g139(.A1(G227gat), .A2(G233gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n341), .B(KEYINPUT64), .Z(new_n342));
  NAND3_X1  g141(.A1(new_n332), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT32), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT33), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G15gat), .B(G43gat), .Z(new_n347));
  XNOR2_X1  g146(.A(G71gat), .B(G99gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n344), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n349), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n343), .B(KEYINPUT32), .C1(new_n345), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT34), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n340), .ZN(new_n355));
  INV_X1    g154(.A(new_n342), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI211_X1 g156(.A(KEYINPUT34), .B(new_n342), .C1(new_n332), .C2(new_n340), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n357), .A2(new_n358), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n350), .A3(new_n352), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n359), .A2(KEYINPUT36), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT36), .B1(new_n359), .B2(new_n361), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n365));
  INV_X1    g164(.A(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G141gat), .ZN(new_n367));
  INV_X1    g166(.A(G141gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G148gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT70), .B(KEYINPUT2), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G155gat), .ZN(new_n373));
  INV_X1    g172(.A(G162gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT71), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n368), .B2(G148gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n366), .A2(KEYINPUT71), .A3(G141gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n369), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n376), .B1(new_n375), .B2(KEYINPUT2), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n372), .A2(new_n377), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT29), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G211gat), .A2(G218gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT22), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(G197gat), .A2(G204gat), .ZN(new_n389));
  AND2_X1   g188(.A1(G197gat), .A2(G204gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G211gat), .B(G218gat), .Z(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G211gat), .B(G218gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G197gat), .B(G204gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n388), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n365), .B1(new_n385), .B2(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(KEYINPUT70), .B(KEYINPUT2), .Z(new_n399));
  XNOR2_X1  g198(.A(G141gat), .B(G148gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n377), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n382), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n384), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n397), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(KEYINPUT76), .A3(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n401), .A2(KEYINPUT72), .A3(new_n402), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT72), .B1(new_n401), .B2(new_n402), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n393), .B2(new_n396), .ZN(new_n410));
  OAI22_X1  g209(.A1(new_n408), .A2(new_n409), .B1(new_n410), .B2(KEYINPUT3), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n398), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G22gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n391), .A2(new_n392), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n394), .B1(new_n388), .B2(new_n395), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n404), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n383), .B1(new_n418), .B2(new_n384), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n419), .A2(new_n420), .A3(new_n413), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n414), .A2(new_n415), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n412), .B2(new_n413), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(new_n415), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT75), .B(KEYINPUT31), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(G50gat), .ZN(new_n428));
  XOR2_X1   g227(.A(G78gat), .B(G106gat), .Z(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n424), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n423), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT78), .ZN(new_n434));
  INV_X1    g233(.A(new_n413), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n405), .A2(new_n406), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT72), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n381), .A2(new_n382), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n375), .A2(new_n376), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n370), .B2(new_n371), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n401), .A2(KEYINPUT72), .A3(new_n402), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n418), .A2(new_n384), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n436), .A2(new_n365), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n435), .B1(new_n445), .B2(new_n407), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n434), .B(G22gat), .C1(new_n446), .C2(new_n421), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT78), .B1(new_n425), .B2(new_n415), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n425), .A2(KEYINPUT77), .A3(new_n415), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n433), .A2(new_n447), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n430), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT79), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n430), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n431), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G8gat), .B(G36gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(G64gat), .ZN(new_n457));
  INV_X1    g256(.A(G92gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(G226gat), .A2(G233gat), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n339), .B2(new_n404), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n331), .B2(new_n308), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n406), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n339), .A2(new_n461), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT29), .B1(new_n331), .B2(new_n308), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n465), .B(new_n397), .C1(new_n466), .C2(new_n461), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n459), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT69), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n464), .A2(new_n467), .A3(new_n459), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT30), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G225gat), .A2(G233gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n283), .B1(new_n286), .B2(new_n268), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n383), .B2(new_n384), .ZN(new_n476));
  INV_X1    g275(.A(new_n403), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(KEYINPUT5), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT4), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n401), .A2(new_n402), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT73), .B1(new_n481), .B2(new_n475), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n275), .A2(new_n270), .ZN(new_n483));
  INV_X1    g282(.A(new_n268), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n269), .A2(G113gat), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n267), .B1(new_n284), .B2(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n483), .A2(new_n484), .B1(new_n486), .B2(new_n281), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT73), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n383), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n480), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n441), .A2(new_n280), .A3(new_n442), .A4(new_n287), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n479), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n491), .A2(new_n480), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT4), .B1(new_n482), .B2(new_n489), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n494), .A2(new_n495), .A3(new_n478), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT74), .B1(new_n487), .B2(new_n383), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n475), .A3(new_n498), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n482), .A2(new_n489), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT5), .B1(new_n500), .B2(new_n474), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n493), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G1gat), .B(G29gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT0), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(G57gat), .ZN(new_n505));
  INV_X1    g304(.A(G85gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT6), .B1(new_n502), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n493), .B(new_n507), .C1(new_n496), .C2(new_n501), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n502), .A2(KEYINPUT6), .A3(new_n508), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n473), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n364), .B1(new_n455), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT80), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n476), .A2(new_n477), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n408), .A2(new_n409), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n518), .A2(new_n480), .A3(new_n280), .A4(new_n287), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n487), .A2(new_n488), .A3(new_n383), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n488), .B1(new_n487), .B2(new_n383), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT4), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n517), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n516), .B1(new_n523), .B2(new_n474), .ZN(new_n524));
  INV_X1    g323(.A(new_n517), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n492), .B2(new_n490), .ZN(new_n526));
  INV_X1    g325(.A(new_n474), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(KEYINPUT80), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT39), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n500), .B2(new_n474), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n531), .A2(new_n507), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT81), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n523), .A2(new_n516), .A3(new_n474), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT80), .B1(new_n526), .B2(new_n527), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n529), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT40), .A4(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n536), .A2(KEYINPUT40), .A3(new_n507), .A4(new_n531), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT81), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT40), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n531), .A2(new_n507), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT39), .B1(new_n524), .B2(new_n528), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n469), .A2(new_n471), .B1(new_n508), .B2(new_n502), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n537), .A2(new_n539), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n334), .A2(new_n337), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n338), .A2(new_n321), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n404), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n460), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n397), .B1(new_n549), .B2(new_n465), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n462), .A2(new_n463), .A3(new_n406), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT37), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT38), .ZN(new_n553));
  INV_X1    g352(.A(new_n459), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n464), .A2(new_n467), .A3(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n552), .A2(new_n553), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT82), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n464), .A2(new_n467), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n459), .B1(new_n560), .B2(KEYINPUT37), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n561), .A2(KEYINPUT82), .A3(new_n553), .A4(new_n556), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n559), .A2(new_n470), .A3(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n512), .A2(KEYINPUT83), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n510), .A2(new_n509), .B1(new_n512), .B2(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(KEYINPUT84), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT84), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n555), .B1(new_n464), .B2(new_n467), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n568), .B2(new_n459), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n569), .A3(new_n556), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT38), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n563), .A2(new_n564), .A3(new_n565), .A4(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n431), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n430), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT79), .B1(new_n450), .B2(new_n430), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n545), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n361), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n360), .B1(new_n352), .B2(new_n350), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n453), .A2(new_n454), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(new_n573), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT35), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n514), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n515), .A2(new_n577), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n472), .B1(new_n565), .B2(new_n564), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n576), .A2(new_n580), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n584), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n261), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT21), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT89), .ZN(new_n592));
  INV_X1    g391(.A(G57gat), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT90), .ZN(new_n594));
  OAI21_X1  g393(.A(G64gat), .B1(KEYINPUT89), .B2(G57gat), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n593), .A2(G64gat), .ZN(new_n596));
  OAI22_X1  g395(.A1(new_n594), .A2(new_n595), .B1(new_n596), .B2(KEYINPUT90), .ZN(new_n597));
  NAND2_X1  g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  OR2_X1    g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT9), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n598), .B(new_n599), .C1(new_n603), .C2(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n236), .B1(new_n591), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G183gat), .ZN(new_n607));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT92), .ZN(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT91), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n609), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n607), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n605), .A2(new_n591), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G211gat), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G85gat), .A2(G92gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT7), .ZN(new_n624));
  NAND2_X1  g423(.A1(G99gat), .A2(G106gat), .ZN(new_n625));
  AOI22_X1  g424(.A1(KEYINPUT8), .A2(new_n625), .B1(new_n506), .B2(new_n458), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G99gat), .B(G106gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n605), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n624), .A2(new_n626), .ZN(new_n633));
  INV_X1    g432(.A(new_n628), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n635), .A2(new_n602), .A3(new_n604), .A4(new_n629), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n632), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n630), .A2(new_n631), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n639), .A2(KEYINPUT10), .A3(new_n602), .A4(new_n604), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n622), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G176gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(G204gat), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n621), .B1(new_n632), .B2(new_n636), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT95), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n645), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n641), .B2(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G190gat), .B(G218gat), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT93), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT94), .ZN(new_n658));
  INV_X1    g457(.A(new_n639), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n230), .A2(new_n237), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n227), .A2(new_n229), .A3(new_n639), .ZN(new_n661));
  AND2_X1   g460(.A1(G232gat), .A2(G233gat), .ZN(new_n662));
  AOI22_X1  g461(.A1(new_n655), .A2(new_n656), .B1(KEYINPUT41), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n658), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n662), .A2(KEYINPUT41), .ZN(new_n666));
  XNOR2_X1  g465(.A(G134gat), .B(G162gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n230), .A2(new_n237), .A3(new_n659), .ZN(new_n669));
  INV_X1    g468(.A(new_n658), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n669), .A2(new_n670), .A3(new_n661), .A4(new_n663), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n665), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n668), .B1(new_n665), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n620), .A2(new_n654), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n590), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n513), .A2(KEYINPUT96), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n513), .A2(KEYINPUT96), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(new_n232), .ZN(G1324gat));
  INV_X1    g481(.A(new_n677), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n472), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(G8gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(G1325gat));
  NOR3_X1   g489(.A1(new_n677), .A2(G15gat), .A3(new_n581), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n364), .B(KEYINPUT97), .Z(new_n692));
  NAND2_X1  g491(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n691), .B1(G15gat), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT98), .Z(G1326gat));
  NOR2_X1   g494(.A1(new_n677), .A2(new_n576), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT43), .B(G22gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(new_n680), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n620), .A2(new_n674), .A3(new_n653), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n590), .A2(new_n202), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT45), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT99), .B(KEYINPUT44), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  AOI211_X1 g504(.A(new_n674), .B(new_n705), .C1(new_n586), .C2(new_n589), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n515), .A2(new_n577), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n583), .A2(new_n585), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n589), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n674), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n620), .A2(new_n261), .A3(new_n653), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n703), .B1(new_n715), .B2(new_n680), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G29gat), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n715), .A2(new_n703), .A3(new_n680), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n702), .B1(new_n717), .B2(new_n718), .ZN(G1328gat));
  NAND4_X1  g518(.A1(new_n590), .A2(new_n203), .A3(new_n472), .A4(new_n700), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(KEYINPUT46), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT102), .Z(new_n722));
  OAI21_X1  g521(.A(G36gat), .B1(new_n715), .B2(new_n473), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(KEYINPUT46), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT101), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(G1329gat));
  INV_X1    g525(.A(new_n715), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n213), .B1(new_n727), .B2(new_n692), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n590), .A2(new_n700), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n581), .A2(G43gat), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n213), .B1(new_n727), .B2(new_n364), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT47), .ZN(new_n734));
  OAI22_X1  g533(.A1(new_n731), .A2(KEYINPUT47), .B1(new_n732), .B2(new_n734), .ZN(G1330gat));
  OAI21_X1  g534(.A(G50gat), .B1(new_n715), .B2(new_n576), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n729), .A2(new_n211), .A3(new_n455), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT48), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n738), .B(new_n740), .ZN(G1331gat));
  NAND4_X1  g540(.A1(new_n620), .A2(new_n261), .A3(new_n674), .A4(new_n653), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n586), .B2(new_n589), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n699), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT89), .B(G57gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1332gat));
  AOI21_X1  g545(.A(new_n473), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT104), .Z(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1333gat));
  NAND2_X1  g550(.A1(new_n743), .A2(new_n692), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n581), .A2(G71gat), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n752), .A2(G71gat), .B1(new_n743), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n743), .A2(new_n455), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  INV_X1    g556(.A(new_n260), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n257), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n759), .A2(new_n620), .A3(new_n654), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n706), .B2(new_n712), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g562(.A(KEYINPUT105), .B(new_n760), .C1(new_n706), .C2(new_n712), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(new_n699), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n506), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n766), .B2(new_n765), .ZN(new_n768));
  INV_X1    g567(.A(new_n620), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n710), .A2(new_n261), .A3(new_n769), .A4(new_n711), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT51), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n680), .A2(G85gat), .A3(new_n654), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT107), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n768), .B1(new_n771), .B2(new_n773), .ZN(G1336gat));
  NAND3_X1  g573(.A1(new_n653), .A2(new_n472), .A3(new_n458), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G92gat), .B1(new_n761), .B2(new_n473), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n472), .A3(new_n764), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(KEYINPUT51), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n770), .B(new_n783), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n775), .B(KEYINPUT108), .Z(new_n785));
  AOI21_X1  g584(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n778), .B1(new_n780), .B2(new_n786), .ZN(G1337gat));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n654), .ZN(new_n788));
  INV_X1    g587(.A(G99gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n789), .A3(new_n580), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n763), .A2(new_n692), .A3(new_n764), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(G1338gat));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n455), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT53), .B1(new_n788), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n713), .A2(new_n455), .A3(new_n760), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n763), .A2(new_n455), .A3(new_n764), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n800), .A2(new_n801), .A3(G106gat), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n800), .B2(G106gat), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n784), .A2(new_n653), .A3(new_n795), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n799), .B1(new_n805), .B2(new_n806), .ZN(G1339gat));
  NOR2_X1   g606(.A1(new_n680), .A2(new_n472), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n638), .A2(new_n640), .A3(new_n622), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT111), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n638), .A2(new_n640), .A3(new_n812), .A4(new_n622), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n811), .A2(new_n642), .A3(KEYINPUT54), .A4(new_n813), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n815));
  AOI21_X1  g614(.A(new_n645), .B1(new_n641), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n816), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n650), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n649), .B1(new_n817), .B2(new_n818), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n824), .A3(new_n820), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n261), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n253), .A2(new_n254), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n239), .B1(new_n238), .B2(new_n241), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n249), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n653), .A2(new_n257), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n674), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n257), .A2(new_n829), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n674), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n825), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n824), .B1(new_n823), .B2(new_n820), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n769), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n676), .A2(new_n261), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n809), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n583), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n261), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n285), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n271), .B2(new_n842), .ZN(G1340gat));
  NOR2_X1   g643(.A1(new_n841), .A2(new_n654), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(new_n269), .ZN(G1341gat));
  NOR2_X1   g645(.A1(new_n841), .A2(new_n769), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(new_n265), .ZN(G1342gat));
  NAND4_X1  g647(.A1(new_n840), .A2(new_n263), .A3(new_n583), .A4(new_n711), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n841), .B2(new_n674), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(G1343gat));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n620), .B1(new_n831), .B2(new_n836), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n675), .A2(new_n759), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n857), .B(new_n455), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n821), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n830), .B1(new_n759), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n836), .B1(new_n862), .B2(new_n711), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n859), .B1(new_n863), .B2(new_n769), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT57), .B1(new_n864), .B2(new_n576), .ZN(new_n865));
  INV_X1    g664(.A(new_n364), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n699), .A2(new_n473), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n860), .A2(new_n865), .A3(new_n759), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G141gat), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n692), .A2(new_n576), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n872), .B(new_n808), .C1(new_n858), .C2(new_n859), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n261), .A2(G141gat), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n876));
  AND2_X1   g675(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n877));
  OAI221_X1 g676(.A(new_n871), .B1(new_n873), .B2(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n873), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(KEYINPUT117), .A3(new_n874), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n873), .B2(new_n875), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n871), .A2(KEYINPUT116), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n885), .A3(G141gat), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n878), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n878), .B(KEYINPUT119), .C1(new_n887), .C2(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1344gat));
  NAND3_X1  g692(.A1(new_n879), .A2(new_n366), .A3(new_n653), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n869), .A2(new_n653), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n839), .B(KEYINPUT120), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n862), .A2(new_n711), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n833), .A2(new_n861), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n620), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n857), .B(new_n455), .C1(new_n897), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n576), .B1(new_n838), .B2(new_n839), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n896), .B(new_n901), .C1(new_n857), .C2(new_n902), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n903), .A2(KEYINPUT121), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n366), .B1(new_n903), .B2(KEYINPUT121), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n895), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n860), .A2(new_n865), .A3(new_n869), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n654), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(KEYINPUT59), .A3(new_n366), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n894), .B1(new_n906), .B2(new_n909), .ZN(G1345gat));
  OAI21_X1  g709(.A(G155gat), .B1(new_n907), .B2(new_n769), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n879), .A2(new_n373), .A3(new_n620), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1346gat));
  OR2_X1    g712(.A1(new_n907), .A2(new_n674), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n374), .B1(new_n914), .B2(KEYINPUT122), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(KEYINPUT122), .B2(new_n914), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n879), .A2(new_n374), .A3(new_n711), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1347gat));
  AOI21_X1  g717(.A(new_n699), .B1(new_n838), .B2(new_n839), .ZN(new_n919));
  INV_X1    g718(.A(new_n583), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n473), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n301), .B1(new_n923), .B2(new_n261), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n680), .A2(new_n472), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT123), .ZN(new_n926));
  AOI211_X1 g725(.A(new_n920), .B(new_n926), .C1(new_n838), .C2(new_n839), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(G169gat), .A3(new_n759), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT124), .Z(G1348gat));
  AOI21_X1  g729(.A(G176gat), .B1(new_n922), .B2(new_n653), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n654), .A2(new_n326), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n927), .B2(new_n932), .ZN(G1349gat));
  AOI21_X1  g732(.A(new_n289), .B1(new_n927), .B2(new_n620), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n620), .A2(new_n309), .A3(new_n311), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n922), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n290), .A3(new_n711), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT125), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n290), .B1(new_n927), .B2(new_n711), .ZN(new_n940));
  XNOR2_X1  g739(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n942), .ZN(G1351gat));
  NAND3_X1  g742(.A1(new_n919), .A2(new_n472), .A3(new_n872), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(new_n261), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n926), .A2(new_n692), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n901), .B(new_n946), .C1(new_n902), .C2(new_n857), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n759), .A2(G197gat), .ZN(new_n948));
  OAI22_X1  g747(.A1(G197gat), .A2(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(G1352gat));
  NOR3_X1   g749(.A1(new_n944), .A2(G204gat), .A3(new_n654), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  OAI21_X1  g751(.A(G204gat), .B1(new_n947), .B2(new_n654), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1353gat));
  OAI21_X1  g753(.A(G211gat), .B1(new_n947), .B2(new_n769), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT63), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n944), .A2(G211gat), .A3(new_n769), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n956), .A2(new_n957), .ZN(G1354gat));
  NOR2_X1   g757(.A1(new_n944), .A2(new_n674), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n711), .A2(G218gat), .ZN(new_n960));
  OAI22_X1  g759(.A1(G218gat), .A2(new_n959), .B1(new_n947), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT127), .Z(G1355gat));
endmodule


