//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943;
  XNOR2_X1  g000(.A(G128), .B(G143), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT13), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  OAI211_X1 g004(.A(new_n188), .B(G134), .C1(KEYINPUT13), .C2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G116), .B(G122), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n187), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n187), .B(new_n195), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(new_n193), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT14), .A3(G122), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(G107), .A3(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(new_n199), .A3(new_n204), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT9), .B(G234), .Z(new_n206));
  INV_X1    g020(.A(G953), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(G217), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n197), .A2(new_n205), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(new_n197), .B2(new_n205), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G902), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G478), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n214), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(G210), .B1(G237), .B2(G902), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT66), .B1(new_n189), .B2(G146), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n189), .A2(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT65), .A2(KEYINPUT0), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(KEYINPUT65), .B2(KEYINPUT0), .ZN(new_n230));
  NOR3_X1   g044(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n226), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n223), .A2(G143), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n234), .A2(new_n225), .A3(KEYINPUT0), .A4(G128), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G125), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT85), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G224), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(G953), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n189), .A2(G146), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n244));
  OAI21_X1  g058(.A(G128), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n226), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G125), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n234), .A2(new_n225), .A3(new_n244), .A4(G128), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT86), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n239), .A2(new_n242), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n242), .B1(new_n239), .B2(new_n250), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT2), .A2(G113), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NOR3_X1   g070(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G116), .B(G119), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G104), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT3), .B1(new_n262), .B2(G107), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n193), .A3(G104), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(G107), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G101), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT80), .B(G101), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n269), .A2(new_n266), .A3(new_n265), .A4(new_n263), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(KEYINPUT4), .A3(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n261), .B(new_n271), .C1(KEYINPUT4), .C2(new_n268), .ZN(new_n272));
  INV_X1    g086(.A(new_n266), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n262), .A2(G107), .ZN(new_n274));
  OAI21_X1  g088(.A(G101), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n258), .A2(new_n260), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n279));
  OR3_X1    g093(.A1(new_n202), .A2(KEYINPUT5), .A3(G119), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(G113), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT82), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n279), .A2(KEYINPUT82), .A3(new_n280), .A4(G113), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n278), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  XOR2_X1   g099(.A(G110), .B(G122), .Z(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n272), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT83), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT6), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT84), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n272), .A2(new_n285), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT84), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n287), .B1(new_n293), .B2(KEYINPUT6), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n295), .A3(KEYINPUT84), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n253), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n286), .B(KEYINPUT8), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n283), .B(new_n284), .C1(new_n258), .C2(new_n260), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n302), .A2(new_n276), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n278), .A2(new_n281), .ZN(new_n304));
  OAI211_X1 g118(.A(KEYINPUT87), .B(new_n301), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT87), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n302), .A2(new_n276), .B1(new_n278), .B2(new_n281), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(new_n300), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n250), .A2(new_n237), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT7), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(new_n241), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n305), .A2(new_n308), .A3(new_n311), .A4(new_n288), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n239), .A2(KEYINPUT7), .A3(new_n242), .A4(new_n250), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n213), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n220), .B1(new_n299), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n252), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n239), .A2(new_n242), .A3(new_n250), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n290), .A2(KEYINPUT84), .A3(new_n295), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n295), .B1(new_n290), .B2(KEYINPUT84), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n311), .A2(new_n288), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(new_n313), .A3(new_n308), .A4(new_n305), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n322), .A2(new_n324), .A3(new_n213), .A4(new_n219), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G952), .ZN(new_n327));
  AOI211_X1 g141(.A(G953), .B(new_n327), .C1(G234), .C2(G237), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI211_X1 g143(.A(new_n213), .B(new_n207), .C1(G234), .C2(G237), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT21), .B(G898), .Z(new_n332));
  OAI21_X1  g146(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G214), .B1(G237), .B2(G902), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n326), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT20), .ZN(new_n336));
  XNOR2_X1  g150(.A(G113), .B(G122), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(new_n262), .ZN(new_n338));
  AND2_X1   g152(.A1(KEYINPUT71), .A2(G237), .ZN(new_n339));
  NOR2_X1   g153(.A1(KEYINPUT71), .A2(G237), .ZN(new_n340));
  OAI211_X1 g154(.A(G214), .B(new_n207), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n189), .A2(KEYINPUT88), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT88), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G143), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G131), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n341), .A2(new_n346), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n346), .B1(new_n341), .B2(new_n343), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT71), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(KEYINPUT71), .A2(G237), .ZN(new_n356));
  AOI21_X1  g170(.A(G953), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n347), .B1(new_n357), .B2(G214), .ZN(new_n358));
  OAI21_X1  g172(.A(G131), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT17), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n351), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(KEYINPUT17), .B(G131), .C1(new_n352), .C2(new_n358), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n247), .A2(KEYINPUT16), .A3(G140), .ZN(new_n363));
  XNOR2_X1  g177(.A(G125), .B(G140), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(KEYINPUT16), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n365), .A2(G146), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(G146), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n361), .A2(new_n362), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n352), .A2(new_n358), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT18), .A2(G131), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT89), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT90), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n374), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT90), .ZN(new_n377));
  NOR4_X1   g191(.A1(new_n352), .A2(new_n358), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(KEYINPUT18), .B(G131), .C1(new_n352), .C2(new_n358), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n364), .B(new_n223), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT91), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n342), .B1(new_n357), .B2(G214), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n350), .B(new_n374), .C1(new_n384), .C2(new_n346), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n377), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n348), .A2(KEYINPUT90), .A3(new_n350), .A4(new_n374), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT91), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n380), .A2(new_n381), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n338), .B(new_n371), .C1(new_n383), .C2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT92), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n389), .B1(new_n388), .B2(new_n390), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n382), .A2(KEYINPUT91), .A3(new_n386), .A4(new_n387), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n370), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(KEYINPUT92), .A3(new_n338), .ZN(new_n398));
  INV_X1    g212(.A(new_n338), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n351), .A2(new_n359), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n364), .B(KEYINPUT19), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n223), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n367), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n383), .B2(new_n391), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n394), .A2(new_n398), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(G475), .A2(G902), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n336), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT93), .B(G475), .Z(new_n409));
  NOR2_X1   g223(.A1(new_n397), .A2(new_n338), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n394), .B2(new_n398), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n411), .B2(G902), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n404), .A2(new_n399), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n397), .A2(KEYINPUT92), .A3(new_n338), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT92), .B1(new_n397), .B2(new_n338), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT20), .A3(new_n406), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n408), .A2(new_n412), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT94), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n408), .A2(new_n412), .A3(new_n417), .A4(KEYINPUT94), .ZN(new_n421));
  AOI211_X1 g235(.A(new_n218), .B(new_n335), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT31), .ZN(new_n423));
  INV_X1    g237(.A(G137), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(G134), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(KEYINPUT67), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n195), .A2(KEYINPUT67), .A3(G137), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(G134), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G131), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT11), .B1(new_n195), .B2(G137), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT11), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n424), .A3(G134), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n425), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n349), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT70), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n246), .A2(new_n438), .A3(new_n248), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n246), .B2(new_n248), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI211_X1 g255(.A(G131), .B(new_n425), .C1(new_n431), .C2(new_n433), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n349), .B1(new_n434), .B2(new_n435), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT69), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n444), .A2(new_n236), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n432), .B1(G134), .B2(new_n424), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n195), .A2(KEYINPUT11), .A3(G137), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n435), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G131), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n436), .ZN(new_n451));
  INV_X1    g265(.A(new_n235), .ZN(new_n452));
  NOR2_X1   g266(.A1(KEYINPUT65), .A2(KEYINPUT0), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n228), .B2(new_n227), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(new_n231), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n452), .B1(new_n455), .B2(new_n226), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT69), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(KEYINPUT30), .B(new_n441), .C1(new_n446), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n246), .A2(new_n248), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n437), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n451), .A2(new_n456), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n458), .A2(new_n261), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n261), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n466), .B(new_n441), .C1(new_n446), .C2(new_n457), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n357), .A2(G210), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n468), .B(new_n469), .Z(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT26), .B(G101), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n470), .B(new_n471), .Z(new_n472));
  NAND3_X1  g286(.A1(new_n465), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT73), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n465), .A2(new_n472), .A3(KEYINPUT73), .A4(new_n467), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n423), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n462), .A2(new_n261), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n467), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT28), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n441), .A2(new_n466), .A3(new_n461), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT28), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n472), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n473), .A2(KEYINPUT31), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n477), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(G472), .A2(G902), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n487), .B(KEYINPUT74), .Z(new_n488));
  OAI21_X1  g302(.A(KEYINPUT32), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n475), .A2(new_n476), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT31), .ZN(new_n491));
  INV_X1    g305(.A(new_n484), .ZN(new_n492));
  INV_X1    g306(.A(new_n485), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT32), .ZN(new_n495));
  INV_X1    g309(.A(new_n488), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n480), .A2(new_n483), .A3(new_n472), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n465), .A2(new_n467), .ZN(new_n499));
  INV_X1    g313(.A(new_n472), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT29), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n441), .B1(new_n446), .B2(new_n457), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n261), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n467), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n506), .A2(KEYINPUT75), .A3(KEYINPUT28), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT75), .B1(new_n506), .B2(KEYINPUT28), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT29), .B(new_n483), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  OAI221_X1 g323(.A(new_n213), .B1(new_n498), .B2(new_n503), .C1(new_n509), .C2(new_n500), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n489), .A2(new_n497), .B1(new_n510), .B2(G472), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n228), .A2(G119), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT23), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n228), .A2(G119), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT76), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(new_n518), .A3(new_n515), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(G110), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n515), .A2(new_n512), .ZN(new_n521));
  XOR2_X1   g335(.A(KEYINPUT24), .B(G110), .Z(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n368), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n364), .A2(new_n223), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n516), .A2(G110), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n521), .A2(new_n522), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n367), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT77), .B(KEYINPUT22), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(G137), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n207), .A2(G221), .A3(G234), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n524), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n524), .B2(new_n528), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n213), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT25), .ZN(new_n536));
  INV_X1    g350(.A(G217), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(G234), .B2(new_n213), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n539), .B(new_n213), .C1(new_n533), .C2(new_n534), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT78), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n538), .A2(G902), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n533), .B2(new_n534), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n542), .B1(new_n541), .B2(new_n544), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n511), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G469), .ZN(new_n549));
  INV_X1    g363(.A(new_n276), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT10), .B(new_n550), .C1(new_n439), .C2(new_n440), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n234), .A2(new_n225), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n245), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n248), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT10), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n456), .B(new_n271), .C1(KEYINPUT4), .C2(new_n268), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n551), .A2(new_n557), .A3(new_n444), .A4(new_n558), .ZN(new_n559));
  XOR2_X1   g373(.A(G110), .B(G140), .Z(new_n560));
  INV_X1    g374(.A(G227), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(G953), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n560), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  OR3_X1    g378(.A1(new_n550), .A2(new_n459), .A3(KEYINPUT81), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT81), .B1(new_n550), .B2(new_n459), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n555), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n451), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(KEYINPUT12), .A3(new_n451), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n564), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n551), .A2(new_n557), .A3(new_n558), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n451), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n563), .B1(new_n574), .B2(new_n559), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n549), .B(new_n213), .C1(new_n572), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(G469), .A2(G902), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n559), .A3(new_n563), .ZN(new_n578));
  INV_X1    g392(.A(new_n559), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n570), .B2(new_n571), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n563), .B(KEYINPUT79), .Z(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n578), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n576), .B(new_n577), .C1(new_n583), .C2(new_n549), .ZN(new_n584));
  INV_X1    g398(.A(new_n206), .ZN(new_n585));
  OAI21_X1  g399(.A(G221), .B1(new_n585), .B2(G902), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n422), .A2(new_n548), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n589), .B(new_n269), .Z(G3));
  OAI21_X1  g404(.A(KEYINPUT33), .B1(new_n211), .B2(KEYINPUT96), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n212), .B(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n592), .A2(new_n215), .A3(G902), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n593), .A2(KEYINPUT97), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(KEYINPUT97), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n214), .A2(new_n215), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n420), .A2(new_n421), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  INV_X1    g413(.A(new_n335), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n600), .A2(new_n420), .A3(new_n421), .A4(new_n597), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT98), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT95), .B1(new_n486), .B2(G902), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n494), .A2(new_n605), .A3(new_n213), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n606), .A3(G472), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n547), .A2(new_n587), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n494), .A2(new_n496), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n601), .A2(new_n603), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  OR2_X1    g427(.A1(new_n418), .A2(new_n217), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n335), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NAND2_X1  g432(.A1(new_n524), .A2(new_n528), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n543), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n541), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT99), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n607), .A2(new_n609), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n607), .A2(KEYINPUT100), .A3(new_n609), .A4(new_n624), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n627), .A2(new_n588), .A3(new_n422), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G110), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  INV_X1    g446(.A(new_n334), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n623), .B(KEYINPUT99), .Z(new_n634));
  INV_X1    g448(.A(new_n326), .ZN(new_n635));
  NOR4_X1   g449(.A1(new_n511), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT102), .B(G900), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n331), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n638), .A2(KEYINPUT103), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(KEYINPUT103), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n329), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n614), .A2(new_n587), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  XOR2_X1   g459(.A(new_n641), .B(KEYINPUT39), .Z(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n584), .A2(new_n586), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n634), .B1(new_n648), .B2(KEYINPUT40), .ZN(new_n649));
  INV_X1    g463(.A(new_n506), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n490), .B1(new_n472), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n213), .ZN(new_n652));
  AOI22_X1  g466(.A1(new_n489), .A2(new_n497), .B1(G472), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT38), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n326), .B(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n649), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n420), .A2(new_n421), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n217), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n656), .A2(new_n334), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G143), .ZN(G45));
  NAND4_X1  g475(.A1(new_n420), .A2(new_n421), .A3(new_n597), .A4(new_n641), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n587), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n636), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G146), .ZN(G48));
  OR2_X1    g479(.A1(new_n572), .A2(new_n575), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n213), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(new_n586), .A3(new_n576), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n601), .A2(new_n548), .A3(new_n603), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT41), .B(G113), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  NAND3_X1  g487(.A1(new_n548), .A2(new_n615), .A3(new_n670), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G116), .ZN(G18));
  NAND2_X1  g489(.A1(new_n489), .A2(new_n497), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n510), .A2(G472), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n634), .A2(new_n669), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n422), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  OAI21_X1  g495(.A(G472), .B1(new_n486), .B2(G902), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n483), .B1(new_n507), .B2(new_n508), .ZN(new_n683));
  AOI211_X1 g497(.A(new_n485), .B(new_n477), .C1(new_n500), .C2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n682), .B1(new_n684), .B2(new_n488), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n541), .A2(new_n544), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n658), .A2(new_n600), .A3(new_n670), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G122), .ZN(G24));
  NOR2_X1   g503(.A1(new_n662), .A2(new_n685), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n635), .A2(new_n633), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n691), .A3(new_n679), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT104), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n247), .ZN(G27));
  NOR2_X1   g508(.A1(new_n326), .A2(new_n633), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n511), .A2(new_n547), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n663), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n663), .A2(KEYINPUT105), .A3(new_n697), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n704));
  INV_X1    g518(.A(new_n686), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n704), .B1(new_n678), .B2(new_n705), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n511), .A2(KEYINPUT106), .A3(new_n686), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n662), .A2(new_n696), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(KEYINPUT42), .A3(new_n588), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G131), .ZN(G33));
  NAND2_X1  g526(.A1(new_n697), .A2(new_n643), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G134), .ZN(G36));
  NAND2_X1  g528(.A1(new_n657), .A2(new_n597), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT43), .B1(new_n657), .B2(new_n597), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n607), .A2(new_n609), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(KEYINPUT44), .A3(new_n720), .A4(new_n624), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n720), .B(new_n624), .C1(new_n717), .C2(new_n718), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n578), .B(KEYINPUT45), .C1(new_n580), .C2(new_n582), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n725), .A2(KEYINPUT107), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n549), .B1(new_n583), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n725), .A2(KEYINPUT107), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n577), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT108), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n730), .A2(new_n735), .A3(KEYINPUT46), .A4(new_n577), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n733), .A2(new_n734), .A3(new_n576), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n586), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n646), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n721), .A2(new_n724), .A3(new_n695), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G137), .ZN(G39));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n737), .A2(KEYINPUT47), .A3(new_n586), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n678), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n547), .A3(new_n709), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G140), .ZN(G42));
  NAND2_X1  g561(.A1(new_n327), .A2(new_n207), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n636), .B1(new_n663), .B2(new_n643), .ZN(new_n750));
  INV_X1    g564(.A(new_n653), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n641), .B(KEYINPUT111), .Z(new_n752));
  NAND3_X1  g566(.A1(new_n541), .A2(new_n622), .A3(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n753), .A2(KEYINPUT112), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(KEYINPUT112), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n587), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n658), .A2(new_n691), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n750), .A2(new_n692), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT53), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n671), .A2(new_n674), .A3(new_n680), .A4(new_n688), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n217), .B1(new_n420), .B2(new_n421), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n610), .B(new_n600), .C1(new_n598), .C2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n629), .A2(new_n589), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n629), .A2(new_n764), .A3(new_n589), .A4(KEYINPUT109), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n408), .A2(new_n412), .A3(new_n417), .A4(new_n641), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n511), .A2(new_n218), .A3(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n624), .B(new_n695), .C1(new_n690), .C2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n713), .B1(new_n772), .B2(new_n587), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n703), .B2(new_n710), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n761), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n769), .A2(new_n774), .A3(KEYINPUT110), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT110), .B1(new_n769), .B2(new_n774), .ZN(new_n779));
  INV_X1    g593(.A(new_n760), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n749), .B(new_n777), .C1(new_n781), .C2(KEYINPUT53), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT113), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n775), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n769), .A2(new_n774), .A3(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI22_X1  g601(.A1(new_n781), .A2(KEYINPUT53), .B1(new_n787), .B2(new_n761), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT54), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n785), .A2(new_n760), .A3(new_n786), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n776), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n793), .A3(new_n749), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n783), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n696), .A2(new_n669), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n328), .B(new_n796), .C1(new_n717), .C2(new_n718), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n706), .A2(new_n707), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n797), .A2(KEYINPUT48), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT116), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT48), .B1(new_n797), .B2(new_n798), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n799), .A2(KEYINPUT116), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n800), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n327), .A2(G953), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n719), .A2(new_n328), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n808), .A2(new_n670), .A3(new_n687), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n691), .ZN(new_n810));
  INV_X1    g624(.A(new_n547), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n796), .A2(new_n653), .A3(new_n811), .A4(new_n328), .ZN(new_n812));
  INV_X1    g626(.A(new_n598), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n806), .A2(new_n807), .A3(new_n810), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT118), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n668), .A2(new_n576), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n743), .B(new_n744), .C1(new_n586), .C2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n808), .A3(new_n687), .A4(new_n695), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT51), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n655), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n334), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n809), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n809), .A2(KEYINPUT50), .A3(new_n824), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n597), .B(new_n812), .C1(new_n420), .C2(new_n421), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT114), .Z(new_n831));
  OR3_X1    g645(.A1(new_n797), .A2(new_n634), .A3(new_n685), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n831), .A2(new_n820), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n822), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n829), .A2(new_n822), .A3(new_n833), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n817), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n748), .B1(new_n795), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n818), .B(KEYINPUT49), .Z(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n705), .A3(new_n586), .A4(new_n334), .ZN(new_n839));
  OR4_X1    g653(.A1(new_n823), .A2(new_n839), .A3(new_n751), .A4(new_n715), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n840), .ZN(G75));
  OAI21_X1  g655(.A(new_n777), .B1(new_n781), .B2(KEYINPUT53), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(G210), .A3(G902), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT56), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n320), .A2(new_n321), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(new_n319), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT55), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(KEYINPUT119), .B2(new_n844), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n845), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n207), .A2(G952), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n843), .A2(new_n844), .A3(new_n850), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(G51));
  OR2_X1    g670(.A1(new_n577), .A2(KEYINPUT57), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n577), .A2(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n790), .A2(new_n791), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n749), .B1(new_n859), .B2(new_n777), .ZN(new_n860));
  AOI211_X1 g674(.A(KEYINPUT54), .B(new_n776), .C1(new_n790), .C2(new_n791), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n857), .B(new_n858), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n666), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n792), .A2(new_n213), .A3(new_n730), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n853), .B1(new_n863), .B2(new_n864), .ZN(G54));
  NOR2_X1   g679(.A1(new_n792), .A2(new_n213), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(KEYINPUT58), .A3(G475), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n405), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n866), .A2(KEYINPUT58), .A3(G475), .A4(new_n416), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n868), .A2(new_n854), .A3(new_n869), .ZN(G60));
  NAND2_X1  g684(.A1(G478), .A2(G902), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT59), .Z(new_n872));
  NOR2_X1   g686(.A1(new_n592), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n860), .B2(new_n861), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n854), .ZN(new_n875));
  INV_X1    g689(.A(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n795), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n875), .B1(new_n877), .B2(new_n592), .ZN(G63));
  NAND2_X1  g692(.A1(G217), .A2(G902), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT120), .Z(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT60), .Z(new_n881));
  NAND2_X1  g695(.A1(new_n842), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n533), .A2(new_n534), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n853), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n842), .A2(new_n621), .A3(new_n881), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(KEYINPUT61), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT61), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  INV_X1    g702(.A(new_n881), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n883), .B1(new_n792), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n885), .A2(new_n890), .A3(new_n854), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n892), .ZN(G66));
  AND2_X1   g707(.A1(new_n332), .A2(G224), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT122), .B1(new_n894), .B2(new_n207), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n769), .A2(G953), .ZN(new_n896));
  MUX2_X1   g710(.A(new_n895), .B(KEYINPUT122), .S(new_n896), .Z(new_n897));
  OAI21_X1  g711(.A(new_n846), .B1(G898), .B2(new_n207), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(G69));
  AND4_X1   g713(.A1(new_n692), .A2(new_n711), .A3(new_n713), .A4(new_n750), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n739), .A2(new_n691), .A3(new_n658), .A4(new_n708), .ZN(new_n901));
  AND4_X1   g715(.A1(new_n740), .A2(new_n900), .A3(new_n746), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n207), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n458), .A2(new_n464), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(new_n401), .Z(new_n905));
  NAND2_X1  g719(.A1(G900), .A2(G953), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(G900), .ZN(new_n908));
  OAI21_X1  g722(.A(G953), .B1(new_n561), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n910));
  INV_X1    g724(.A(new_n648), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n598), .A2(new_n763), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n598), .B2(new_n763), .ZN(new_n914));
  AND4_X1   g728(.A1(new_n911), .A2(new_n913), .A3(new_n697), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n660), .A2(new_n750), .A3(new_n692), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n660), .A2(new_n750), .A3(KEYINPUT62), .A4(new_n692), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n740), .A3(new_n746), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n920), .A2(new_n740), .A3(KEYINPUT125), .A4(new_n746), .ZN(new_n924));
  AOI21_X1  g738(.A(G953), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n905), .B(KEYINPUT123), .Z(new_n926));
  OAI211_X1 g740(.A(new_n907), .B(new_n910), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G72));
  INV_X1    g743(.A(new_n499), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n902), .A2(new_n769), .ZN(new_n931));
  NAND2_X1  g745(.A1(G472), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT63), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n500), .B(new_n930), .C1(new_n931), .C2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n923), .A2(new_n769), .A3(new_n924), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n930), .B1(new_n936), .B2(new_n933), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n472), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n937), .B2(new_n472), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n854), .B(new_n935), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n490), .A2(new_n501), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n788), .A2(new_n933), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n941), .A2(new_n943), .ZN(G57));
endmodule


