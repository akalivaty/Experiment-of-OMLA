//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G57gat), .ZN(new_n204));
  INV_X1    g003(.A(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT5), .ZN(new_n208));
  NAND2_X1  g007(.A1(G225gat), .A2(G233gat), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n209), .B(KEYINPUT76), .Z(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT68), .ZN(new_n212));
  INV_X1    g011(.A(G113gat), .ZN(new_n213));
  INV_X1    g012(.A(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g015(.A1(G113gat), .A2(G120gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G127gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G134gat), .ZN(new_n220));
  INV_X1    g019(.A(G134gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G127gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n212), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT1), .B1(new_n213), .B2(new_n214), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n225), .A2(KEYINPUT68), .A3(new_n217), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n221), .A2(G127gat), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n226), .A2(new_n217), .B1(new_n229), .B2(KEYINPUT67), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT74), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(G155gat), .B2(G162gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(G141gat), .B(G148gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(G155gat), .B2(G162gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G155gat), .B(G162gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G155gat), .A2(G162gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT2), .ZN(new_n245));
  INV_X1    g044(.A(G141gat), .ZN(new_n246));
  INV_X1    g045(.A(G148gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G141gat), .A2(G148gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n241), .A3(new_n236), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n243), .A2(KEYINPUT3), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n250), .A2(new_n241), .A3(new_n236), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n241), .B1(new_n250), .B2(new_n236), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT75), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n251), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT75), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n260), .A3(new_n254), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n253), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n224), .A2(new_n227), .B1(new_n232), .B2(new_n230), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n263), .A3(KEYINPUT4), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n211), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n255), .A2(new_n256), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n234), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n268), .B1(KEYINPUT4), .B2(new_n211), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT77), .B1(new_n259), .B2(new_n263), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT77), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n234), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n270), .A2(new_n272), .A3(new_n210), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n208), .B1(new_n266), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n263), .B1(new_n267), .B2(KEYINPUT3), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n260), .B1(new_n259), .B2(new_n254), .ZN(new_n277));
  AOI211_X1 g076(.A(KEYINPUT75), .B(KEYINPUT3), .C1(new_n243), .C2(new_n251), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n263), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT78), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n280), .A2(new_n282), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT78), .B1(new_n286), .B2(new_n264), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n210), .A2(KEYINPUT5), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n285), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n207), .B1(new_n275), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n264), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n281), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n258), .A2(new_n261), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n294), .A2(new_n276), .B1(new_n280), .B2(new_n283), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n295), .A3(new_n288), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n264), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n297), .A2(new_n211), .B1(new_n273), .B2(new_n269), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n206), .B(new_n296), .C1(new_n298), .C2(new_n208), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT6), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n291), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT6), .B(new_n207), .C1(new_n275), .C2(new_n290), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT22), .ZN(new_n307));
  NAND2_X1  g106(.A1(G211gat), .A2(G218gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n312), .A2(KEYINPUT73), .A3(new_n308), .ZN(new_n313));
  XNOR2_X1  g112(.A(G197gat), .B(G204gat), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n309), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n309), .B2(new_n314), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(KEYINPUT23), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(KEYINPUT23), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(KEYINPUT66), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT24), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT24), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(G183gat), .A3(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR3_X1   g128(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n332), .A2(G169gat), .A3(G176gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT66), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT25), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n322), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n324), .A2(new_n326), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(G169gat), .B2(G176gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n340), .A3(new_n318), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT25), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(KEYINPUT27), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT27), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G183gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n345), .A3(new_n338), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT28), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n343), .A2(new_n345), .A3(new_n348), .A4(new_n338), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT26), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n319), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n318), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n347), .A2(new_n323), .A3(new_n349), .A4(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n342), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(G226gat), .A3(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n355), .A2(new_n358), .B1(G226gat), .B2(G233gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n317), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n355), .A2(new_n358), .ZN(new_n361));
  NAND2_X1  g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n317), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n364), .A3(new_n356), .ZN(new_n365));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(G64gat), .ZN(new_n367));
  INV_X1    g166(.A(G92gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n360), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT30), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n360), .A2(new_n365), .A3(KEYINPUT30), .A4(new_n369), .ZN(new_n373));
  INV_X1    g172(.A(new_n369), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n357), .A2(new_n359), .A3(new_n317), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n364), .B1(new_n363), .B2(new_n356), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n372), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n303), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n309), .A2(new_n314), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n312), .A2(new_n308), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n358), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n381), .A2(new_n382), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n254), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n267), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n258), .B2(new_n261), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(new_n364), .ZN(new_n389));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n358), .B1(new_n277), .B2(new_n278), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n317), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n358), .B1(new_n315), .B2(new_n316), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n254), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n390), .B1(new_n396), .B2(new_n267), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n392), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n392), .B(new_n397), .C1(new_n388), .C2(new_n364), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n391), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G22gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n397), .B1(new_n388), .B2(new_n364), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT79), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n404), .A2(new_n399), .B1(new_n390), .B2(new_n389), .ZN(new_n405));
  INV_X1    g204(.A(G22gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT31), .ZN(new_n409));
  INV_X1    g208(.A(G50gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n402), .A2(new_n407), .A3(KEYINPUT80), .A4(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(new_n405), .B2(new_n406), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n415), .A2(new_n411), .B1(new_n402), .B2(new_n407), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n380), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n370), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT37), .B1(new_n375), .B2(new_n376), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT37), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n360), .A2(new_n365), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n374), .A3(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(KEYINPUT81), .B(KEYINPUT38), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n418), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n419), .A2(new_n374), .A3(new_n423), .A4(new_n421), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n301), .A2(new_n425), .A3(new_n302), .A4(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT80), .B1(new_n401), .B2(G22gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n411), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n405), .A2(new_n406), .ZN(new_n430));
  AOI221_X4 g229(.A(G22gat), .B1(new_n389), .B2(new_n390), .C1(new_n404), .C2(new_n399), .ZN(new_n431));
  OAI22_X1  g230(.A1(new_n428), .A2(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT40), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n211), .B1(new_n293), .B2(new_n295), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n270), .A2(new_n272), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(new_n211), .A3(new_n280), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT39), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n206), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n210), .B1(new_n285), .B2(new_n287), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(KEYINPUT39), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n433), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(KEYINPUT39), .A3(new_n436), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT39), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n442), .A2(new_n444), .A3(KEYINPUT40), .A4(new_n206), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n441), .A2(new_n291), .A3(new_n445), .A4(new_n378), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n427), .A2(new_n432), .A3(new_n446), .A4(new_n412), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT36), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT32), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n355), .A2(new_n263), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n234), .A2(new_n342), .A3(new_n354), .A4(new_n336), .ZN(new_n451));
  NAND2_X1  g250(.A1(G227gat), .A2(G233gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n452), .B(KEYINPUT64), .Z(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT69), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT69), .A4(new_n453), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n449), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n456), .B2(new_n457), .ZN(new_n461));
  XNOR2_X1  g260(.A(G15gat), .B(G43gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n458), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT71), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n467));
  INV_X1    g266(.A(new_n453), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n466), .B1(new_n469), .B2(KEYINPUT34), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT34), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n467), .A2(KEYINPUT71), .A3(new_n471), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(KEYINPUT34), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n464), .ZN(new_n475));
  AOI221_X4 g274(.A(new_n449), .B1(new_n475), .B2(new_n460), .C1(new_n456), .C2(new_n457), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n465), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n474), .ZN(new_n478));
  INV_X1    g277(.A(new_n458), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n456), .A2(new_n457), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n459), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n481), .A3(new_n475), .ZN(new_n482));
  INV_X1    g281(.A(new_n476), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n448), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n474), .B1(new_n465), .B2(new_n476), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(new_n483), .A3(new_n478), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(KEYINPUT36), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n417), .A2(new_n447), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n413), .A2(new_n416), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n378), .B1(new_n301), .B2(new_n302), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n477), .A2(new_n484), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n491), .A2(KEYINPUT35), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n493), .A2(new_n492), .A3(new_n432), .A4(new_n412), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n490), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n490), .A2(new_n494), .A3(new_n497), .A4(KEYINPUT82), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n410), .A2(G43gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n410), .A2(G43gat), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n504), .A2(KEYINPUT15), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507));
  INV_X1    g306(.A(G43gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT83), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT83), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G43gat), .ZN(new_n511));
  AOI21_X1  g310(.A(G50gat), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n507), .B1(new_n512), .B2(new_n503), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514));
  OR3_X1    g313(.A1(new_n514), .A2(G29gat), .A3(G36gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(G29gat), .B2(G36gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(G29gat), .A2(G36gat), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n506), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n504), .A2(KEYINPUT15), .A3(new_n505), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT17), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n506), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT83), .B(G43gat), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n504), .B1(new_n526), .B2(G50gat), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n520), .B1(new_n527), .B2(new_n507), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n524), .B(new_n525), .C1(new_n528), .C2(new_n506), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n406), .A2(G15gat), .ZN(new_n530));
  INV_X1    g329(.A(G15gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(G1gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT16), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(G1gat), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT84), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n536), .B2(G1gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(G8gat), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G8gat), .ZN(new_n541));
  OAI221_X1 g340(.A(new_n535), .B1(new_n538), .B2(new_n541), .C1(G1gat), .C2(new_n536), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n523), .A2(new_n529), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT85), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n519), .A2(new_n522), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n540), .A2(KEYINPUT85), .A3(new_n542), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT88), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT18), .A4(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n525), .B1(new_n528), .B2(new_n506), .ZN(new_n555));
  INV_X1    g354(.A(new_n549), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT85), .B1(new_n540), .B2(new_n542), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n559), .A3(new_n550), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT89), .A4(new_n549), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n553), .B(KEYINPUT13), .Z(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n550), .A3(new_n553), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT18), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT88), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n554), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n564), .A2(KEYINPUT86), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n565), .B1(new_n564), .B2(KEYINPUT86), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G113gat), .B(G141gat), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT11), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G169gat), .ZN(new_n573));
  INV_X1    g372(.A(G197gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT12), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n567), .B(new_n570), .C1(KEYINPUT87), .C2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n554), .A2(new_n566), .A3(KEYINPUT87), .A4(new_n563), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n575), .B(KEYINPUT12), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n554), .A2(new_n563), .A3(new_n566), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n568), .A2(new_n569), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT7), .B1(new_n205), .B2(new_n368), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(G85gat), .A3(G92gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G99gat), .B(G106gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  AOI22_X1  g390(.A1(KEYINPUT8), .A2(new_n591), .B1(new_n205), .B2(new_n368), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n590), .B1(new_n589), .B2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n523), .A2(new_n529), .A3(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n597), .A2(KEYINPUT93), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(KEYINPUT93), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT41), .ZN(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI22_X1  g402(.A1(new_n555), .A2(new_n596), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G190gat), .B(G218gat), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT94), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n606), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n603), .A2(new_n601), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n604), .B1(new_n598), .B2(new_n599), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n607), .B1(new_n617), .B2(new_n611), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n616), .B1(new_n613), .B2(new_n618), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G57gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(G64gat), .ZN(new_n623));
  INV_X1    g422(.A(G64gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(G57gat), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT9), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(G71gat), .A2(G78gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT90), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(new_n622), .B2(G64gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n622), .A2(G64gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n624), .A2(KEYINPUT90), .A3(G57gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT9), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n628), .B1(new_n627), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT92), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n629), .A2(new_n626), .B1(new_n635), .B2(new_n637), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT92), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n643), .A3(KEYINPUT21), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n644), .B1(new_n556), .B2(new_n557), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(new_n337), .ZN(new_n646));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT91), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n641), .A2(KEYINPUT21), .ZN(new_n652));
  XNOR2_X1  g451(.A(G127gat), .B(G155gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G211gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n646), .A2(new_n650), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n651), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n651), .B2(new_n656), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n590), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT95), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n630), .A2(new_n661), .A3(new_n638), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n593), .B2(new_n594), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n589), .A2(new_n592), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n660), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n641), .A2(new_n665), .A3(new_n666), .A4(new_n661), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n663), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n640), .A2(new_n643), .A3(new_n595), .A4(KEYINPUT10), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(G230gat), .A2(G233gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n663), .A2(new_n667), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(G230gat), .A3(G233gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G204gat), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT96), .B(G176gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n673), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT97), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT97), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n673), .A2(new_n675), .A3(new_n682), .A4(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n673), .A2(new_n675), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n679), .B(KEYINPUT98), .Z(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n621), .A2(new_n659), .A3(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n502), .A2(new_n585), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n303), .B(KEYINPUT99), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g494(.A(KEYINPUT16), .B(G8gat), .Z(new_n696));
  NAND3_X1  g495(.A1(new_n691), .A2(new_n378), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  INV_X1    g499(.A(new_n502), .ZN(new_n701));
  INV_X1    g500(.A(new_n690), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n584), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G8gat), .B1(new_n703), .B2(new_n379), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n699), .A2(new_n700), .A3(new_n704), .ZN(G1325gat));
  XNOR2_X1  g504(.A(new_n489), .B(KEYINPUT100), .ZN(new_n706));
  OAI21_X1  g505(.A(G15gat), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n531), .A3(new_n493), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n707), .A2(KEYINPUT101), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1326gat));
  INV_X1    g512(.A(new_n491), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n691), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  INV_X1    g516(.A(new_n659), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n689), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n621), .ZN(new_n720));
  AND4_X1   g519(.A1(new_n501), .A2(new_n500), .A3(new_n584), .A4(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(G29gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n722), .A3(new_n693), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n621), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n500), .A2(new_n501), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n619), .A2(new_n620), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n498), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n727), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n719), .A2(new_n585), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n729), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G29gat), .B1(new_n734), .B2(new_n692), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n723), .A2(new_n725), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n726), .A2(new_n735), .A3(new_n736), .ZN(G1328gat));
  INV_X1    g536(.A(new_n721), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n738), .A2(G36gat), .A3(new_n379), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n734), .B2(new_n379), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(G1329gat));
  AND3_X1   g543(.A1(new_n721), .A2(new_n493), .A3(new_n526), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n526), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n734), .B2(new_n489), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(KEYINPUT47), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n706), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n729), .A2(new_n732), .A3(new_n750), .A4(new_n733), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n751), .A2(KEYINPUT103), .A3(new_n747), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT103), .B1(new_n751), .B2(new_n747), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n752), .A2(new_n753), .A3(new_n745), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n749), .B1(new_n754), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n491), .A2(G50gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n721), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n729), .A2(new_n732), .A3(new_n714), .A4(new_n733), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G50gat), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n760), .B(new_n762), .C1(new_n759), .C2(new_n758), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n758), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT104), .B1(new_n764), .B2(new_n756), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n761), .A2(G50gat), .B1(new_n721), .B2(new_n757), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT48), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n763), .B1(new_n765), .B2(new_n768), .ZN(G1331gat));
  NAND2_X1  g568(.A1(new_n585), .A2(new_n688), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n770), .A2(new_n718), .A3(new_n730), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n498), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n693), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g573(.A(new_n379), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT106), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1333gat));
  NAND2_X1  g578(.A1(new_n772), .A2(new_n750), .ZN(new_n780));
  INV_X1    g579(.A(new_n493), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(G71gat), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n780), .A2(G71gat), .B1(new_n772), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n772), .A2(new_n714), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT107), .B(G78gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1335gat));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n659), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n729), .A2(new_n732), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n692), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n584), .B(new_n659), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n498), .A2(new_n730), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n795), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n498), .A2(new_n730), .A3(new_n797), .A4(new_n793), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n688), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n693), .A2(new_n205), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n790), .B1(new_n799), .B2(new_n800), .ZN(G1336gat));
  OAI21_X1  g600(.A(G92gat), .B1(new_n789), .B2(new_n379), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n796), .A2(new_n798), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n688), .A2(new_n368), .A3(new_n378), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT109), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT52), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n802), .B(new_n808), .C1(new_n803), .C2(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1337gat));
  NAND4_X1  g609(.A1(new_n729), .A2(new_n732), .A3(new_n750), .A4(new_n788), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT110), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G99gat), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n811), .A2(KEYINPUT110), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n781), .A2(G99gat), .ZN(new_n815));
  OAI22_X1  g614(.A1(new_n813), .A2(new_n814), .B1(new_n799), .B2(new_n815), .ZN(G1338gat));
  NOR2_X1   g615(.A1(new_n491), .A2(G106gat), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n796), .A2(new_n688), .A3(new_n798), .A4(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(KEYINPUT112), .ZN(new_n819));
  XNOR2_X1  g618(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n820));
  XOR2_X1   g619(.A(KEYINPUT111), .B(G106gat), .Z(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n789), .B2(new_n491), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n820), .B1(new_n819), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(G1339gat));
  NOR3_X1   g624(.A1(new_n714), .A2(new_n378), .A3(new_n781), .ZN(new_n826));
  INV_X1    g625(.A(new_n672), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n669), .A2(new_n827), .A3(new_n670), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n669), .A2(new_n670), .A3(KEYINPUT114), .A4(new_n827), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n830), .A2(new_n673), .A3(KEYINPUT54), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n827), .B1(new_n669), .B2(new_n670), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n679), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n832), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n684), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n578), .B2(new_n583), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n567), .A2(new_n570), .A3(new_n577), .ZN(new_n842));
  INV_X1    g641(.A(new_n575), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n562), .B1(new_n560), .B2(new_n561), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n551), .A2(new_n553), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n842), .A2(new_n688), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n621), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n840), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n730), .A2(new_n850), .A3(new_n846), .A4(new_n842), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n659), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n690), .A2(new_n584), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n693), .B(new_n826), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G113gat), .B1(new_n854), .B2(new_n585), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT115), .Z(new_n856));
  XOR2_X1   g655(.A(new_n854), .B(KEYINPUT116), .Z(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n213), .A3(new_n584), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(G1340gat));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n214), .A3(new_n688), .ZN(new_n860));
  OAI21_X1  g659(.A(G120gat), .B1(new_n854), .B2(new_n689), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1341gat));
  NOR2_X1   g661(.A1(new_n854), .A2(new_n718), .ZN(new_n863));
  NOR2_X1   g662(.A1(KEYINPUT117), .A2(G127gat), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT118), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n863), .B(new_n865), .ZN(G1342gat));
  NOR2_X1   g665(.A1(new_n854), .A2(new_n621), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT119), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n867), .A2(new_n868), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(G134gat), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n870), .B(new_n872), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n874), .B(new_n714), .C1(new_n852), .C2(new_n853), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n693), .A2(new_n379), .A3(new_n489), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n840), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n838), .A2(new_n684), .A3(KEYINPUT120), .A4(new_n839), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n584), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n730), .B1(new_n880), .B2(new_n847), .ZN(new_n881));
  AND4_X1   g680(.A1(new_n730), .A2(new_n850), .A3(new_n846), .A4(new_n842), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n718), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n702), .A2(new_n585), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n491), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n875), .B(new_n876), .C1(new_n885), .C2(new_n874), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886), .B2(new_n585), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT58), .B1(new_n887), .B2(KEYINPUT123), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n706), .A2(new_n714), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n852), .A2(new_n853), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n692), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n584), .A2(new_n246), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT122), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n891), .A2(new_n379), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n887), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n888), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n896), .B(new_n887), .C1(KEYINPUT123), .C2(KEYINPUT58), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(G1344gat));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n874), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT57), .B1(new_n892), .B2(new_n491), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n688), .A3(new_n876), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n905), .B2(G148gat), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n886), .A2(new_n689), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(KEYINPUT59), .A3(new_n247), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n379), .A3(new_n893), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n688), .A2(new_n247), .ZN(new_n910));
  OAI22_X1  g709(.A1(new_n906), .A2(new_n908), .B1(new_n909), .B2(new_n910), .ZN(G1345gat));
  OAI21_X1  g710(.A(G155gat), .B1(new_n886), .B2(new_n718), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n718), .A2(G155gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n886), .B2(new_n621), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n621), .A2(G162gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n909), .B2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n892), .A2(new_n693), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n714), .A2(new_n379), .A3(new_n781), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n585), .ZN(new_n923));
  NAND2_X1  g722(.A1(KEYINPUT125), .A2(G169gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g724(.A(KEYINPUT125), .B(G169gat), .Z(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n923), .B2(new_n926), .ZN(G1348gat));
  INV_X1    g726(.A(new_n922), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n688), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n343), .A2(new_n345), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n928), .A2(new_n931), .A3(new_n659), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n337), .B1(new_n922), .B2(new_n718), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n934), .B(new_n935), .ZN(G1350gat));
  NOR2_X1   g735(.A1(new_n922), .A2(new_n621), .ZN(new_n937));
  NAND2_X1  g736(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g738(.A(KEYINPUT61), .B(G190gat), .Z(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n937), .B2(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n889), .A2(new_n379), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n920), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n584), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n750), .A2(new_n693), .A3(new_n379), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n904), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n585), .A2(new_n574), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1352gat));
  XOR2_X1   g748(.A(KEYINPUT126), .B(G204gat), .Z(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n943), .A2(new_n689), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n904), .A2(new_n688), .A3(new_n946), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n950), .B2(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n944), .A2(new_n310), .A3(new_n659), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n904), .A2(new_n659), .A3(new_n946), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  NAND4_X1  g759(.A1(new_n904), .A2(G218gat), .A3(new_n730), .A4(new_n946), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n311), .B1(new_n943), .B2(new_n621), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n961), .A2(new_n965), .A3(new_n962), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1355gat));
endmodule


