//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n607, new_n608, new_n609, new_n610,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n193), .A2(G227), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n192), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT75), .A3(G104), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n196), .A2(KEYINPUT75), .A3(KEYINPUT3), .A4(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G107), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G101), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n196), .A2(G104), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(new_n203), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n211), .B1(new_n214), .B2(KEYINPUT1), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n206), .A2(new_n210), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT10), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n209), .B1(new_n201), .B2(new_n205), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT77), .A3(new_n220), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n225), .ZN(new_n228));
  INV_X1    g042(.A(new_n217), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT1), .B1(new_n215), .B2(G146), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n214), .A2(KEYINPUT66), .A3(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(G128), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n219), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n229), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT10), .B1(new_n228), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n227), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G137), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G134), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT11), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(G134), .B2(new_n239), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n244), .A2(KEYINPUT11), .A3(G137), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n241), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT11), .B1(new_n244), .B2(G137), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n242), .A2(new_n239), .A3(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(new_n241), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n201), .A2(new_n203), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT76), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G101), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n204), .B1(new_n199), .B2(new_n200), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT76), .B1(new_n258), .B2(new_n207), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n201), .B2(new_n205), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n258), .A2(new_n207), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT0), .B(G128), .Z(new_n264));
  OR2_X1    g078(.A1(new_n264), .A2(new_n219), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n219), .A2(new_n266), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n263), .A2(new_n260), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n238), .A2(new_n254), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n254), .B1(new_n238), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n195), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n238), .A2(new_n254), .A3(new_n269), .ZN(new_n273));
  INV_X1    g087(.A(new_n195), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n223), .A2(new_n226), .B1(new_n236), .B2(new_n228), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT12), .B1(new_n253), .B2(KEYINPUT78), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n275), .A2(new_n254), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n276), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n225), .A2(KEYINPUT77), .A3(new_n220), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT77), .B1(new_n225), .B2(new_n220), .ZN(new_n280));
  OAI21_X1  g094(.A(G128), .B1(new_n230), .B2(new_n231), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT66), .B1(new_n214), .B2(KEYINPUT1), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n235), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n217), .ZN(new_n284));
  OAI22_X1  g098(.A1(new_n279), .A2(new_n280), .B1(new_n284), .B2(new_n225), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n278), .B1(new_n285), .B2(new_n253), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n273), .B(new_n274), .C1(new_n277), .C2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(G902), .B1(new_n272), .B2(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(KEYINPUT79), .B(G469), .Z(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n273), .B1(new_n277), .B2(new_n286), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n195), .B(KEYINPUT74), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n227), .A2(new_n237), .B1(new_n262), .B2(new_n268), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n195), .B1(new_n294), .B2(new_n254), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n238), .A2(new_n269), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n253), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n291), .A2(new_n293), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G469), .B1(new_n298), .B2(G902), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n191), .B1(new_n290), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(G116), .B(G119), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT5), .ZN(new_n302));
  INV_X1    g116(.A(G116), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n303), .A2(KEYINPUT5), .A3(G119), .ZN(new_n304));
  INV_X1    g118(.A(G113), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT2), .B(G113), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n302), .A2(new_n306), .B1(new_n308), .B2(new_n301), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n309), .A2(new_n225), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n301), .B(new_n307), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n263), .B2(new_n260), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n310), .B1(new_n262), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(G110), .B(G122), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(new_n314), .B(KEYINPUT80), .Z(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT6), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT81), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n262), .A2(new_n312), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n317), .B1(new_n321), .B2(new_n310), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT6), .A4(new_n315), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n267), .B1(new_n264), .B2(new_n219), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G125), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n236), .B2(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n193), .A2(G224), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n313), .A2(KEYINPUT6), .A3(new_n318), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n320), .A2(new_n324), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT82), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n328), .B1(new_n332), .B2(KEYINPUT7), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n332), .B2(KEYINPUT7), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n327), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n327), .A2(KEYINPUT7), .A3(new_n328), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n314), .B(KEYINPUT8), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n309), .A2(new_n225), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n310), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(G902), .B1(new_n340), .B2(new_n315), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n331), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(G210), .B1(G237), .B2(G902), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n331), .A2(new_n341), .A3(new_n343), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G214), .B1(G237), .B2(G902), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n300), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G475), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT16), .ZN(new_n351));
  INV_X1    g165(.A(G125), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G140), .ZN(new_n353));
  INV_X1    g167(.A(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G125), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n355), .A3(KEYINPUT71), .ZN(new_n356));
  OR3_X1    g170(.A1(new_n354), .A2(KEYINPUT71), .A3(G125), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n351), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(new_n354), .A3(G125), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT72), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(G146), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G237), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n193), .A3(G214), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n215), .ZN(new_n366));
  NOR2_X1   g180(.A1(G237), .A2(G953), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(G143), .A3(G214), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G131), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT17), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(new_n251), .A3(new_n368), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n360), .B(KEYINPUT72), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n213), .B1(new_n374), .B2(new_n358), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n369), .A2(KEYINPUT17), .A3(G131), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n363), .A2(new_n373), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n366), .A2(new_n368), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n213), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n356), .A2(new_n357), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(new_n213), .ZN(new_n383));
  INV_X1    g197(.A(new_n378), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n369), .A2(KEYINPUT83), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT83), .B1(new_n369), .B2(new_n384), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n379), .B(new_n383), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n377), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n202), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n377), .A2(new_n387), .A3(new_n390), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n350), .B1(new_n394), .B2(new_n190), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n350), .A2(new_n190), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT84), .ZN(new_n398));
  INV_X1    g212(.A(new_n393), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n370), .A2(new_n372), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n380), .A2(KEYINPUT19), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n382), .B2(KEYINPUT19), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n363), .B(new_n400), .C1(G146), .C2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n390), .B1(new_n403), .B2(new_n387), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n398), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n387), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n391), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(new_n408), .B2(new_n393), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n405), .B1(new_n409), .B2(KEYINPUT20), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n393), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n406), .A3(new_n412), .A4(new_n398), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n193), .A2(G952), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(G234), .B2(G237), .ZN(new_n416));
  INV_X1    g230(.A(G234), .ZN(new_n417));
  OAI211_X1 g231(.A(G902), .B(G953), .C1(new_n417), .C2(new_n364), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n418), .B(KEYINPUT88), .Z(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT21), .B(G898), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n303), .B2(G122), .ZN(new_n426));
  INV_X1    g240(.A(G122), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT86), .A3(G116), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n303), .A2(G122), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n196), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n196), .B1(new_n429), .B2(new_n430), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n424), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n433), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT87), .A3(new_n431), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT13), .B1(new_n211), .B2(G143), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n244), .ZN(new_n438));
  XNOR2_X1  g252(.A(G128), .B(G143), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n434), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n430), .B(KEYINPUT14), .ZN(new_n442));
  INV_X1    g256(.A(new_n429), .ZN(new_n443));
  OAI21_X1  g257(.A(G107), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n439), .B(new_n244), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n431), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G217), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n188), .A2(new_n447), .A3(G953), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n441), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n441), .B2(new_n446), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n190), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G478), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT15), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n441), .A2(new_n446), .ZN(new_n455));
  INV_X1    g269(.A(new_n448), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n441), .A2(new_n446), .A3(new_n448), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n453), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n190), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  AND4_X1   g276(.A1(new_n396), .A2(new_n414), .A3(new_n423), .A4(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n349), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT73), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n367), .A2(G210), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT27), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT26), .B(G101), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT67), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT28), .ZN(new_n472));
  AOI211_X1 g286(.A(G131), .B(new_n240), .C1(new_n248), .C2(new_n249), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n251), .B1(new_n250), .B2(new_n241), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n325), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT65), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n239), .B2(G134), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT64), .B1(new_n244), .B2(G137), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT64), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n239), .A3(G134), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n244), .A2(KEYINPUT65), .A3(G137), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n477), .A2(new_n478), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G131), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n252), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n475), .B1(new_n236), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n311), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n475), .B(new_n311), .C1(new_n236), .C2(new_n484), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n472), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n483), .A2(new_n252), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n490), .A2(new_n284), .B1(new_n253), .B2(new_n325), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT28), .B1(new_n491), .B2(new_n311), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n471), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n475), .B(KEYINPUT30), .C1(new_n236), .C2(new_n484), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n486), .B(new_n494), .C1(new_n491), .C2(KEYINPUT30), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n488), .A2(new_n469), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n495), .A2(KEYINPUT31), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT31), .B1(new_n495), .B2(new_n496), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT68), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(G472), .A2(G902), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n493), .B(KEYINPUT68), .C1(new_n497), .C2(new_n498), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT69), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT32), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n501), .A2(new_n507), .A3(new_n502), .A4(new_n503), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n495), .A2(new_n488), .ZN(new_n510));
  INV_X1    g324(.A(new_n469), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n489), .A2(new_n471), .A3(new_n492), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n513), .A2(KEYINPUT29), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n489), .A2(new_n492), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT29), .A3(new_n469), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n190), .ZN(new_n518));
  OAI21_X1  g332(.A(G472), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n501), .A2(KEYINPUT32), .A3(new_n502), .A4(new_n503), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n509), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n447), .B1(G234), .B2(new_n190), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT22), .B(G137), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n187), .A2(new_n417), .A3(G953), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT23), .B1(new_n211), .B2(G119), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT70), .B1(new_n211), .B2(G119), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n211), .B(G119), .C1(KEYINPUT70), .C2(KEYINPUT23), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(G119), .B(G128), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT24), .B(G110), .Z(new_n535));
  OAI22_X1  g349(.A1(new_n533), .A2(G110), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n363), .A2(new_n381), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n533), .A2(G110), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n534), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n363), .B2(new_n375), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n528), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n542), .ZN(new_n544));
  INV_X1    g358(.A(new_n528), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n537), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n525), .B1(new_n547), .B2(G902), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n543), .A2(new_n546), .A3(KEYINPUT25), .A4(new_n190), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n524), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n547), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n523), .A2(G902), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n465), .B1(new_n522), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n553), .ZN(new_n555));
  AOI211_X1 g369(.A(KEYINPUT73), .B(new_n555), .C1(new_n509), .C2(new_n521), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n464), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT89), .B(G101), .Z(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(G3));
  NAND2_X1  g373(.A1(new_n300), .A2(new_n553), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n501), .A2(new_n190), .A3(new_n503), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G472), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n505), .A2(new_n563), .A3(new_n508), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n565), .A3(KEYINPUT90), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT90), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n560), .B2(new_n564), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n347), .A2(new_n348), .A3(new_n423), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n395), .B1(new_n410), .B2(new_n413), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n459), .A2(KEYINPUT33), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT33), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n457), .A2(new_n573), .A3(new_n458), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(G478), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n459), .A2(new_n452), .A3(new_n190), .ZN(new_n576));
  NAND2_X1  g390(.A1(G478), .A2(G902), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n571), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n569), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n566), .A2(new_n568), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT34), .B(G104), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G6));
  INV_X1    g398(.A(new_n569), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n405), .A2(KEYINPUT20), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n411), .A2(new_n412), .A3(new_n398), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n395), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n454), .A2(new_n461), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n566), .A2(new_n568), .A3(new_n585), .A4(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT35), .B(G107), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G9));
  OAI21_X1  g408(.A(KEYINPUT91), .B1(new_n538), .B2(new_n542), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT91), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n544), .A2(new_n596), .A3(new_n537), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n598), .B1(new_n595), .B2(new_n597), .ZN(new_n600));
  INV_X1    g414(.A(new_n552), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n550), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n349), .A2(new_n565), .A3(new_n463), .A4(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT37), .B(G110), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G12));
  XOR2_X1   g420(.A(KEYINPUT92), .B(G900), .Z(new_n607));
  AOI21_X1  g421(.A(new_n416), .B1(new_n420), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n590), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n522), .A2(new_n349), .A3(new_n603), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G128), .ZN(G30));
  AND2_X1   g425(.A1(new_n495), .A2(new_n496), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n487), .A2(new_n488), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(new_n471), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n614), .B2(G902), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n520), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n509), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(KEYINPUT94), .Z(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n347), .B(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n462), .B1(new_n414), .B2(new_n396), .ZN(new_n623));
  INV_X1    g437(.A(new_n348), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n603), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n608), .B(KEYINPUT39), .Z(new_n626));
  NAND2_X1  g440(.A1(new_n300), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n623), .B(new_n625), .C1(new_n627), .C2(KEYINPUT40), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(KEYINPUT40), .B2(new_n627), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n618), .A2(new_n622), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G143), .ZN(G45));
  NOR3_X1   g445(.A1(new_n570), .A2(new_n578), .A3(new_n608), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n522), .A2(new_n349), .A3(new_n603), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G146), .ZN(G48));
  AOI21_X1  g448(.A(new_n555), .B1(new_n509), .B2(new_n521), .ZN(new_n635));
  INV_X1    g449(.A(new_n191), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n272), .A2(new_n287), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n190), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT95), .B1(new_n638), .B2(G469), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT95), .ZN(new_n640));
  INV_X1    g454(.A(G469), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n288), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n636), .B(new_n290), .C1(new_n639), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT96), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n638), .A2(KEYINPUT95), .A3(G469), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n640), .B1(new_n288), .B2(new_n641), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n647), .A2(new_n648), .A3(new_n636), .A4(new_n290), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n635), .A2(new_n581), .A3(new_n644), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT41), .B(G113), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G15));
  NOR2_X1   g466(.A1(new_n569), .A2(new_n590), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n635), .A2(new_n653), .A3(new_n644), .A4(new_n649), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G116), .ZN(G18));
  NAND2_X1  g469(.A1(new_n463), .A2(new_n603), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n509), .B2(new_n521), .ZN(new_n657));
  INV_X1    g471(.A(new_n347), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n624), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n657), .A2(new_n644), .A3(new_n659), .A4(new_n649), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G119), .ZN(G21));
  AND3_X1   g475(.A1(new_n331), .A2(new_n341), .A3(new_n343), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n343), .B1(new_n331), .B2(new_n341), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n623), .B(new_n348), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n347), .A2(KEYINPUT97), .A3(new_n348), .A4(new_n623), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n499), .A2(new_n502), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n423), .A2(new_n563), .A3(new_n553), .A4(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n668), .A2(new_n649), .A3(new_n644), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G122), .ZN(G24));
  AND4_X1   g486(.A1(new_n563), .A2(new_n632), .A3(new_n603), .A4(new_n669), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n644), .A2(new_n673), .A3(new_n659), .A4(new_n649), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G125), .ZN(G27));
  NAND2_X1  g489(.A1(new_n299), .A2(KEYINPUT98), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n641), .A2(KEYINPUT98), .A3(G902), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n298), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n290), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n345), .A2(new_n348), .A3(new_n346), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n636), .A3(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n504), .A2(new_n506), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n519), .A2(new_n520), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n553), .B(new_n632), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT42), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n288), .A2(new_n289), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n676), .B2(new_n678), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n689), .A2(new_n191), .A3(new_n681), .ZN(new_n690));
  INV_X1    g504(.A(new_n632), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(KEYINPUT42), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n635), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n251), .ZN(G33));
  NAND3_X1  g509(.A1(new_n690), .A2(new_n635), .A3(new_n609), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G134), .ZN(G36));
  XOR2_X1   g511(.A(new_n681), .B(KEYINPUT104), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n579), .A2(new_n570), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n703));
  AOI22_X1  g517(.A1(new_n579), .A2(new_n570), .B1(new_n703), .B2(KEYINPUT43), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(KEYINPUT103), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n701), .B2(new_n704), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n550), .A2(new_n602), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n565), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n712), .B1(new_n709), .B2(new_n711), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n698), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(G469), .B1(new_n298), .B2(KEYINPUT45), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n291), .A2(new_n293), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n295), .A2(new_n297), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n720));
  OR3_X1    g534(.A1(new_n719), .A2(KEYINPUT99), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT99), .B1(new_n719), .B2(new_n720), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n716), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n641), .A2(new_n190), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT100), .B1(new_n725), .B2(KEYINPUT46), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n688), .B1(new_n725), .B2(KEYINPUT46), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT100), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n728), .B(new_n729), .C1(new_n723), .C2(new_n724), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n726), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n636), .A3(new_n626), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT101), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n731), .A2(KEYINPUT101), .A3(new_n636), .A4(new_n626), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n715), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT105), .B(G137), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G39));
  NOR3_X1   g552(.A1(new_n522), .A2(new_n691), .A3(new_n553), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n682), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n731), .A2(new_n636), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n731), .A2(KEYINPUT47), .A3(new_n636), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT106), .B(G140), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G42));
  NAND2_X1  g561(.A1(new_n647), .A2(new_n290), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT107), .Z(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(KEYINPUT49), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(KEYINPUT108), .Z(new_n751));
  XNOR2_X1  g565(.A(new_n617), .B(KEYINPUT94), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n553), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n749), .A2(KEYINPUT49), .ZN(new_n755));
  NOR4_X1   g569(.A1(new_n622), .A2(new_n191), .A3(new_n624), .A4(new_n699), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n751), .A2(new_n754), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n571), .A2(new_n462), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n566), .A2(new_n568), .A3(new_n585), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n604), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n557), .A2(new_n582), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n557), .A2(KEYINPUT109), .A3(new_n582), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n690), .A2(new_n673), .ZN(new_n766));
  INV_X1    g580(.A(new_n608), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n588), .A2(new_n462), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n710), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n522), .A2(new_n300), .A3(new_n682), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n690), .A2(new_n635), .A3(new_n609), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT110), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n769), .A2(new_n300), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n774), .B1(new_n509), .B2(new_n521), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n775), .A2(new_n682), .B1(new_n690), .B2(new_n673), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n696), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n650), .A2(new_n671), .A3(new_n654), .A4(new_n660), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n694), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n764), .A2(new_n765), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n603), .A2(new_n608), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n299), .A2(KEYINPUT98), .B1(new_n298), .B2(new_n677), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n784), .B(new_n636), .C1(new_n785), .C2(new_n688), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT112), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n680), .A2(new_n788), .A3(new_n636), .A4(new_n784), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n666), .A2(new_n667), .B1(new_n509), .B2(new_n616), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n674), .A2(new_n610), .A3(new_n633), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n783), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n674), .A2(new_n610), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n790), .A2(new_n791), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT52), .A4(new_n633), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n758), .B1(new_n782), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n779), .A2(new_n781), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n557), .A2(KEYINPUT109), .A3(new_n582), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT109), .B1(new_n557), .B2(new_n582), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n803), .A2(new_n804), .A3(new_n761), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n795), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n783), .B1(new_n790), .B2(new_n791), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n674), .A2(new_n610), .A3(KEYINPUT111), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n633), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n794), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n802), .A2(new_n805), .A3(new_n811), .A4(KEYINPUT53), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n800), .A2(new_n801), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n782), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n794), .A2(new_n798), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(KEYINPUT113), .A3(KEYINPUT53), .A4(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n802), .A2(new_n805), .A3(KEYINPUT53), .A4(new_n815), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n811), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n758), .B1(new_n820), .B2(new_n782), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n816), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n813), .B1(new_n822), .B2(KEYINPUT54), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n644), .A2(new_n649), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(KEYINPUT116), .A3(new_n682), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n644), .A2(new_n649), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(new_n681), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n416), .B1(new_n701), .B2(new_n704), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT117), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n829), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n563), .A2(new_n669), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n603), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n824), .A2(new_n624), .A3(new_n621), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n553), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n831), .B2(new_n832), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n824), .A2(KEYINPUT115), .A3(new_n624), .A4(new_n621), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n843), .A2(KEYINPUT50), .A3(new_n845), .A4(new_n846), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n754), .A2(new_n416), .A3(new_n829), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n571), .A2(new_n579), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n849), .A2(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n743), .A2(new_n744), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n749), .A2(new_n636), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n698), .B(new_n845), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n840), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT48), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n553), .B1(new_n684), .B2(new_n685), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n838), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n415), .B(KEYINPUT118), .Z(new_n864));
  NOR3_X1   g678(.A1(new_n827), .A2(new_n624), .A3(new_n658), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n845), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n754), .A2(new_n829), .A3(new_n416), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n866), .B1(new_n867), .B2(new_n580), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT119), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n870), .B(new_n866), .C1(new_n867), .C2(new_n580), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n860), .A2(new_n863), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n840), .A2(new_n853), .A3(KEYINPUT51), .A4(new_n856), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n838), .A2(KEYINPUT48), .A3(new_n862), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n823), .A2(new_n859), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(G952), .A2(G953), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n757), .B1(new_n876), .B2(new_n877), .ZN(G75));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n800), .A2(new_n812), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(G902), .ZN(new_n881));
  INV_X1    g695(.A(G210), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n320), .A2(new_n324), .A3(new_n330), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n329), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT55), .Z(new_n886));
  AND2_X1   g700(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n883), .A2(new_n886), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n193), .A2(G952), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G51));
  NAND3_X1  g704(.A1(new_n800), .A2(new_n801), .A3(new_n812), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT120), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n800), .A2(new_n812), .A3(new_n893), .A4(new_n801), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n880), .A2(KEYINPUT54), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n724), .B(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n637), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n880), .A2(G902), .A3(new_n723), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n889), .B1(new_n899), .B2(new_n900), .ZN(G54));
  INV_X1    g715(.A(new_n411), .ZN(new_n902));
  NAND2_X1  g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(new_n881), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n889), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n881), .A2(new_n902), .A3(new_n903), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(G60));
  AND2_X1   g722(.A1(new_n572), .A2(new_n574), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n577), .B(KEYINPUT59), .Z(new_n910));
  OAI21_X1  g724(.A(new_n909), .B1(new_n823), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n889), .B1(new_n896), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT60), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n800), .B2(new_n812), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(new_n551), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n599), .A2(new_n600), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n889), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT121), .B1(new_n917), .B2(new_n920), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n918), .B(new_n921), .C1(new_n923), .C2(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(G66));
  INV_X1    g741(.A(new_n421), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n193), .B1(new_n928), .B2(G224), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n762), .A2(new_n763), .ZN(new_n930));
  INV_X1    g744(.A(new_n761), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n765), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n780), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n934), .B2(new_n193), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n884), .B1(G898), .B2(new_n193), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n935), .B(new_n936), .Z(G69));
  AOI21_X1  g751(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n807), .A2(new_n633), .A3(new_n809), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n734), .A2(new_n735), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n861), .B1(new_n666), .B2(new_n667), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n687), .A2(new_n693), .A3(new_n696), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n745), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n715), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n942), .A2(new_n944), .A3(new_n193), .A4(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n494), .B1(new_n491), .B2(KEYINPUT30), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT122), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n402), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(G900), .B2(G953), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n947), .A2(KEYINPUT126), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n950), .B(KEYINPUT123), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n630), .A2(new_n633), .A3(new_n809), .A4(new_n807), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT62), .Z(new_n960));
  INV_X1    g774(.A(new_n745), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n554), .A2(new_n556), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n580), .B1(new_n571), .B2(new_n462), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n682), .A2(new_n300), .A3(new_n626), .A4(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT124), .B1(new_n946), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT124), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n736), .A2(new_n968), .A3(new_n965), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n960), .B(new_n961), .C1(new_n967), .C2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n958), .B1(new_n970), .B2(new_n193), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n938), .B1(new_n956), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n193), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(KEYINPUT125), .A3(new_n957), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n938), .B1(new_n947), .B2(new_n951), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n971), .A2(KEYINPUT125), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(G72));
  NAND4_X1  g792(.A1(new_n942), .A2(new_n944), .A3(new_n946), .A4(new_n933), .ZN(new_n979));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(KEYINPUT127), .A3(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(new_n488), .A3(new_n511), .A4(new_n495), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT127), .B1(new_n979), .B2(new_n981), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n905), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n510), .A2(new_n469), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n946), .A2(KEYINPUT124), .A3(new_n966), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n968), .B1(new_n736), .B2(new_n965), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n745), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n989), .A2(new_n933), .A3(new_n960), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n986), .B1(new_n990), .B2(new_n981), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n513), .A2(new_n612), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n822), .A2(new_n981), .A3(new_n992), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n985), .A2(new_n991), .A3(new_n993), .ZN(G57));
endmodule


