//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n561, new_n562, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n615, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT68), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n460), .B1(new_n449), .B2(new_n456), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g037(.A(G113), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT70), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(G113), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n465), .B(new_n467), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G101), .A3(G2104), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT71), .B1(new_n469), .B2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n469), .A2(G2104), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n475), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G137), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n478), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(new_n468), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(G2105), .A3(new_n479), .ZN(new_n492));
  INV_X1    g067(.A(G124), .ZN(new_n493));
  OAI221_X1 g068(.A(new_n488), .B1(new_n482), .B2(new_n489), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  OR3_X1    g071(.A1(new_n496), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(new_n471), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n491), .A2(G138), .A3(new_n475), .A4(new_n479), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(KEYINPUT4), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(new_n475), .B2(G114), .ZN(new_n501));
  NOR2_X1   g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT72), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n502), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n504), .A2(new_n506), .A3(new_n507), .A4(G2104), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n491), .A2(G126), .A3(G2105), .A4(new_n479), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n500), .A2(new_n511), .ZN(G164));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(KEYINPUT73), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(KEYINPUT6), .A3(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n514), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n520), .A2(G651), .B1(G50), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n518), .B1(new_n523), .B2(new_n525), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT74), .B(G88), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND2_X1  g107(.A1(new_n528), .A2(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n526), .A2(G51), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n515), .A2(new_n517), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n537), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n533), .A2(new_n535), .A3(new_n536), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  XNOR2_X1  g115(.A(KEYINPUT76), .B(G52), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n528), .A2(G90), .B1(new_n526), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT77), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n537), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT75), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n537), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n522), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n526), .A2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n523), .A2(new_n525), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n537), .A2(new_n552), .A3(G81), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n551), .A2(new_n553), .A3(KEYINPUT78), .ZN(new_n554));
  AOI21_X1  g129(.A(KEYINPUT78), .B1(new_n551), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n526), .B2(G53), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n526), .A2(new_n564), .A3(G53), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n566), .A2(new_n567), .B1(G91), .B2(new_n528), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n518), .A2(KEYINPUT79), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n515), .A2(new_n517), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(G65), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n522), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n568), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n528), .A2(G91), .ZN(new_n578));
  INV_X1    g153(.A(new_n567), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n565), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT80), .B1(new_n580), .B2(new_n574), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G299));
  NAND2_X1  g157(.A1(new_n528), .A2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n526), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n537), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  AOI22_X1  g161(.A1(new_n537), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n522), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n526), .A2(G48), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n528), .A2(G86), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G305));
  XOR2_X1   g166(.A(KEYINPUT81), .B(G47), .Z(new_n592));
  NAND2_X1  g167(.A1(new_n526), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n537), .A2(new_n552), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n537), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI221_X1 g171(.A(new_n593), .B1(new_n594), .B2(new_n595), .C1(new_n596), .C2(new_n522), .ZN(G290));
  NAND3_X1  g172(.A1(new_n528), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n598), .A2(new_n601), .B1(G54), .B2(new_n526), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n569), .A2(G66), .A3(new_n571), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT82), .Z(new_n605));
  OAI21_X1  g180(.A(G651), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G171), .B2(new_n608), .ZN(G284));
  XOR2_X1   g185(.A(G284), .B(KEYINPUT83), .Z(G321));
  INV_X1    g186(.A(G299), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n608), .ZN(new_n613));
  NAND2_X1  g188(.A1(G168), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT84), .Z(G297));
  INV_X1    g191(.A(new_n615), .ZN(G280));
  INV_X1    g192(.A(new_n607), .ZN(new_n618));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G860), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT85), .Z(G148));
  NAND2_X1  g196(.A1(new_n556), .A2(new_n608), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n607), .A2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g200(.A(new_n492), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G123), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n483), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n469), .A2(new_n464), .A3(G2105), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n637), .A2(KEYINPUT87), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n637), .A2(KEYINPUT87), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n632), .B(new_n640), .C1(new_n638), .C2(new_n636), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT88), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2443), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT89), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n652), .B(new_n654), .Z(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(G14), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  AOI21_X1  g236(.A(KEYINPUT18), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n668), .A2(new_n669), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n674), .B1(KEYINPUT20), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n677), .B(new_n678), .C1(KEYINPUT20), .C2(new_n676), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT90), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT91), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(G6), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G305), .B2(G16), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT32), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI211_X1 g268(.A(KEYINPUT32), .B(new_n689), .C1(G305), .C2(G16), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n693), .A2(G1981), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G1981), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n692), .B2(new_n694), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n688), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n688), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n696), .A2(new_n698), .B1(G1976), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n688), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n688), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT94), .B(G1971), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n703), .A2(G1976), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n704), .A2(new_n705), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G25), .ZN(new_n712));
  OAI21_X1  g287(.A(KEYINPUT92), .B1(new_n712), .B2(G29), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n712), .A2(KEYINPUT92), .A3(G29), .ZN(new_n714));
  OR2_X1    g289(.A1(G95), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT93), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n626), .A2(G119), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n483), .A2(G131), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n713), .B(new_n714), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT35), .B(G1991), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n711), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n696), .A2(new_n698), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n703), .A2(G1976), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n728), .A2(new_n710), .A3(new_n709), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(KEYINPUT34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT95), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT95), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n730), .A2(new_n733), .A3(KEYINPUT34), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n688), .A2(G24), .ZN(new_n735));
  INV_X1    g310(.A(G290), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(new_n688), .ZN(new_n737));
  INV_X1    g312(.A(G1986), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n727), .A2(new_n732), .A3(new_n734), .A4(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(KEYINPUT36), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT97), .Z(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n741), .A2(KEYINPUT36), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n740), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(G5), .A2(G16), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G301), .B2(new_n688), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1961), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  NAND2_X1  g325(.A1(G164), .A2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G27), .B2(G29), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n749), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n688), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n688), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT104), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n752), .A2(new_n750), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n722), .B1(new_n761), .B2(G28), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(G28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(KEYINPUT105), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n631), .B2(new_n722), .ZN(new_n767));
  AND2_X1   g342(.A1(KEYINPUT24), .A2(G34), .ZN(new_n768));
  NOR2_X1   g343(.A1(KEYINPUT24), .A2(G34), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n768), .A2(new_n769), .A3(G29), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n485), .B2(G29), .ZN(new_n771));
  INV_X1    g346(.A(G2084), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n767), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n758), .A2(new_n759), .A3(new_n760), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n722), .A2(G35), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G162), .B2(new_n722), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT29), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(G2090), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(G2090), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT101), .B(KEYINPUT26), .ZN(new_n780));
  AND3_X1   g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n491), .A2(G129), .A3(G2105), .A4(new_n479), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n491), .A2(G141), .A3(new_n475), .A4(new_n479), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n475), .A2(G105), .A3(G2104), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT102), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G29), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G29), .B2(G32), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT27), .B(G1996), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n778), .B(new_n779), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n753), .A2(new_n774), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n722), .A2(G26), .ZN(new_n793));
  OR2_X1    g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n795));
  INV_X1    g370(.A(G140), .ZN(new_n796));
  INV_X1    g371(.A(G128), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n795), .B1(new_n482), .B2(new_n796), .C1(new_n492), .C2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n793), .B1(new_n798), .B2(G29), .ZN(new_n799));
  MUX2_X1   g374(.A(new_n793), .B(new_n799), .S(KEYINPUT28), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2067), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G4), .B2(G16), .ZN(new_n803));
  OR3_X1    g378(.A1(new_n802), .A2(G4), .A3(G16), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n803), .B(new_n804), .C1(new_n607), .C2(new_n688), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1348), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n688), .A2(G19), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n556), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1341), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n801), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n688), .A2(KEYINPUT23), .A3(G20), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT23), .ZN(new_n814));
  INV_X1    g389(.A(G20), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(G16), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n813), .B(new_n816), .C1(new_n612), .C2(new_n688), .ZN(new_n817));
  INV_X1    g392(.A(G1956), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n792), .A2(new_n812), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(G115), .A2(G2104), .ZN(new_n821));
  INV_X1    g396(.A(G127), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n471), .B2(new_n822), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n483), .A2(G139), .B1(new_n823), .B2(G2105), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT25), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT100), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n824), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n722), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n722), .B2(G33), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G2072), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n789), .A2(new_n790), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n833), .B(new_n834), .C1(new_n772), .C2(new_n771), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT103), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n820), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n746), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT31), .B(G11), .Z(new_n839));
  AOI21_X1  g414(.A(new_n744), .B1(new_n740), .B2(new_n745), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G311));
  INV_X1    g416(.A(new_n840), .ZN(new_n842));
  INV_X1    g417(.A(new_n839), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n842), .A2(new_n843), .A3(new_n746), .A4(new_n837), .ZN(G150));
  NAND2_X1  g419(.A1(new_n528), .A2(G93), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n526), .A2(G55), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n537), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n845), .B(new_n846), .C1(new_n522), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  OR2_X1    g425(.A1(new_n847), .A2(new_n522), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n556), .A2(new_n845), .A3(new_n851), .A4(new_n846), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n848), .B(new_n550), .C1(new_n554), .C2(new_n555), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n607), .A2(new_n619), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n860));
  AOI21_X1  g435(.A(G860), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n857), .A2(new_n858), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n850), .B1(new_n862), .B2(new_n863), .ZN(G145));
  OAI21_X1  g439(.A(KEYINPUT4), .B1(new_n482), .B2(new_n496), .ZN(new_n865));
  INV_X1    g440(.A(new_n498), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n509), .A2(new_n510), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT107), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n871));
  NAND2_X1  g446(.A1(G164), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n787), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n786), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n786), .A2(new_n875), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n870), .B(new_n872), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n798), .ZN(new_n880));
  INV_X1    g455(.A(new_n798), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n874), .A2(new_n881), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT108), .B1(new_n827), .B2(KEYINPUT100), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G142), .ZN(new_n886));
  NOR2_X1   g461(.A1(G106), .A2(G2105), .ZN(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(new_n475), .B2(G118), .ZN(new_n888));
  OAI22_X1  g463(.A1(new_n482), .A2(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(G130), .B2(new_n626), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(new_n635), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n721), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n829), .B1(new_n883), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n885), .B(new_n892), .C1(new_n894), .C2(new_n827), .ZN(new_n895));
  INV_X1    g470(.A(new_n892), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n874), .A2(new_n881), .A3(new_n878), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n881), .B1(new_n874), .B2(new_n878), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n893), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n827), .B1(new_n899), .B2(KEYINPUT100), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n883), .A2(new_n884), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n902), .A3(KEYINPUT109), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n904), .B(new_n896), .C1(new_n900), .C2(new_n901), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n485), .B(new_n631), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n494), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(KEYINPUT110), .B(G37), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT111), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n910), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n895), .A2(new_n902), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n908), .A2(new_n909), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT40), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT40), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n908), .A2(new_n916), .A3(new_n909), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(G395));
  INV_X1    g493(.A(KEYINPUT113), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n854), .B(new_n623), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n576), .B1(new_n568), .B2(new_n575), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n580), .A2(KEYINPUT80), .A3(new_n574), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n618), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n577), .A2(new_n581), .A3(new_n607), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(KEYINPUT112), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT112), .ZN(new_n930));
  NAND3_X1  g505(.A1(G299), .A2(new_n930), .A3(new_n618), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n924), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT41), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n923), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n919), .A2(new_n920), .ZN(new_n935));
  XNOR2_X1  g510(.A(G303), .B(G288), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n936), .A2(G305), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(G305), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n736), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n736), .B1(new_n937), .B2(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n935), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n929), .A2(new_n931), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n922), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n934), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n934), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n921), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n929), .A2(new_n931), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n933), .B1(new_n948), .B2(KEYINPUT41), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n944), .B1(new_n949), .B2(new_n922), .ZN(new_n950));
  INV_X1    g525(.A(new_n942), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n934), .A2(new_n942), .A3(new_n944), .ZN(new_n953));
  INV_X1    g528(.A(new_n921), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n947), .A2(G868), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n848), .A2(new_n608), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n960), .B2(new_n957), .ZN(G295));
  OAI21_X1  g536(.A(new_n958), .B1(new_n960), .B2(new_n957), .ZN(G331));
  AND3_X1   g537(.A1(G301), .A2(new_n853), .A3(new_n852), .ZN(new_n963));
  AOI21_X1  g538(.A(G301), .B1(new_n852), .B2(new_n853), .ZN(new_n964));
  OAI21_X1  g539(.A(G286), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(G171), .A2(new_n854), .ZN(new_n966));
  NAND3_X1  g541(.A1(G301), .A2(new_n853), .A3(new_n852), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(G168), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n948), .B1(new_n969), .B2(new_n924), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n937), .A2(new_n938), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G290), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n939), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n965), .A2(new_n968), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n927), .A2(new_n928), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT41), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n970), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n943), .A2(new_n968), .A3(new_n965), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n973), .B(new_n979), .C1(new_n969), .C2(new_n949), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n978), .A2(KEYINPUT43), .A3(new_n909), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n969), .B2(new_n949), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n974), .ZN(new_n983));
  INV_X1    g558(.A(G37), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n980), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(new_n986), .B2(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n978), .A2(new_n990), .A3(new_n909), .A4(new_n980), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n988), .A2(new_n994), .ZN(G397));
  INV_X1    g570(.A(new_n787), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(G1996), .ZN(new_n997));
  INV_X1    g572(.A(G2067), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n798), .B(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1996), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n787), .A2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n997), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n720), .B(new_n725), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n500), .B2(new_n511), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n477), .A2(G40), .A3(new_n484), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1011), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(new_n738), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT115), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n1017));
  AND4_X1   g592(.A1(G40), .A2(new_n484), .A3(new_n474), .A4(new_n476), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT45), .B(new_n1006), .C1(new_n500), .C2(new_n511), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1009), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1009), .A2(KEYINPUT116), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n750), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1007), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT50), .B(new_n1006), .C1(new_n500), .C2(new_n511), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1010), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(G1961), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1020), .A2(new_n1025), .A3(G2078), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1026), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(G171), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1032), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1036));
  AOI21_X1  g611(.A(G301), .B1(new_n1036), .B2(new_n1031), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1017), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(G171), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(G301), .A3(new_n1031), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(KEYINPUT54), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1020), .A2(new_n757), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT50), .B1(new_n869), .B2(new_n1006), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1029), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n772), .B(new_n1018), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G286), .A2(G8), .ZN(new_n1048));
  XOR2_X1   g623(.A(new_n1048), .B(KEYINPUT123), .Z(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT124), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT124), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n772), .A2(new_n1030), .B1(new_n1020), .B2(new_n757), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1052), .B(new_n1049), .C1(new_n1053), .C2(new_n1042), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1051), .A2(new_n1054), .A3(KEYINPUT51), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1053), .A2(new_n1049), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT124), .B(new_n1057), .C1(new_n1047), .C2(new_n1050), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1971), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1018), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G2090), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G303), .A2(G8), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(KEYINPUT55), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G305), .A2(G1981), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n588), .A2(new_n697), .A3(new_n589), .A4(new_n590), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(KEYINPUT49), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1007), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1042), .B1(new_n1070), .B2(new_n1018), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT49), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n700), .A2(G1976), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT52), .ZN(new_n1077));
  INV_X1    g652(.A(G1976), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT52), .B1(G288), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1071), .A2(new_n1075), .A3(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1074), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1065), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1061), .B2(G2090), .ZN(new_n1084));
  INV_X1    g659(.A(G2090), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1030), .A2(KEYINPUT117), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(G8), .B(new_n1082), .C1(new_n1087), .C2(new_n1060), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1066), .A2(new_n1081), .A3(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1038), .A2(new_n1041), .A3(new_n1059), .A4(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT118), .B1(new_n566), .B2(new_n567), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n568), .B(new_n575), .C1(new_n1092), .C2(KEYINPUT57), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n579), .B2(new_n565), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1094), .B(new_n1096), .C1(new_n580), .C2(new_n574), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1061), .A2(new_n818), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1009), .A2(new_n1018), .A3(new_n1019), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1098), .B(new_n1101), .C1(new_n1030), .C2(G1956), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1091), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(KEYINPUT121), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(KEYINPUT61), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1105), .A2(KEYINPUT122), .A3(KEYINPUT61), .A4(new_n1106), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G1348), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1061), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1070), .A2(new_n998), .A3(new_n1018), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT119), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(KEYINPUT119), .B(new_n1114), .C1(new_n1030), .C2(G1348), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT60), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1114), .B1(new_n1030), .B2(G1348), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n1116), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1118), .A2(new_n618), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1126));
  OAI211_X1 g701(.A(KEYINPUT60), .B(new_n607), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT58), .B(G1341), .Z(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1010), .B2(new_n1007), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1020), .B2(G1996), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n557), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT59), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1111), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1121), .A2(new_n618), .A3(new_n1116), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1102), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1104), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1137), .B(KEYINPUT120), .Z(new_n1138));
  AOI21_X1  g713(.A(new_n1090), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1059), .A2(KEYINPUT62), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1055), .A2(new_n1141), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1140), .A2(new_n1037), .A3(new_n1089), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1088), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1074), .A2(new_n1078), .A3(new_n700), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1068), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1144), .A2(new_n1081), .B1(new_n1146), .B2(new_n1071), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1053), .A2(new_n1042), .A3(G286), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1066), .A2(new_n1081), .A3(new_n1088), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(G8), .B1(new_n1087), .B2(new_n1060), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1150), .B1(new_n1152), .B2(new_n1065), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1153), .A2(new_n1088), .A3(new_n1081), .A4(new_n1148), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1143), .A2(new_n1147), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1016), .B1(new_n1139), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1003), .A2(new_n725), .A3(new_n721), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n881), .A2(new_n998), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1013), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT46), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1013), .B2(G1996), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1011), .B1(new_n996), .B2(new_n1000), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1011), .A2(KEYINPUT46), .A3(new_n1001), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT47), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1165), .B(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1011), .A2(new_n738), .A3(new_n736), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT48), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1160), .B(new_n1168), .C1(new_n1012), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1157), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g747(.A1(new_n461), .A2(G227), .ZN(new_n1174));
  INV_X1    g748(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g749(.A(new_n1175), .B1(new_n989), .B2(new_n991), .ZN(new_n1176));
  NOR2_X1   g750(.A1(G401), .A2(G229), .ZN(new_n1177));
  AND3_X1   g751(.A1(new_n1176), .A2(new_n914), .A3(new_n1177), .ZN(G308));
  NAND3_X1  g752(.A1(new_n1176), .A2(new_n914), .A3(new_n1177), .ZN(G225));
endmodule


