//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n465), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(new_n472), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT68), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n473), .A2(G136), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT67), .ZN(new_n488));
  INV_X1    g063(.A(G100), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n489), .A2(new_n464), .A3(KEYINPUT69), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT69), .B1(new_n489), .B2(new_n464), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G112), .B2(new_n464), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n486), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n479), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n462), .A2(new_n464), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n473), .A2(new_n502), .A3(G138), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT72), .B1(new_n505), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT5), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(new_n509), .B1(new_n505), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .A3(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT70), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT70), .A2(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(KEYINPUT6), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n510), .A2(new_n516), .A3(G88), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n516), .A2(G543), .A3(new_n519), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(new_n518), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  OAI221_X1 g100(.A(new_n520), .B1(new_n521), .B2(new_n522), .C1(new_n523), .C2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(G166));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n510), .A2(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n510), .A2(new_n516), .A3(G89), .A4(new_n519), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n516), .A2(G51), .A3(G543), .A4(new_n519), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(G168));
  NAND4_X1  g110(.A1(new_n510), .A2(new_n516), .A3(G90), .A4(new_n519), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT74), .B(G52), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n516), .A2(G543), .A3(new_n519), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n505), .A2(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n507), .B1(KEYINPUT5), .B2(new_n508), .ZN(new_n540));
  NOR3_X1   g115(.A1(new_n505), .A2(KEYINPUT72), .A3(G543), .ZN(new_n541));
  OAI211_X1 g116(.A(G64), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n525), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n536), .B(new_n538), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  NOR3_X1   g122(.A1(new_n547), .A2(KEYINPUT73), .A3(new_n525), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(G171));
  NAND4_X1  g124(.A1(new_n516), .A2(G43), .A3(G543), .A4(new_n519), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n510), .A2(new_n516), .A3(G81), .A4(new_n519), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(new_n525), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(new_n521), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(G53), .A3(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n561), .B(KEYINPUT9), .C1(new_n521), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n516), .A2(new_n519), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT76), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n570), .A2(KEYINPUT76), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n571), .B(new_n572), .C1(new_n568), .C2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(G91), .A2(new_n569), .B1(new_n574), .B2(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n566), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  NAND3_X1  g152(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(G286));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n526), .A2(new_n579), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n523), .A2(new_n525), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n560), .A2(G50), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT77), .A4(new_n520), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(G303));
  NAND4_X1  g159(.A1(new_n510), .A2(new_n516), .A3(G87), .A4(new_n519), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n521), .ZN(G288));
  NAND4_X1  g163(.A1(new_n510), .A2(new_n516), .A3(G86), .A4(new_n519), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n516), .A2(G48), .A3(G543), .A4(new_n519), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n510), .A2(G61), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(new_n524), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT78), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n525), .B1(new_n593), .B2(new_n594), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  NOR3_X1   g174(.A1(new_n591), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(G305));
  NAND4_X1  g176(.A1(new_n510), .A2(new_n516), .A3(G85), .A4(new_n519), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n521), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n510), .A2(G60), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n525), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND4_X1  g184(.A1(new_n510), .A2(new_n516), .A3(G92), .A4(new_n519), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n568), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n560), .A2(G54), .B1(new_n615), .B2(G651), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n618), .B2(G171), .ZN(G284));
  OAI21_X1  g195(.A(new_n619), .B1(new_n618), .B2(G171), .ZN(G321));
  NAND2_X1  g196(.A1(G299), .A2(new_n618), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n618), .B2(G168), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(new_n618), .B2(G168), .ZN(G280));
  INV_X1    g199(.A(new_n617), .ZN(new_n625));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n631));
  XNOR2_X1  g206(.A(G323), .B(new_n631), .ZN(G282));
  NAND2_X1  g207(.A1(new_n485), .A2(G123), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(G135), .B2(new_n473), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT80), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n638), .A2(G2096), .ZN(new_n646));
  NAND4_X1  g221(.A1(new_n639), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(G156));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT82), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2451), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n652), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2454), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2096), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n682), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n683), .A2(KEYINPUT20), .A3(new_n682), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n684), .B1(new_n682), .B2(new_n680), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT84), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  XNOR2_X1  g272(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT91), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G26), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n480), .A2(new_n483), .A3(G128), .ZN(new_n703));
  INV_X1    g278(.A(G104), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(new_n464), .A3(KEYINPUT89), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G104), .B2(G2105), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G116), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n470), .B1(new_n709), .B2(G2105), .ZN(new_n710));
  AOI22_X1  g285(.A1(G140), .A2(new_n473), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n702), .B1(G29), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G2067), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT31), .B(G11), .Z(new_n716));
  NOR2_X1   g291(.A1(new_n638), .A2(new_n700), .ZN(new_n717));
  INV_X1    g292(.A(G28), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n719));
  AOI21_X1  g294(.A(G29), .B1(new_n718), .B2(KEYINPUT30), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n716), .B(new_n717), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NOR2_X1   g297(.A1(G168), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n722), .B2(G21), .ZN(new_n724));
  INV_X1    g299(.A(G1966), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n700), .B1(KEYINPUT24), .B2(G34), .ZN(new_n728));
  OAI22_X1  g303(.A1(G160), .A2(new_n700), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G2084), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(G2084), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n721), .A2(new_n726), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G19), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n554), .B2(G16), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n715), .B(new_n732), .C1(G1341), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(G1341), .ZN(new_n736));
  AND3_X1   g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT26), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n473), .A2(G141), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n480), .A2(new_n483), .A3(G129), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(new_n700), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n700), .B2(G32), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI22_X1  g323(.A1(new_n748), .A2(KEYINPUT92), .B1(new_n725), .B2(new_n724), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n736), .B(new_n749), .C1(KEYINPUT92), .C2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n722), .A2(G20), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT23), .Z(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G299), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1956), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n735), .A2(new_n750), .A3(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n746), .A2(new_n747), .ZN(new_n756));
  NOR2_X1   g331(.A1(G29), .A2(G33), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT25), .Z(new_n759));
  INV_X1    g334(.A(G139), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n499), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n462), .A2(G127), .ZN(new_n762));
  NAND2_X1  g337(.A1(G115), .A2(G2104), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n464), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n757), .B1(new_n765), .B2(G29), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G2072), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n700), .A2(G27), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT94), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n700), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G2078), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(G2078), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n756), .A2(new_n767), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n625), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G4), .B2(G16), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G5), .A2(G16), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT93), .Z(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G301), .B2(new_n722), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1961), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n777), .B(new_n781), .C1(new_n774), .C2(new_n776), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n700), .A2(G35), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G162), .B2(new_n700), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2090), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n755), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n700), .A2(G25), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n485), .A2(G119), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n791));
  INV_X1    g366(.A(G107), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G2105), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G131), .B2(new_n473), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n789), .B1(new_n796), .B2(new_n700), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT35), .B(G1991), .Z(new_n798));
  XOR2_X1   g373(.A(new_n797), .B(new_n798), .Z(new_n799));
  NOR2_X1   g374(.A1(new_n608), .A2(new_n722), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n722), .B2(G24), .ZN(new_n801));
  INV_X1    g376(.A(G1986), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n799), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n722), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n722), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G1971), .Z(new_n808));
  AND2_X1   g383(.A1(new_n722), .A2(G6), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G305), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT32), .B(G1981), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT85), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n810), .A2(new_n812), .ZN(new_n814));
  MUX2_X1   g389(.A(G23), .B(G288), .S(G16), .Z(new_n815));
  XOR2_X1   g390(.A(KEYINPUT33), .B(G1976), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT86), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n808), .A2(new_n813), .A3(new_n814), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n805), .B1(new_n819), .B2(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT87), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT87), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT88), .B(KEYINPUT36), .Z(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n788), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n826), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n827), .A2(new_n829), .ZN(G311));
  OR2_X1    g405(.A1(new_n824), .A2(new_n826), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n831), .A2(new_n828), .A3(new_n788), .ZN(G150));
  XOR2_X1   g407(.A(KEYINPUT97), .B(G860), .Z(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n617), .A2(new_n626), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n552), .A2(new_n525), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n551), .A2(new_n550), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n510), .A2(new_n516), .A3(G93), .A4(new_n519), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n516), .A2(G55), .A3(G543), .A4(new_n519), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n510), .A2(G67), .ZN(new_n843));
  AND2_X1   g418(.A1(G80), .A2(G543), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n524), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n838), .A2(new_n839), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n844), .B1(new_n510), .B2(G67), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n841), .B(new_n840), .C1(new_n847), .C2(new_n525), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n553), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n837), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n834), .B1(new_n852), .B2(KEYINPUT39), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(KEYINPUT39), .B2(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n848), .A2(new_n834), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT37), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  INV_X1    g434(.A(new_n742), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n703), .B(new_n711), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n712), .A2(new_n742), .A3(new_n741), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n501), .A2(new_n503), .ZN(new_n865));
  INV_X1    g440(.A(new_n498), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n862), .A2(new_n863), .A3(G164), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n765), .B1(new_n870), .B2(KEYINPUT98), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n868), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n859), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n862), .A2(new_n863), .A3(G164), .ZN(new_n875));
  AOI21_X1  g450(.A(G164), .B1(new_n862), .B2(new_n863), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT98), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n765), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n877), .A2(new_n873), .A3(new_n859), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n870), .A2(new_n765), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n858), .B1(new_n874), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n873), .A3(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT99), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n884), .A2(KEYINPUT101), .A3(new_n880), .A4(new_n879), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  INV_X1    g461(.A(G118), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n886), .B1(new_n887), .B2(G2105), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n888), .B1(G142), .B2(new_n473), .ZN(new_n889));
  INV_X1    g464(.A(G130), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n484), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT100), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n641), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n795), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n882), .A2(new_n885), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT102), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n882), .A2(new_n897), .A3(new_n885), .A4(new_n894), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n638), .B(G160), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(G162), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n874), .A2(new_n881), .ZN(new_n901));
  INV_X1    g476(.A(new_n894), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n896), .A2(new_n898), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n902), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n894), .B1(new_n874), .B2(new_n881), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G37), .B1(new_n907), .B2(new_n900), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n904), .A2(KEYINPUT40), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT40), .B1(new_n904), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(G395));
  AND2_X1   g486(.A1(new_n846), .A2(new_n849), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n628), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G299), .A2(new_n617), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n566), .A2(new_n612), .A3(new_n575), .A4(new_n616), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR3_X1    g491(.A1(new_n913), .A2(KEYINPUT103), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n913), .A2(new_n916), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n914), .A2(KEYINPUT41), .A3(new_n915), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n914), .B2(new_n915), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT103), .B1(new_n913), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n917), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(KEYINPUT105), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n926));
  OAI221_X1 g501(.A(new_n917), .B1(new_n926), .B2(KEYINPUT42), .C1(new_n918), .C2(new_n922), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n604), .A2(new_n607), .A3(KEYINPUT104), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT104), .B1(new_n604), .B2(new_n607), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n929), .B(new_n930), .C1(new_n597), .C2(new_n600), .ZN(new_n931));
  INV_X1    g506(.A(new_n600), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n599), .B1(new_n591), .B2(new_n598), .ZN(new_n933));
  INV_X1    g508(.A(new_n930), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n932), .B(new_n933), .C1(new_n934), .C2(new_n928), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n526), .B(G288), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n931), .A2(new_n935), .A3(new_n937), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(new_n926), .B2(KEYINPUT42), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n925), .A2(new_n927), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n925), .B2(new_n927), .ZN(new_n944));
  OAI21_X1  g519(.A(G868), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n848), .A2(new_n618), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(G295));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n946), .ZN(G331));
  NAND3_X1  g523(.A1(new_n939), .A2(KEYINPUT108), .A3(new_n940), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n931), .A2(new_n935), .A3(new_n937), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n937), .B1(new_n931), .B2(new_n935), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(G286), .B1(new_n546), .B2(new_n548), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n544), .A2(new_n545), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT73), .B1(new_n547), .B2(new_n525), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n536), .A2(new_n538), .ZN(new_n957));
  NAND4_X1  g532(.A1(G168), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n954), .A2(new_n958), .A3(new_n846), .A4(new_n849), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n912), .A2(KEYINPUT107), .A3(new_n954), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n954), .A2(new_n958), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n963), .A2(new_n964), .A3(new_n850), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n964), .B1(new_n963), .B2(new_n850), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n961), .B(new_n962), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(new_n916), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n850), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n959), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n921), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n949), .B(new_n953), .C1(new_n968), .C2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(new_n916), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n967), .B2(new_n921), .ZN(new_n974));
  AOI21_X1  g549(.A(G37), .B1(new_n974), .B2(new_n941), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT110), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(KEYINPUT43), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n965), .A2(new_n966), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n962), .A2(new_n961), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n921), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n973), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n941), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G37), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n953), .A2(new_n949), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(new_n974), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n981), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n980), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT43), .B1(new_n988), .B2(new_n990), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n972), .A2(new_n975), .A3(new_n992), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n995), .B1(new_n998), .B2(new_n981), .ZN(new_n999));
  AOI211_X1 g574(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n996), .C2(new_n997), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n994), .B1(new_n999), .B2(new_n1000), .ZN(G397));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(G164), .B2(G1384), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G160), .A2(G40), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n743), .B(G1996), .Z(new_n1006));
  XNOR2_X1  g581(.A(new_n712), .B(new_n714), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(new_n795), .B(new_n798), .Z(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n802), .B2(new_n608), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n608), .A2(new_n802), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT111), .Z(new_n1013));
  OAI21_X1  g588(.A(new_n1005), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n865), .B2(new_n866), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT113), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1019), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1004), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1961), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n867), .A2(KEYINPUT45), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1003), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1016), .A2(KEYINPUT112), .A3(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G2078), .ZN(new_n1030));
  INV_X1    g605(.A(G40), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n465), .A2(new_n475), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1023), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1025), .A2(new_n1003), .A3(new_n1032), .ZN(new_n1036));
  OR3_X1    g611(.A1(new_n1036), .A2(KEYINPUT125), .A3(G2078), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT125), .B1(new_n1036), .B2(G2078), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(KEYINPUT53), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(G301), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1004), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT53), .B1(new_n1041), .B2(new_n1030), .ZN(new_n1042));
  INV_X1    g617(.A(new_n463), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n464), .B1(new_n1043), .B2(KEYINPUT126), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(KEYINPUT126), .B2(new_n1043), .ZN(new_n1045));
  NOR4_X1   g620(.A1(new_n475), .A2(new_n1034), .A3(new_n1031), .A4(G2078), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1048));
  NOR4_X1   g623(.A1(new_n1042), .A2(G171), .A3(new_n1023), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1015), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  INV_X1    g626(.A(G2084), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1021), .A2(new_n1052), .A3(new_n1022), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1036), .A2(new_n725), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G286), .A2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1055), .A2(KEYINPUT51), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G8), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1056), .B(KEYINPUT124), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g638(.A(new_n1051), .B(G168), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1058), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1035), .A2(G301), .A3(new_n1039), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1042), .A2(new_n1023), .A3(new_n1048), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1067), .B(KEYINPUT54), .C1(G301), .C2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n580), .A2(new_n583), .A3(G8), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(KEYINPUT55), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n580), .A2(new_n583), .A3(G8), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1971), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1079));
  INV_X1    g654(.A(G2090), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1021), .A2(new_n1080), .A3(new_n1022), .ZN(new_n1081));
  OAI211_X1 g656(.A(G8), .B(new_n1078), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1016), .A2(new_n1032), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(G1976), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G288), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT52), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1051), .B1(new_n1016), .B2(new_n1032), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT52), .B1(G288), .B2(new_n1085), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1088), .B(new_n1089), .C1(new_n1085), .C2(G288), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  OR3_X1    g666(.A1(new_n591), .A2(new_n598), .A3(G1981), .ZN(new_n1092));
  OAI21_X1  g667(.A(G1981), .B1(new_n591), .B2(new_n598), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT49), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT115), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1092), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1091), .B1(new_n1088), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1082), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n867), .A2(new_n1024), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT50), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1022), .A2(new_n1102), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1041), .A2(G1971), .B1(new_n1103), .B2(G2090), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1078), .B1(new_n1104), .B2(G8), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1050), .A2(new_n1066), .A3(new_n1069), .A4(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1041), .A2(new_n1108), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n575), .B2(KEYINPUT118), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(G299), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n566), .B(new_n575), .C1(KEYINPUT118), .C2(KEYINPUT57), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1116));
  NOR4_X1   g691(.A1(new_n1110), .A2(new_n1115), .A3(KEYINPUT120), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1041), .A2(new_n1108), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1118), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(G1348), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1083), .A2(G2067), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI22_X1  g701(.A1(new_n1117), .A2(new_n1123), .B1(new_n617), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1110), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1120), .A2(KEYINPUT123), .A3(new_n1128), .A4(new_n1121), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1131), .A2(KEYINPUT61), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1132), .B(new_n1134), .C1(new_n1117), .C2(new_n1123), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1126), .A2(KEYINPUT60), .A3(new_n617), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1125), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1032), .B1(new_n1101), .B2(KEYINPUT50), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT60), .B(new_n1137), .C1(new_n1139), .C2(G1348), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1142), .A3(new_n625), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT121), .B(G1996), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1041), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT58), .B(G1341), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1016), .B2(new_n1032), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n554), .B(new_n1144), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1148), .B1(new_n1041), .B2(new_n1145), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n553), .ZN(new_n1152));
  AND4_X1   g727(.A1(new_n1136), .A2(new_n1143), .A3(new_n1149), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1129), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1110), .A2(new_n1128), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1135), .A2(new_n1153), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1107), .B1(new_n1130), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(G171), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1161), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1061), .A2(new_n1059), .A3(new_n1056), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1062), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT51), .B1(new_n1055), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1163), .B1(new_n1165), .B2(new_n1064), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1163), .B(KEYINPUT62), .C1(new_n1165), .C2(new_n1064), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1162), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(G8), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1171), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1055), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n1082), .A4(new_n1099), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1055), .A2(G168), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1100), .A2(new_n1105), .A3(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1174), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1082), .ZN(new_n1179));
  NOR2_X1   g754(.A1(G288), .A2(G1976), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT116), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1092), .B1(new_n1098), .B2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1179), .A2(new_n1099), .B1(new_n1088), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1170), .A2(new_n1178), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1014), .B1(new_n1159), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1013), .A2(KEYINPUT48), .A3(new_n1005), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1005), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1186), .B1(new_n1187), .B2(new_n1010), .ZN(new_n1188));
  AOI21_X1  g763(.A(KEYINPUT48), .B1(new_n1013), .B2(new_n1005), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OR3_X1    g765(.A1(new_n1187), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1191));
  OAI21_X1  g766(.A(KEYINPUT46), .B1(new_n1187), .B2(G1996), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1007), .A2(new_n744), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1191), .A2(new_n1192), .B1(new_n1005), .B2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT47), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n796), .A2(new_n798), .ZN(new_n1196));
  OAI22_X1  g771(.A1(new_n1008), .A2(new_n1196), .B1(G2067), .B2(new_n712), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1190), .B(new_n1195), .C1(new_n1005), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1185), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g774(.A1(new_n904), .A2(new_n908), .ZN(new_n1201));
  INV_X1    g775(.A(new_n1201), .ZN(new_n1202));
  NOR3_X1   g776(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1203));
  NAND3_X1  g777(.A1(new_n998), .A2(new_n696), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g778(.A1(new_n1202), .A2(new_n1204), .ZN(G308));
  NAND4_X1  g779(.A1(new_n1201), .A2(new_n696), .A3(new_n998), .A4(new_n1203), .ZN(G225));
endmodule


