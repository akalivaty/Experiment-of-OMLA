//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1154, new_n1155, new_n1156, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND3_X1  g0013(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n206), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n213), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(new_n210), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n218), .B(new_n226), .C1(KEYINPUT1), .C2(new_n224), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G68), .Z(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  OAI21_X1  g0044(.A(G20), .B1(new_n207), .B2(G50), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT8), .B(G58), .Z(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(G20), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n246), .A2(new_n248), .B1(G150), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT69), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  NAND4_X1  g0055(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT70), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n255), .A4(new_n256), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G20), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G13), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n251), .A2(new_n261), .B1(new_n215), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n263), .B(KEYINPUT71), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n259), .A2(new_n267), .A3(new_n264), .A4(new_n260), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n266), .B1(new_n215), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G1), .A3(G13), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT68), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G222), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(G1698), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n279), .B1(new_n280), .B2(new_n275), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n277), .A2(new_n274), .A3(new_n278), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n273), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n272), .A2(new_n287), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(G226), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G179), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n270), .B(new_n293), .C1(new_n294), .C2(new_n292), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(G200), .B2(new_n292), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n270), .A2(KEYINPUT9), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n270), .A2(KEYINPUT9), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n298), .A2(new_n303), .A3(new_n299), .A4(new_n300), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n295), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT77), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G33), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n307), .A2(new_n309), .A3(G226), .A4(G1698), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n307), .A2(new_n309), .A3(G223), .A4(new_n276), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G87), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n313), .A2(new_n273), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n272), .A2(G232), .A3(new_n287), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT76), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n289), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n272), .A2(new_n287), .A3(KEYINPUT76), .A4(G232), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n314), .A2(new_n320), .A3(G190), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n313), .A2(new_n273), .ZN(new_n323));
  AOI21_X1  g0123(.A(G200), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n306), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT16), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G20), .ZN(new_n328));
  INV_X1    g0128(.A(G159), .ZN(new_n329));
  INV_X1    g0129(.A(new_n249), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n275), .B2(G20), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n307), .A2(new_n309), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT7), .A3(new_n262), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n202), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n326), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n275), .A2(new_n332), .A3(G20), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT7), .B1(new_n334), .B2(new_n262), .ZN(new_n339));
  OAI21_X1  g0139(.A(G68), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n327), .A2(G20), .B1(G159), .B2(new_n249), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(KEYINPUT16), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n337), .A2(new_n342), .A3(new_n261), .ZN(new_n343));
  MUX2_X1   g0143(.A(new_n264), .B(new_n268), .S(new_n246), .Z(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n314), .B2(new_n320), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n322), .A2(new_n296), .A3(new_n323), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT77), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n325), .A2(new_n343), .A3(new_n344), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT17), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n343), .A2(new_n344), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT17), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(new_n325), .A4(new_n348), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n343), .A2(new_n344), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n314), .A2(G179), .A3(new_n320), .ZN(new_n355));
  AOI21_X1  g0155(.A(G169), .B1(new_n322), .B2(new_n323), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT18), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n357), .A3(KEYINPUT18), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n350), .A2(new_n353), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT15), .B(G87), .Z(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n248), .ZN(new_n364));
  INV_X1    g0164(.A(new_n246), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n364), .B1(new_n262), .B2(new_n280), .C1(new_n365), .C2(new_n330), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n261), .B1(new_n280), .B2(new_n265), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n280), .B2(new_n268), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n290), .A2(G244), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n275), .A2(G232), .A3(new_n276), .ZN(new_n371));
  INV_X1    g0171(.A(G107), .ZN(new_n372));
  INV_X1    g0172(.A(G238), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n371), .B1(new_n372), .B2(new_n275), .C1(new_n282), .C2(new_n373), .ZN(new_n374));
  AOI211_X1 g0174(.A(new_n289), .B(new_n370), .C1(new_n374), .C2(new_n273), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G190), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n369), .B(new_n376), .C1(new_n345), .C2(new_n375), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n375), .A2(G169), .ZN(new_n378));
  INV_X1    g0178(.A(G179), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n368), .A3(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n305), .A2(new_n362), .A3(new_n377), .A4(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n289), .B1(new_n290), .B2(G238), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n307), .A2(new_n309), .A3(G232), .A4(G1698), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n307), .A2(new_n309), .A3(G226), .A4(new_n276), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G97), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT72), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n387), .A2(new_n388), .A3(new_n273), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n388), .B1(new_n387), .B2(new_n273), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n383), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT13), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n393), .B(new_n383), .C1(new_n389), .C2(new_n390), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(KEYINPUT73), .A3(new_n394), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n389), .A2(new_n390), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT73), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(new_n393), .A4(new_n383), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n294), .B1(KEYINPUT75), .B2(KEYINPUT14), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n395), .A2(new_n401), .A3(new_n398), .A4(new_n399), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n392), .A2(G179), .A3(new_n394), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n248), .A2(G77), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n262), .B2(G68), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(KEYINPUT74), .B1(G50), .B2(new_n249), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(KEYINPUT74), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n261), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT11), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n268), .A2(new_n202), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n265), .A2(new_n202), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT12), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n410), .A2(KEYINPUT11), .A3(new_n261), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n413), .A2(new_n415), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n406), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n419), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n395), .A2(G200), .A3(new_n398), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n392), .A2(G190), .A3(new_n394), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G283), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n307), .A2(new_n309), .A3(G250), .A4(G1698), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n307), .A2(new_n309), .A3(G244), .A4(new_n276), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT4), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n426), .B(new_n427), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT78), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n275), .A2(KEYINPUT78), .A3(G244), .A4(new_n276), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n429), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n434), .B2(KEYINPUT79), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT79), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n432), .A2(new_n433), .A3(new_n436), .A4(new_n429), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n272), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT5), .B(G41), .ZN(new_n439));
  INV_X1    g0239(.A(G45), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G1), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(G274), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n273), .B1(new_n439), .B2(new_n441), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(G257), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G190), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n286), .A2(G33), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n259), .A2(new_n264), .A3(new_n260), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G97), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT6), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n453), .A2(new_n451), .A3(G107), .ZN(new_n454));
  XNOR2_X1  g0254(.A(G97), .B(G107), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n456), .A2(new_n262), .B1(new_n280), .B2(new_n330), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n372), .B1(new_n333), .B2(new_n335), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n261), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n265), .A2(new_n451), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n452), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n434), .A2(KEYINPUT79), .ZN(new_n462));
  INV_X1    g0262(.A(new_n430), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n462), .A2(new_n437), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n445), .B1(new_n464), .B2(new_n272), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n461), .B1(new_n465), .B2(G200), .ZN(new_n466));
  OAI211_X1 g0266(.A(G179), .B(new_n445), .C1(new_n464), .C2(new_n272), .ZN(new_n467));
  OAI21_X1  g0267(.A(G169), .B1(new_n438), .B2(new_n446), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT80), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n452), .A2(new_n459), .A3(new_n471), .A4(new_n460), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n448), .A2(new_n466), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n275), .A2(G257), .A3(new_n276), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n275), .A2(G264), .A3(G1698), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n334), .A2(G303), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(new_n273), .B1(new_n444), .B2(G270), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n442), .ZN(new_n480));
  INV_X1    g0280(.A(G116), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n450), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n265), .A2(new_n481), .ZN(new_n483));
  AOI21_X1  g0283(.A(G20), .B1(G33), .B2(G283), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n247), .A2(G97), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n484), .A2(new_n485), .B1(G20), .B2(new_n481), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n257), .A2(KEYINPUT20), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT20), .B1(new_n257), .B2(new_n486), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n480), .B(G169), .C1(new_n482), .C2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT21), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n480), .A2(new_n379), .ZN(new_n492));
  OR2_X1    g0292(.A1(new_n482), .A2(new_n489), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n493), .A2(KEYINPUT21), .A3(G169), .A4(new_n480), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n480), .A2(G200), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n482), .A2(new_n489), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n496), .B(new_n497), .C1(new_n296), .C2(new_n480), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n275), .A2(G238), .A3(new_n276), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n275), .A2(G244), .A3(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G116), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n273), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n272), .B(G250), .C1(G1), .C2(new_n440), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n441), .A2(G274), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G200), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n275), .A2(new_n262), .A3(G68), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT81), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n275), .A2(KEYINPUT81), .A3(new_n262), .A4(G68), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n248), .A2(new_n515), .A3(G97), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  INV_X1    g0317(.A(G87), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n517), .A2(new_n518), .B1(new_n386), .B2(new_n262), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n516), .B1(new_n519), .B2(new_n515), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n513), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n363), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n521), .A2(new_n261), .B1(new_n265), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g0323(.A1(new_n450), .A2(new_n518), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n507), .B1(new_n503), .B2(new_n273), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G190), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n510), .A2(new_n523), .A3(new_n524), .A4(new_n526), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n450), .A2(new_n522), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n523), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(new_n379), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(G169), .B2(new_n525), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n527), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n450), .A2(new_n372), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n265), .A2(new_n372), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n535), .B(KEYINPUT25), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n307), .A2(new_n309), .A3(new_n262), .A4(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n275), .A2(new_n541), .A3(new_n262), .A4(G87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT24), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n502), .A2(G20), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT82), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n262), .B2(G107), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT23), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT23), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n546), .B(new_n549), .C1(new_n262), .C2(G107), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n545), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n543), .A2(new_n544), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n544), .B1(new_n543), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n261), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT83), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(KEYINPUT83), .B(new_n261), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n538), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G257), .ZN(new_n559));
  INV_X1    g0359(.A(G294), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n282), .A2(new_n559), .B1(new_n247), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G250), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n277), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n273), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n443), .B1(new_n444), .B2(G264), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(new_n296), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n345), .B1(new_n564), .B2(new_n565), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n533), .B1(new_n558), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n566), .A2(new_n294), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G179), .B2(new_n566), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n558), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n474), .A2(new_n499), .A3(new_n570), .A4(new_n573), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n382), .A2(new_n425), .A3(new_n574), .ZN(G372));
  NOR2_X1   g0375(.A1(new_n382), .A2(new_n425), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n494), .B(new_n495), .C1(new_n558), .C2(new_n572), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n474), .A2(new_n570), .A3(new_n577), .ZN(new_n578));
  AOI211_X1 g0378(.A(G179), .B(new_n507), .C1(new_n503), .C2(new_n273), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n294), .B2(new_n509), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n529), .ZN(new_n581));
  INV_X1    g0381(.A(new_n461), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n467), .B2(new_n468), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n510), .A2(new_n526), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n524), .A2(new_n523), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n584), .A2(new_n585), .B1(new_n580), .B2(new_n529), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT26), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n469), .A2(new_n473), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT26), .B1(new_n589), .B2(new_n533), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n578), .A2(new_n581), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n576), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g0392(.A(new_n592), .B(KEYINPUT84), .Z(new_n593));
  NAND2_X1  g0393(.A1(new_n360), .A2(new_n361), .ZN(new_n594));
  INV_X1    g0394(.A(new_n381), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n406), .B2(new_n419), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n350), .A2(new_n353), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n424), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n302), .A2(new_n304), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n295), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n593), .A2(new_n601), .ZN(G369));
  NAND2_X1  g0402(.A1(new_n494), .A2(new_n495), .ZN(new_n603));
  INV_X1    g0403(.A(G13), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(G20), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n286), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT85), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT27), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(G213), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(G343), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(new_n497), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n603), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n616), .B1(new_n617), .B2(new_n615), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(G330), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n556), .A2(new_n557), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(new_n537), .A3(new_n569), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n558), .B2(new_n614), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n573), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n558), .A2(new_n572), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n614), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n613), .B1(new_n494), .B2(new_n495), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n623), .A2(new_n628), .B1(new_n624), .B2(new_n614), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(G399));
  INV_X1    g0430(.A(new_n211), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(G41), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NOR4_X1   g0433(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G1), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n217), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT28), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT86), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n574), .B2(new_n613), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT30), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n479), .A2(new_n525), .A3(new_n564), .A4(new_n565), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n467), .B2(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n479), .A2(new_n525), .A3(new_n564), .A4(new_n565), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n447), .A2(KEYINPUT30), .A3(G179), .A4(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n566), .A2(new_n379), .A3(new_n509), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n465), .A2(new_n480), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n642), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n647), .A2(KEYINPUT31), .A3(new_n613), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT31), .B1(new_n647), .B2(new_n613), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n621), .A2(new_n586), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n651), .A2(new_n617), .A3(new_n624), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n652), .A2(KEYINPUT86), .A3(new_n474), .A4(new_n614), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n639), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(G330), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n586), .A2(new_n469), .A3(new_n587), .A4(new_n473), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n583), .A2(new_n586), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT26), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n578), .A2(new_n581), .A3(new_n656), .A4(new_n658), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n659), .A2(KEYINPUT29), .A3(new_n614), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT29), .B1(new_n591), .B2(new_n614), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT87), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(KEYINPUT29), .A3(new_n614), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT87), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n655), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n637), .B1(new_n666), .B2(G1), .ZN(G364));
  AOI21_X1  g0467(.A(new_n286), .B1(new_n605), .B2(G45), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n633), .A2(KEYINPUT88), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT88), .ZN(new_n670));
  INV_X1    g0470(.A(new_n668), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n632), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(G355), .A2(KEYINPUT89), .ZN(new_n674));
  NAND2_X1  g0474(.A1(G355), .A2(KEYINPUT89), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n674), .A2(new_n211), .A3(new_n275), .A4(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n243), .A2(new_n440), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n631), .A2(new_n275), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n217), .B2(G45), .ZN(new_n679));
  OAI221_X1 g0479(.A(new_n676), .B1(G116), .B2(new_n211), .C1(new_n677), .C2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(G13), .A2(G33), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G20), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n255), .B1(G20), .B2(new_n294), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n673), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n262), .A2(new_n296), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n379), .A3(G200), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n262), .A2(G190), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n379), .A2(G200), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n689), .A2(G87), .B1(new_n693), .B2(G77), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n379), .A2(new_n345), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n690), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n694), .B1(new_n202), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n687), .ZN(new_n698));
  INV_X1    g0498(.A(new_n690), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n699), .A2(G179), .A3(new_n345), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI221_X1 g0501(.A(new_n275), .B1(new_n215), .B2(new_n698), .C1(new_n701), .C2(new_n372), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT91), .ZN(new_n703));
  OAI21_X1  g0503(.A(G20), .B1(G179), .B2(G200), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n699), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n703), .B1(new_n699), .B2(new_n704), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI211_X1 g0508(.A(new_n697), .B(new_n702), .C1(new_n708), .C2(G97), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n687), .A2(new_n691), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n699), .A2(G179), .A3(G200), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G159), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n711), .A2(new_n201), .B1(new_n713), .B2(KEYINPUT32), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(KEYINPUT32), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n708), .A2(G294), .ZN(new_n716));
  INV_X1    g0516(.A(new_n710), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n275), .B1(new_n717), .B2(G322), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(G329), .ZN(new_n719));
  INV_X1    g0519(.A(G283), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n718), .B(new_n719), .C1(new_n701), .C2(new_n720), .ZN(new_n721));
  XOR2_X1   g0521(.A(KEYINPUT33), .B(G317), .Z(new_n722));
  INV_X1    g0522(.A(G311), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n722), .A2(new_n696), .B1(new_n692), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G303), .ZN(new_n725));
  INV_X1    g0525(.A(G326), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n688), .A2(new_n725), .B1(new_n698), .B2(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n721), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n709), .A2(new_n715), .B1(new_n716), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n684), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n686), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT92), .Z(new_n732));
  INV_X1    g0532(.A(new_n683), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n732), .B1(new_n618), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n619), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n673), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n618), .A2(G330), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(G396));
  NAND2_X1  g0538(.A1(new_n591), .A2(new_n614), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n377), .B1(new_n369), .B2(new_n614), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n381), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n595), .A2(new_n614), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n739), .B(new_n743), .Z(new_n744));
  INV_X1    g0544(.A(new_n655), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n673), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n744), .B2(new_n745), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n684), .A2(new_n681), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n747), .B1(G77), .B2(new_n751), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n688), .A2(new_n372), .B1(new_n710), .B2(new_n560), .ZN(new_n753));
  INV_X1    g0553(.A(new_n698), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n275), .B(new_n753), .C1(G303), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n708), .A2(G97), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G87), .A2(new_n700), .B1(new_n712), .B2(G311), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n696), .A2(new_n720), .B1(new_n692), .B2(new_n481), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT93), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n755), .A2(new_n756), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT94), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n701), .A2(new_n202), .ZN(new_n762));
  INV_X1    g0562(.A(new_n712), .ZN(new_n763));
  INV_X1    g0563(.A(G132), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n275), .B1(new_n215), .B2(new_n688), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n762), .B(new_n765), .C1(new_n708), .C2(G58), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n754), .A2(G137), .B1(new_n693), .B2(G159), .ZN(new_n769));
  INV_X1    g0569(.A(G150), .ZN(new_n770));
  INV_X1    g0570(.A(G143), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n769), .B1(new_n770), .B2(new_n696), .C1(new_n711), .C2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT34), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT95), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n766), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n761), .B1(new_n768), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n752), .B1(new_n776), .B2(new_n684), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n743), .B2(new_n682), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT96), .Z(new_n779));
  NOR2_X1   g0579(.A1(new_n749), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(G384));
  OAI21_X1  g0581(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n217), .A2(new_n782), .B1(G50), .B2(new_n202), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(G1), .A3(new_n604), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT35), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n481), .B(new_n214), .C1(new_n456), .C2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n785), .B2(new_n456), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n788));
  OAI21_X1  g0588(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n787), .B2(new_n788), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT39), .ZN(new_n791));
  INV_X1    g0591(.A(new_n611), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n354), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n349), .A2(new_n358), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT37), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n349), .A2(new_n358), .A3(new_n793), .A4(KEYINPUT37), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(new_n362), .C2(new_n793), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(KEYINPUT100), .A3(KEYINPUT38), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(KEYINPUT38), .B1(new_n798), .B2(KEYINPUT100), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n791), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT38), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n597), .A2(new_n594), .ZN(new_n804));
  INV_X1    g0604(.A(new_n793), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n796), .A2(new_n797), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n793), .B1(new_n597), .B2(new_n594), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n796), .A2(new_n797), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n809), .A2(new_n810), .A3(KEYINPUT38), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n802), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n406), .A2(new_n419), .A3(new_n614), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT99), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n591), .A2(new_n614), .A3(new_n743), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n421), .A2(new_n614), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT98), .B1(new_n406), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n406), .A2(KEYINPUT98), .A3(new_n822), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n822), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n420), .A2(new_n424), .A3(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n821), .A2(new_n742), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n812), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n360), .A2(new_n361), .A3(new_n611), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n820), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n662), .A2(new_n576), .A3(new_n665), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n833), .A2(new_n601), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n832), .B(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n801), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n836), .A2(KEYINPUT40), .A3(new_n799), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n406), .A2(KEYINPUT98), .A3(new_n822), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n828), .B1(new_n823), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n654), .A2(new_n839), .A3(new_n743), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n812), .A2(new_n654), .A3(new_n839), .A4(new_n743), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT40), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n843), .A2(KEYINPUT101), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT101), .B1(new_n843), .B2(new_n844), .ZN(new_n846));
  OAI211_X1 g0646(.A(G330), .B(new_n842), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n576), .A2(new_n655), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n843), .A2(new_n844), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT101), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n843), .A2(KEYINPUT101), .A3(new_n844), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n841), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n576), .A2(new_n654), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n847), .A2(new_n848), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n835), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n835), .A2(new_n855), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT102), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n856), .B1(new_n286), .B2(new_n605), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n857), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(KEYINPUT102), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n790), .B1(new_n859), .B2(new_n861), .ZN(G367));
  INV_X1    g0662(.A(new_n678), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n234), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n685), .B1(new_n211), .B2(new_n522), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n747), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT107), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n698), .A2(new_n723), .B1(new_n692), .B2(new_n720), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n689), .A2(G116), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT46), .Z(new_n870));
  INV_X1    g0670(.A(new_n696), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n868), .B(new_n870), .C1(G294), .C2(new_n871), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n872), .B1(new_n372), .B2(new_n707), .C1(new_n725), .C2(new_n711), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n700), .A2(G97), .ZN(new_n874));
  INV_X1    g0674(.A(G317), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n874), .B(new_n334), .C1(new_n763), .C2(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT108), .Z(new_n877));
  NOR2_X1   g0677(.A1(new_n707), .A2(new_n202), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n275), .B1(new_n710), .B2(new_n770), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(G137), .B2(new_n712), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n754), .A2(G143), .B1(new_n693), .B2(G50), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n689), .A2(G58), .B1(new_n871), .B2(G159), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n700), .A2(G77), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n873), .A2(new_n877), .B1(new_n878), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT47), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n730), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n867), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n614), .A2(new_n585), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n890), .A2(new_n581), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n890), .A2(new_n586), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(KEYINPUT103), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(KEYINPUT103), .B2(new_n891), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n889), .B1(new_n894), .B2(new_n733), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n626), .A2(new_n628), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n474), .A2(new_n577), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n896), .A2(KEYINPUT42), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n474), .B1(new_n582), .B2(new_n614), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n583), .A2(new_n613), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n589), .B1(new_n901), .B2(new_n573), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n614), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT42), .B1(new_n896), .B2(new_n897), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n898), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n894), .B(KEYINPUT43), .Z(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT104), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n898), .A2(new_n903), .A3(new_n904), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n894), .A2(KEYINPUT43), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n907), .A2(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n905), .A2(KEYINPUT104), .A3(new_n906), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n627), .A2(new_n901), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT105), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT105), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n911), .A2(new_n917), .A3(new_n914), .A4(new_n912), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n913), .A2(new_n915), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n899), .A2(new_n900), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n629), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT45), .Z(new_n924));
  NOR2_X1   g0724(.A1(new_n629), .A2(new_n922), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT44), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n627), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n927), .B(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n627), .B(KEYINPUT106), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n626), .B(new_n628), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n930), .B1(new_n735), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n666), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n666), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n632), .B(KEYINPUT41), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n671), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n895), .B1(new_n921), .B2(new_n936), .ZN(G387));
  NAND2_X1  g0737(.A1(new_n932), .A2(new_n671), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n626), .A2(new_n733), .ZN(new_n939));
  INV_X1    g0739(.A(new_n685), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n863), .B1(new_n231), .B2(G45), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n246), .A2(new_n943), .A3(new_n215), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n944), .B(new_n440), .C1(new_n202), .C2(new_n280), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n943), .B1(new_n246), .B2(new_n215), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n634), .B1(new_n942), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n942), .B1(new_n631), .B2(new_n334), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n948), .A2(new_n949), .B1(new_n372), .B2(new_n631), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n712), .A2(G150), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n689), .A2(G77), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n874), .A2(new_n951), .A3(new_n275), .A4(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n707), .A2(new_n522), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n365), .A2(new_n696), .B1(new_n202), .B2(new_n692), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n698), .A2(new_n329), .B1(new_n710), .B2(new_n215), .ZN(new_n956));
  NOR4_X1   g0756(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT110), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n711), .A2(new_n875), .B1(new_n725), .B2(new_n692), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT111), .ZN(new_n960));
  AOI22_X1  g0760(.A1(G322), .A2(new_n754), .B1(new_n871), .B2(G311), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT48), .Z(new_n963));
  OAI22_X1  g0763(.A1(new_n707), .A2(new_n720), .B1(new_n560), .B2(new_n688), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n334), .B1(new_n701), .B2(new_n481), .C1(new_n726), .C2(new_n763), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n965), .B2(new_n966), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n958), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n747), .B1(new_n940), .B2(new_n950), .C1(new_n970), .C2(new_n730), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n632), .B(KEYINPUT113), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n933), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n932), .A2(new_n666), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n938), .B1(new_n939), .B2(new_n971), .C1(new_n974), .C2(new_n975), .ZN(G393));
  OAI22_X1  g0776(.A1(new_n696), .A2(new_n725), .B1(new_n692), .B2(new_n560), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n708), .B2(G116), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT115), .Z(new_n979));
  OAI22_X1  g0779(.A1(new_n698), .A2(new_n875), .B1(new_n710), .B2(new_n723), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT52), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n334), .B1(new_n720), .B2(new_n688), .C1(new_n701), .C2(new_n372), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G322), .B2(new_n712), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n979), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n707), .A2(new_n280), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n365), .A2(new_n692), .B1(new_n215), .B2(new_n696), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT114), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n275), .B1(new_n202), .B2(new_n688), .C1(new_n701), .C2(new_n518), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G143), .B2(new_n712), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n698), .A2(new_n770), .B1(new_n710), .B2(new_n329), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT51), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n730), .B1(new_n984), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n239), .A2(new_n678), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n940), .B1(G97), .B2(new_n631), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n673), .B(new_n994), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n922), .B2(new_n733), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n929), .A2(new_n933), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n973), .B1(new_n929), .B2(new_n933), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n998), .B1(new_n668), .B2(new_n929), .C1(new_n999), .C2(new_n1000), .ZN(G390));
  NAND2_X1  g0801(.A1(new_n821), .A2(new_n742), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n819), .B1(new_n1002), .B2(new_n839), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n659), .A2(new_n614), .A3(new_n741), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n742), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n1005), .A2(new_n839), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n836), .A2(new_n817), .A3(new_n818), .A4(new_n799), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n814), .A2(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n654), .A2(new_n839), .A3(G330), .A4(new_n743), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n833), .A2(new_n601), .A3(new_n848), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n654), .A2(G330), .A3(new_n743), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n839), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1005), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n1009), .A3(new_n1016), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n839), .A2(new_n743), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n655), .A2(new_n1018), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1002), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NOR3_X1   g0821(.A1(new_n819), .A2(new_n800), .A3(new_n801), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n802), .B(new_n813), .C1(new_n829), .C2(new_n819), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n1024), .A3(new_n1009), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1011), .A2(new_n1012), .A3(new_n1021), .A4(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1026), .A2(new_n973), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1011), .A2(new_n1025), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1028), .A2(new_n668), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n814), .A2(new_n682), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n762), .B1(G294), .B2(new_n712), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT118), .Z(new_n1036));
  OAI21_X1  g0836(.A(new_n334), .B1(new_n688), .B2(new_n518), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n871), .A2(G107), .B1(new_n693), .B2(G97), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n720), .B2(new_n698), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n985), .B1(G116), .B2(new_n717), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT119), .ZN(new_n1042));
  XOR2_X1   g0842(.A(KEYINPUT54), .B(G143), .Z(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(G137), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n1044), .A2(new_n692), .B1(new_n1045), .B2(new_n696), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n708), .B2(G159), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT116), .Z(new_n1048));
  NOR2_X1   g0848(.A1(new_n688), .A2(new_n770), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT53), .ZN(new_n1050));
  INV_X1    g0850(.A(G128), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n698), .A2(new_n1051), .B1(new_n710), .B2(new_n764), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G125), .B2(new_n712), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n275), .B1(new_n701), .B2(new_n215), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1050), .B(new_n1053), .C1(KEYINPUT117), .C2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(KEYINPUT117), .B2(new_n1054), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1040), .A2(new_n1042), .B1(new_n1048), .B2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n747), .B1(new_n246), .B2(new_n751), .C1(new_n1057), .C2(new_n730), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1034), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1033), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(KEYINPUT120), .ZN(new_n1062));
  OR3_X1    g0862(.A1(new_n1033), .A2(KEYINPUT120), .A3(new_n1059), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1032), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(G378));
  NOR2_X1   g0865(.A1(new_n270), .A2(new_n611), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n305), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n305), .A2(new_n1067), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OR3_X1    g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1071), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n853), .B2(G330), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1074), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n847), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n832), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n847), .A2(new_n1076), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n851), .A2(new_n852), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1080), .A2(G330), .A3(new_n842), .A4(new_n1074), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n832), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1078), .A2(KEYINPUT123), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1026), .A2(new_n1012), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT123), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT57), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n1026), .B2(new_n1012), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1082), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n973), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1084), .A2(new_n671), .A3(new_n1088), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1076), .A2(new_n681), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n747), .B1(G50), .B2(new_n751), .ZN(new_n1100));
  INV_X1    g0900(.A(G41), .ZN(new_n1101));
  AOI21_X1  g0901(.A(G50), .B1(new_n247), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n275), .B2(G41), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n689), .A2(G77), .B1(new_n754), .B2(G116), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n201), .B2(new_n701), .C1(new_n720), .C2(new_n763), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1101), .B(new_n334), .C1(new_n696), .C2(new_n451), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n522), .A2(new_n692), .B1(new_n372), .B2(new_n710), .ZN(new_n1107));
  OR4_X1    g0907(.A1(new_n878), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT58), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1103), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n1109), .B2(new_n1108), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n710), .A2(new_n1051), .B1(new_n692), .B2(new_n1045), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G125), .B2(new_n754), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n689), .A2(new_n1043), .B1(new_n871), .B2(G132), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(new_n770), .C2(new_n707), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT122), .Z(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n247), .B(new_n1101), .C1(new_n701), .C2(new_n329), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G124), .B2(new_n712), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1111), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1100), .B1(new_n1123), .B2(new_n684), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1099), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1098), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1097), .A2(new_n1127), .ZN(G375));
  OR2_X1    g0928(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n935), .A3(new_n1029), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n334), .B1(new_n693), .B2(G150), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n701), .B2(new_n201), .C1(new_n1051), .C2(new_n763), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n689), .A2(G159), .B1(new_n754), .B2(G132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n696), .B2(new_n1044), .C1(new_n711), .C2(new_n1045), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(G50), .C2(new_n708), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n275), .B1(new_n754), .B2(G294), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1136), .B(new_n883), .C1(new_n725), .C2(new_n763), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n688), .A2(new_n451), .B1(new_n692), .B2(new_n372), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n481), .A2(new_n696), .B1(new_n710), .B2(new_n720), .ZN(new_n1139));
  NOR4_X1   g0939(.A1(new_n1137), .A2(new_n954), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n684), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1141), .B(new_n747), .C1(G68), .C2(new_n751), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1014), .B2(new_n681), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1021), .B2(new_n671), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1130), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT124), .Z(G381));
  NAND2_X1  g0946(.A1(new_n1031), .A2(new_n1060), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(G375), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(G390), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n780), .ZN(new_n1150));
  OR2_X1    g0950(.A1(G393), .A2(G396), .ZN(new_n1151));
  NOR4_X1   g0951(.A1(G381), .A2(new_n1150), .A3(G387), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1148), .A2(new_n1152), .ZN(G407));
  NAND2_X1  g0953(.A1(new_n1148), .A2(new_n612), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(G407), .A2(new_n1154), .A3(G213), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT125), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1155), .B(new_n1156), .ZN(G409));
  INV_X1    g0957(.A(G213), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(G343), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT60), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1129), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1129), .A2(new_n1161), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1162), .A2(new_n973), .A3(new_n1029), .A4(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1164), .A2(G384), .A3(new_n1144), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G384), .B1(new_n1164), .B2(new_n1144), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1095), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1168), .A2(new_n1064), .A3(new_n1126), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n668), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1099), .B2(new_n1124), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1084), .A2(new_n1085), .A3(new_n935), .A4(new_n1088), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1147), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1160), .B(new_n1167), .C1(new_n1169), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT62), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1097), .A2(G378), .A3(new_n1127), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1173), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT62), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1178), .A2(new_n1179), .A3(new_n1160), .A4(new_n1167), .ZN(new_n1180));
  OAI211_X1 g0980(.A(G2897), .B(new_n1159), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1166), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1164), .A2(G384), .A3(new_n1144), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1159), .A2(G2897), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1181), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1126), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1173), .B1(new_n1187), .B2(G378), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1186), .B1(new_n1188), .B2(new_n1159), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT61), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1175), .A2(new_n1180), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(G387), .A2(new_n1149), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G390), .B(new_n895), .C1(new_n921), .C2(new_n936), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(G393), .B(G396), .Z(new_n1195));
  INV_X1    g0995(.A(KEYINPUT126), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G387), .B2(new_n1149), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1195), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1192), .A2(new_n1199), .A3(new_n1196), .A4(new_n1193), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1191), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1178), .A2(new_n1160), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT61), .B1(new_n1204), .B2(new_n1186), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT63), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1174), .A2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1178), .A2(KEYINPUT63), .A3(new_n1160), .A4(new_n1167), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1201), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1203), .A2(new_n1209), .ZN(G405));
  NAND2_X1  g1010(.A1(new_n1167), .A2(KEYINPUT127), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1198), .A2(new_n1200), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1167), .A2(KEYINPUT127), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(G375), .A2(new_n1031), .A3(new_n1060), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n1176), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1214), .B(new_n1217), .ZN(G402));
endmodule


