

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575;

  XNOR2_X1 U320 ( .A(n365), .B(n364), .ZN(n366) );
  AND2_X1 U321 ( .A1(G229GAT), .A2(G233GAT), .ZN(n288) );
  NOR2_X1 U322 ( .A1(n554), .A2(n395), .ZN(n397) );
  NOR2_X1 U323 ( .A1(n466), .A2(n517), .ZN(n404) );
  XNOR2_X1 U324 ( .A(n420), .B(KEYINPUT55), .ZN(n421) );
  XNOR2_X1 U325 ( .A(n363), .B(n288), .ZN(n364) );
  XNOR2_X1 U326 ( .A(n422), .B(n421), .ZN(n442) );
  XNOR2_X1 U327 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U328 ( .A(n443), .B(KEYINPUT123), .ZN(n555) );
  XNOR2_X1 U329 ( .A(n372), .B(n371), .ZN(n560) );
  XNOR2_X1 U330 ( .A(n444), .B(G176GAT), .ZN(n445) );
  XNOR2_X1 U331 ( .A(n446), .B(n445), .ZN(G1349GAT) );
  XOR2_X1 U332 ( .A(G141GAT), .B(KEYINPUT24), .Z(n290) );
  NAND2_X1 U333 ( .A1(G228GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U334 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U335 ( .A(KEYINPUT21), .B(G218GAT), .Z(n292) );
  XNOR2_X1 U336 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U338 ( .A(G197GAT), .B(n293), .Z(n313) );
  XOR2_X1 U339 ( .A(n294), .B(n313), .Z(n296) );
  XNOR2_X1 U340 ( .A(G50GAT), .B(G22GAT), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U342 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n298) );
  XNOR2_X1 U343 ( .A(KEYINPUT91), .B(KEYINPUT23), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U345 ( .A(n300), .B(n299), .Z(n309) );
  XNOR2_X1 U346 ( .A(G155GAT), .B(KEYINPUT90), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n301), .B(KEYINPUT2), .ZN(n302) );
  XOR2_X1 U348 ( .A(n302), .B(KEYINPUT3), .Z(n304) );
  XNOR2_X1 U349 ( .A(G148GAT), .B(G162GAT), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n408) );
  XOR2_X1 U351 ( .A(G204GAT), .B(G106GAT), .Z(n306) );
  XNOR2_X1 U352 ( .A(KEYINPUT73), .B(G78GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U354 ( .A(KEYINPUT74), .B(n307), .ZN(n356) );
  XOR2_X1 U355 ( .A(n408), .B(n356), .Z(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n455) );
  XOR2_X1 U357 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n311) );
  XNOR2_X1 U358 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U360 ( .A(KEYINPUT19), .B(n312), .Z(n439) );
  XNOR2_X1 U361 ( .A(n439), .B(n313), .ZN(n324) );
  XOR2_X1 U362 ( .A(G190GAT), .B(KEYINPUT78), .Z(n328) );
  XOR2_X1 U363 ( .A(KEYINPUT79), .B(n328), .Z(n315) );
  XOR2_X1 U364 ( .A(G169GAT), .B(G8GAT), .Z(n358) );
  XNOR2_X1 U365 ( .A(n358), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U367 ( .A(n316), .B(G92GAT), .Z(n322) );
  XNOR2_X1 U368 ( .A(G176GAT), .B(G64GAT), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n317), .B(KEYINPUT76), .ZN(n351) );
  XOR2_X1 U370 ( .A(n351), .B(KEYINPUT94), .Z(n319) );
  NAND2_X1 U371 ( .A1(G226GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U373 ( .A(G36GAT), .B(n320), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n466) );
  XOR2_X1 U376 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n326) );
  XNOR2_X1 U377 ( .A(G218GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U379 ( .A(n327), .B(KEYINPUT9), .Z(n330) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(n328), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n336) );
  XOR2_X1 U382 ( .A(KEYINPUT75), .B(G92GAT), .Z(n332) );
  XNOR2_X1 U383 ( .A(G99GAT), .B(G85GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n345) );
  XOR2_X1 U385 ( .A(G134GAT), .B(n345), .Z(n334) );
  NAND2_X1 U386 ( .A1(G232GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U388 ( .A(n336), .B(n335), .Z(n344) );
  XOR2_X1 U389 ( .A(KEYINPUT8), .B(G50GAT), .Z(n338) );
  XNOR2_X1 U390 ( .A(G43GAT), .B(G36GAT), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U392 ( .A(KEYINPUT7), .B(n339), .Z(n369) );
  XOR2_X1 U393 ( .A(KEYINPUT65), .B(KEYINPUT10), .Z(n341) );
  XNOR2_X1 U394 ( .A(G162GAT), .B(KEYINPUT64), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n369), .B(n342), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n554) );
  XOR2_X1 U398 ( .A(n345), .B(KEYINPUT32), .Z(n347) );
  NAND2_X1 U399 ( .A1(G230GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n355) );
  XOR2_X1 U401 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n349) );
  XNOR2_X1 U402 ( .A(G148GAT), .B(KEYINPUT33), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U404 ( .A(G71GAT), .B(KEYINPUT13), .Z(n376) );
  XOR2_X1 U405 ( .A(n350), .B(n376), .Z(n353) );
  XOR2_X1 U406 ( .A(G120GAT), .B(G57GAT), .Z(n410) );
  XNOR2_X1 U407 ( .A(n410), .B(n351), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n355), .B(n354), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n564) );
  XNOR2_X1 U411 ( .A(KEYINPUT41), .B(n564), .ZN(n541) );
  XOR2_X1 U412 ( .A(KEYINPUT29), .B(G197GAT), .Z(n360) );
  XOR2_X1 U413 ( .A(G22GAT), .B(G15GAT), .Z(n389) );
  XNOR2_X1 U414 ( .A(n358), .B(n389), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n365) );
  XOR2_X1 U416 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n362) );
  XNOR2_X1 U417 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n366), .B(KEYINPUT66), .ZN(n372) );
  XOR2_X1 U420 ( .A(G1GAT), .B(G113GAT), .Z(n368) );
  XNOR2_X1 U421 ( .A(G29GAT), .B(G141GAT), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n409) );
  XOR2_X1 U423 ( .A(n409), .B(KEYINPUT67), .Z(n370) );
  NAND2_X1 U424 ( .A1(n541), .A2(n560), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n373), .B(KEYINPUT46), .ZN(n394) );
  XOR2_X1 U426 ( .A(G64GAT), .B(G78GAT), .Z(n375) );
  XNOR2_X1 U427 ( .A(G127GAT), .B(G155GAT), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U429 ( .A(n377), .B(n376), .Z(n379) );
  XNOR2_X1 U430 ( .A(G183GAT), .B(G211GAT), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n393) );
  XOR2_X1 U432 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n381) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U435 ( .A(KEYINPUT81), .B(KEYINPUT15), .Z(n383) );
  XNOR2_X1 U436 ( .A(KEYINPUT82), .B(KEYINPUT80), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U438 ( .A(n385), .B(n384), .Z(n391) );
  XOR2_X1 U439 ( .A(KEYINPUT79), .B(G57GAT), .Z(n387) );
  XNOR2_X1 U440 ( .A(G1GAT), .B(G8GAT), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U444 ( .A(n393), .B(n392), .ZN(n528) );
  NAND2_X1 U445 ( .A1(n394), .A2(n528), .ZN(n395) );
  XNOR2_X1 U446 ( .A(KEYINPUT47), .B(KEYINPUT109), .ZN(n396) );
  XNOR2_X1 U447 ( .A(n397), .B(n396), .ZN(n402) );
  INV_X1 U448 ( .A(n560), .ZN(n489) );
  XNOR2_X1 U449 ( .A(n489), .B(KEYINPUT71), .ZN(n550) );
  XOR2_X1 U450 ( .A(n554), .B(KEYINPUT36), .Z(n573) );
  NOR2_X1 U451 ( .A1(n573), .A2(n528), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n398), .B(KEYINPUT45), .ZN(n399) );
  NAND2_X1 U453 ( .A1(n399), .A2(n564), .ZN(n400) );
  NOR2_X1 U454 ( .A1(n550), .A2(n400), .ZN(n401) );
  NOR2_X1 U455 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U456 ( .A(KEYINPUT48), .B(n403), .ZN(n517) );
  XNOR2_X1 U457 ( .A(n404), .B(KEYINPUT54), .ZN(n419) );
  XOR2_X1 U458 ( .A(KEYINPUT1), .B(KEYINPUT92), .Z(n406) );
  XNOR2_X1 U459 ( .A(G85GAT), .B(KEYINPUT5), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U461 ( .A(n408), .B(n407), .ZN(n418) );
  XOR2_X1 U462 ( .A(n410), .B(n409), .Z(n412) );
  NAND2_X1 U463 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U465 ( .A(n413), .B(KEYINPUT4), .Z(n416) );
  XNOR2_X1 U466 ( .A(G134GAT), .B(G127GAT), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n414), .B(KEYINPUT0), .ZN(n431) );
  XNOR2_X1 U468 ( .A(n431), .B(KEYINPUT6), .ZN(n415) );
  XNOR2_X1 U469 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U470 ( .A(n418), .B(n417), .ZN(n454) );
  XNOR2_X1 U471 ( .A(KEYINPUT93), .B(n454), .ZN(n457) );
  NAND2_X1 U472 ( .A1(n419), .A2(n457), .ZN(n558) );
  NOR2_X1 U473 ( .A1(n455), .A2(n558), .ZN(n422) );
  XNOR2_X1 U474 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n420) );
  XOR2_X1 U475 ( .A(G71GAT), .B(G15GAT), .Z(n424) );
  XNOR2_X1 U476 ( .A(G169GAT), .B(G113GAT), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n438) );
  XOR2_X1 U478 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n426) );
  XNOR2_X1 U479 ( .A(G99GAT), .B(KEYINPUT86), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U481 ( .A(G176GAT), .B(KEYINPUT20), .Z(n428) );
  XNOR2_X1 U482 ( .A(G120GAT), .B(KEYINPUT83), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U484 ( .A(n430), .B(n429), .Z(n436) );
  XOR2_X1 U485 ( .A(n431), .B(G190GAT), .Z(n433) );
  NAND2_X1 U486 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(n434), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n441) );
  INV_X1 U491 ( .A(n439), .ZN(n440) );
  XOR2_X1 U492 ( .A(n441), .B(n440), .Z(n449) );
  INV_X1 U493 ( .A(n449), .ZN(n521) );
  NAND2_X1 U494 ( .A1(n442), .A2(n521), .ZN(n443) );
  NAND2_X1 U495 ( .A1(n555), .A2(n541), .ZN(n446) );
  XOR2_X1 U496 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n444) );
  XNOR2_X1 U497 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n465) );
  INV_X1 U498 ( .A(n457), .ZN(n507) );
  NOR2_X1 U499 ( .A1(n449), .A2(n466), .ZN(n447) );
  NOR2_X1 U500 ( .A1(n455), .A2(n447), .ZN(n448) );
  XOR2_X1 U501 ( .A(KEYINPUT25), .B(n448), .Z(n452) );
  XNOR2_X1 U502 ( .A(n466), .B(KEYINPUT27), .ZN(n456) );
  NAND2_X1 U503 ( .A1(n455), .A2(n449), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n450), .B(KEYINPUT26), .ZN(n559) );
  NOR2_X1 U505 ( .A1(n456), .A2(n559), .ZN(n451) );
  NOR2_X1 U506 ( .A1(n452), .A2(n451), .ZN(n453) );
  NOR2_X1 U507 ( .A1(n454), .A2(n453), .ZN(n460) );
  XNOR2_X1 U508 ( .A(n455), .B(KEYINPUT28), .ZN(n519) );
  OR2_X1 U509 ( .A1(n521), .A2(n519), .ZN(n458) );
  OR2_X1 U510 ( .A1(n457), .A2(n456), .ZN(n516) );
  NOR2_X1 U511 ( .A1(n458), .A2(n516), .ZN(n459) );
  NOR2_X1 U512 ( .A1(n460), .A2(n459), .ZN(n474) );
  NOR2_X1 U513 ( .A1(n554), .A2(n528), .ZN(n461) );
  XOR2_X1 U514 ( .A(KEYINPUT16), .B(n461), .Z(n462) );
  NOR2_X1 U515 ( .A1(n474), .A2(n462), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(KEYINPUT95), .ZN(n491) );
  NAND2_X1 U517 ( .A1(n550), .A2(n564), .ZN(n478) );
  NOR2_X1 U518 ( .A1(n491), .A2(n478), .ZN(n472) );
  NAND2_X1 U519 ( .A1(n507), .A2(n472), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n465), .B(n464), .ZN(G1324GAT) );
  INV_X1 U521 ( .A(n466), .ZN(n509) );
  NAND2_X1 U522 ( .A1(n509), .A2(n472), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n467), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U524 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n469) );
  NAND2_X1 U525 ( .A1(n472), .A2(n521), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(n471) );
  XOR2_X1 U527 ( .A(G15GAT), .B(KEYINPUT96), .Z(n470) );
  XNOR2_X1 U528 ( .A(n471), .B(n470), .ZN(G1326GAT) );
  NAND2_X1 U529 ( .A1(n519), .A2(n472), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U531 ( .A(G29GAT), .B(KEYINPUT39), .Z(n481) );
  XOR2_X1 U532 ( .A(KEYINPUT98), .B(KEYINPUT37), .Z(n477) );
  NOR2_X1 U533 ( .A1(n573), .A2(n474), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n475), .A2(n528), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(n505) );
  NOR2_X1 U536 ( .A1(n505), .A2(n478), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT38), .B(n479), .ZN(n486) );
  NAND2_X1 U538 ( .A1(n507), .A2(n486), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1328GAT) );
  NAND2_X1 U540 ( .A1(n486), .A2(n509), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT40), .B(KEYINPUT99), .Z(n484) );
  NAND2_X1 U543 ( .A1(n486), .A2(n521), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U545 ( .A(G43GAT), .B(n485), .ZN(G1330GAT) );
  NAND2_X1 U546 ( .A1(n486), .A2(n519), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n487), .B(KEYINPUT100), .ZN(n488) );
  XNOR2_X1 U548 ( .A(G50GAT), .B(n488), .ZN(G1331GAT) );
  XNOR2_X1 U549 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n494) );
  NAND2_X1 U550 ( .A1(n541), .A2(n489), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT101), .B(n490), .Z(n504) );
  NOR2_X1 U552 ( .A1(n504), .A2(n491), .ZN(n492) );
  XNOR2_X1 U553 ( .A(KEYINPUT102), .B(n492), .ZN(n501) );
  NAND2_X1 U554 ( .A1(n507), .A2(n501), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1332GAT) );
  XOR2_X1 U556 ( .A(G64GAT), .B(KEYINPUT103), .Z(n496) );
  NAND2_X1 U557 ( .A1(n501), .A2(n509), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1333GAT) );
  NAND2_X1 U559 ( .A1(n501), .A2(n521), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n499) );
  XNOR2_X1 U562 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U564 ( .A(KEYINPUT104), .B(n500), .Z(n503) );
  NAND2_X1 U565 ( .A1(n501), .A2(n519), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  NOR2_X1 U567 ( .A1(n505), .A2(n504), .ZN(n506) );
  XOR2_X1 U568 ( .A(KEYINPUT107), .B(n506), .Z(n512) );
  NAND2_X1 U569 ( .A1(n507), .A2(n512), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G85GAT), .B(n508), .ZN(G1336GAT) );
  NAND2_X1 U571 ( .A1(n509), .A2(n512), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n510), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U573 ( .A1(n521), .A2(n512), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n514) );
  NAND2_X1 U576 ( .A1(n512), .A2(n519), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U578 ( .A(G106GAT), .B(n515), .Z(G1339GAT) );
  NOR2_X1 U579 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U580 ( .A(KEYINPUT110), .B(n518), .Z(n536) );
  NOR2_X1 U581 ( .A1(n536), .A2(n519), .ZN(n520) );
  NAND2_X1 U582 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U583 ( .A(n522), .B(KEYINPUT111), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n550), .A2(n531), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n523), .B(KEYINPUT112), .ZN(n524) );
  XNOR2_X1 U586 ( .A(G113GAT), .B(n524), .ZN(G1340GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n526) );
  NAND2_X1 U588 ( .A1(n531), .A2(n541), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U590 ( .A(G120GAT), .B(n527), .Z(G1341GAT) );
  INV_X1 U591 ( .A(n528), .ZN(n568) );
  NAND2_X1 U592 ( .A1(n531), .A2(n568), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(KEYINPUT50), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G127GAT), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n533) );
  NAND2_X1 U596 ( .A1(n531), .A2(n554), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n535) );
  XOR2_X1 U598 ( .A(G134GAT), .B(KEYINPUT115), .Z(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1343GAT) );
  NOR2_X1 U600 ( .A1(n559), .A2(n536), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n537), .B(KEYINPUT116), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n560), .A2(n548), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G141GAT), .B(n538), .ZN(G1344GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n540) );
  XNOR2_X1 U605 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n545) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n548), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1345GAT) );
  NAND2_X1 U611 ( .A1(n548), .A2(n568), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT120), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  NAND2_X1 U614 ( .A1(n548), .A2(n554), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n555), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(KEYINPUT124), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n552), .ZN(G1348GAT) );
  NAND2_X1 U619 ( .A1(n555), .A2(n568), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT58), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G190GAT), .B(n557), .ZN(G1351GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n562) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n569), .A2(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(n563), .ZN(G1352GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n566) );
  INV_X1 U630 ( .A(n569), .ZN(n572) );
  OR2_X1 U631 ( .A1(n572), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(G204GAT), .B(n567), .Z(G1353GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(KEYINPUT126), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G211GAT), .B(n571), .ZN(G1354GAT) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT62), .B(n574), .Z(n575) );
  XNOR2_X1 U639 ( .A(G218GAT), .B(n575), .ZN(G1355GAT) );
endmodule

