//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT86), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT77), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(G141gat), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n207), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(G141gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT78), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT78), .A4(new_n209), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n214), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n207), .A2(G148gat), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT2), .B1(new_n225), .B2(new_n209), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n226), .A2(new_n217), .A3(new_n219), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT79), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n227), .B1(new_n214), .B2(new_n222), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT79), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(new_n224), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT29), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT74), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G211gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(G218gat), .ZN(new_n239));
  INV_X1    g038(.A(G218gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(G211gat), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT74), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT73), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT72), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n238), .ZN(new_n246));
  NAND2_X1  g045(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n240), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n244), .B1(new_n248), .B2(KEYINPUT22), .ZN(new_n249));
  AND2_X1   g048(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n251));
  OAI21_X1  g050(.A(G218gat), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT22), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(KEYINPUT73), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G197gat), .B(G204gat), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n243), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n252), .A2(KEYINPUT73), .A3(new_n253), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT73), .B1(new_n252), .B2(new_n253), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n243), .B(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(KEYINPUT75), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT75), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n256), .B1(new_n249), .B2(new_n254), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n265), .B2(new_n243), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n259), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n203), .B1(new_n234), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT29), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n232), .B1(new_n231), .B2(new_n224), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n212), .A2(new_n213), .B1(new_n218), .B2(new_n221), .ZN(new_n271));
  NOR4_X1   g070(.A1(new_n271), .A2(KEYINPUT79), .A3(new_n227), .A4(KEYINPUT3), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n269), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n262), .A2(KEYINPUT75), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n255), .A2(new_n264), .A3(new_n243), .A4(new_n257), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n258), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(KEYINPUT86), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n202), .B1(new_n268), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n267), .A2(KEYINPUT85), .A3(new_n269), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT85), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(new_n276), .B2(KEYINPUT29), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n281), .A3(new_n224), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n223), .A2(new_n228), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n263), .A2(new_n266), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT84), .B1(new_n265), .B2(new_n243), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT84), .ZN(new_n289));
  INV_X1    g088(.A(new_n243), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n269), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n231), .B1(new_n293), .B2(new_n224), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n273), .A2(new_n276), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n202), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(KEYINPUT87), .B(G22gat), .Z(new_n298));
  NAND3_X1  g097(.A1(new_n285), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G78gat), .B(G106gat), .ZN(new_n300));
  INV_X1    g099(.A(G50gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n287), .B(new_n291), .C1(new_n263), .C2(new_n266), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT3), .B1(new_n307), .B2(new_n269), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n295), .B1(new_n308), .B2(new_n231), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n278), .A2(new_n284), .B1(new_n309), .B2(new_n202), .ZN(new_n310));
  OR2_X1    g109(.A1(KEYINPUT87), .A2(G22gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G22gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(KEYINPUT88), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n282), .A2(new_n283), .ZN(new_n317));
  INV_X1    g116(.A(new_n202), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n234), .A2(new_n203), .A3(new_n267), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT86), .B1(new_n273), .B2(new_n276), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n297), .B(new_n316), .C1(new_n317), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n304), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n285), .B2(new_n297), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n305), .B1(new_n310), .B2(new_n316), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n297), .B1(new_n317), .B2(new_n321), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n315), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT89), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n313), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n230), .A2(new_n233), .ZN(new_n332));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(KEYINPUT1), .ZN(new_n334));
  XOR2_X1   g133(.A(G127gat), .B(G134gat), .Z(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n336), .B1(new_n283), .B2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g136(.A(new_n336), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT4), .B1(new_n283), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n231), .A2(new_n340), .A3(new_n336), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n332), .A2(new_n337), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n343));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n342), .A2(KEYINPUT81), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n337), .B1(new_n270), .B2(new_n272), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n339), .A2(new_n341), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n343), .A4(new_n344), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G1gat), .B(G29gat), .Z(new_n352));
  XNOR2_X1  g151(.A(G57gat), .B(G85gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n344), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n231), .B(new_n336), .ZN(new_n359));
  INV_X1    g158(.A(new_n344), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n343), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n351), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n351), .A2(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n356), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT6), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n345), .A2(new_n350), .B1(new_n358), .B2(new_n361), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(new_n357), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(KEYINPUT82), .A3(new_n357), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT24), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(G183gat), .A3(G190gat), .ZN(new_n375));
  INV_X1    g174(.A(G183gat), .ZN(new_n376));
  INV_X1    g175(.A(G190gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n375), .B1(new_n378), .B2(new_n374), .ZN(new_n379));
  NOR2_X1   g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT23), .ZN(new_n384));
  NAND2_X1  g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT23), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(G169gat), .B2(G176gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT25), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n380), .B(KEYINPUT64), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n379), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT65), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n391), .B(new_n393), .C1(new_n388), .C2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT27), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G183gat), .ZN(new_n397));
  AOI21_X1  g196(.A(G190gat), .B1(new_n397), .B2(KEYINPUT66), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT27), .B(G183gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(KEYINPUT66), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT28), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(G190gat), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n400), .A2(new_n401), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n378), .B1(KEYINPUT26), .B2(new_n383), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT26), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n383), .B2(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n389), .B(new_n395), .C1(new_n403), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n269), .ZN(new_n409));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n410), .B(KEYINPUT76), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n389), .A2(new_n395), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n403), .A2(new_n407), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n411), .B(new_n267), .C1(new_n413), .C2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n410), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n412), .B1(new_n408), .B2(new_n269), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n276), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G64gat), .B(G92gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n422), .B(new_n423), .Z(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n417), .A2(new_n420), .A3(new_n424), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(KEYINPUT30), .A3(new_n427), .ZN(new_n428));
  OR3_X1    g227(.A1(new_n421), .A2(KEYINPUT30), .A3(new_n425), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n368), .A2(new_n373), .A3(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(G15gat), .B(G43gat), .Z(new_n433));
  XNOR2_X1  g232(.A(G71gat), .B(G99gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G227gat), .A2(G233gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n416), .A2(new_n336), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n408), .A2(new_n338), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT32), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n441), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n408), .A2(new_n338), .ZN(new_n446));
  OAI211_X1 g245(.A(G227gat), .B(G233gat), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT67), .B(KEYINPUT33), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(KEYINPUT68), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT68), .ZN(new_n450));
  INV_X1    g249(.A(new_n448), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n450), .B1(new_n442), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n444), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n447), .A2(KEYINPUT32), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n437), .A2(new_n448), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n439), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT34), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n439), .B2(KEYINPUT71), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n457), .B(new_n459), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n453), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n460), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n437), .B1(new_n447), .B2(KEYINPUT32), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT68), .B1(new_n447), .B2(new_n448), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n442), .A2(new_n450), .A3(new_n451), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n454), .A2(new_n455), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n331), .A2(new_n432), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT35), .ZN(new_n471));
  INV_X1    g270(.A(new_n469), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n324), .B1(new_n323), .B2(new_n325), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT89), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n475), .B2(new_n313), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT35), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n432), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n425), .B1(new_n421), .B2(KEYINPUT37), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n421), .A2(KEYINPUT37), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n411), .B1(new_n413), .B2(new_n416), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT37), .B1(new_n485), .B2(new_n267), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n418), .A2(new_n419), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(new_n276), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n480), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n427), .B1(new_n489), .B2(new_n481), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(new_n368), .B2(new_n373), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n346), .A2(new_n347), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n360), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n357), .B1(new_n494), .B2(KEYINPUT39), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT39), .B1(new_n359), .B2(new_n360), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n493), .B2(new_n360), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  OAI22_X1  g298(.A1(new_n495), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n501), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(new_n431), .A3(new_n367), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n331), .A2(new_n492), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n306), .A2(new_n312), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(new_n473), .B2(new_n474), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n371), .B1(new_n363), .B2(new_n364), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n367), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT82), .B1(new_n369), .B2(new_n357), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n371), .B1(new_n510), .B2(new_n370), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n511), .A3(new_n430), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n460), .B1(new_n453), .B2(new_n456), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n466), .A2(new_n462), .A3(new_n467), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT36), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT36), .B1(new_n514), .B2(new_n515), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n505), .B(new_n513), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n479), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n522), .A2(new_n523), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(new_n523), .B2(new_n522), .ZN(new_n525));
  OR3_X1    g324(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n528), .B(KEYINPUT95), .Z(new_n531));
  OAI21_X1  g330(.A(KEYINPUT96), .B1(new_n527), .B2(KEYINPUT15), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n527), .A2(KEYINPUT96), .A3(KEYINPUT15), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(G29gat), .B2(G36gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n522), .A2(new_n526), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n531), .A2(new_n532), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT17), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  INV_X1    g341(.A(G85gat), .ZN(new_n543));
  INV_X1    g342(.A(G92gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(KEYINPUT8), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g345(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n546), .A2(G85gat), .A3(G92gat), .A4(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n546), .A2(new_n547), .B1(G85gat), .B2(G92gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT100), .ZN(new_n552));
  XNOR2_X1  g351(.A(G99gat), .B(G106gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n551), .A2(new_n554), .ZN(new_n556));
  INV_X1    g355(.A(new_n545), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT99), .B(KEYINPUT7), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n543), .B2(new_n544), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n559), .B2(new_n548), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n553), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n561), .A3(KEYINPUT100), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n539), .A2(new_n541), .A3(new_n555), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n555), .ZN(new_n564));
  AND2_X1   g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n537), .A2(new_n564), .B1(KEYINPUT41), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n566), .A2(KEYINPUT101), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(KEYINPUT101), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n563), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n565), .A2(KEYINPUT41), .ZN(new_n572));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n571), .B(new_n574), .Z(new_n575));
  XOR2_X1   g374(.A(G57gat), .B(G64gat), .Z(new_n576));
  INV_X1    g375(.A(G71gat), .ZN(new_n577));
  INV_X1    g376(.A(G78gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n576), .B1(KEYINPUT9), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G71gat), .B(G78gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT21), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  XNOR2_X1  g385(.A(G15gat), .B(G22gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT16), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(G1gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(G1gat), .B2(new_n587), .ZN(new_n590));
  INV_X1    g389(.A(G8gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n582), .B2(new_n583), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n586), .B(new_n593), .Z(new_n594));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT98), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n594), .B(new_n600), .Z(new_n601));
  NOR2_X1   g400(.A1(new_n575), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT10), .ZN(new_n603));
  AOI211_X1 g402(.A(new_n603), .B(new_n582), .C1(new_n562), .C2(new_n555), .ZN(new_n604));
  INV_X1    g403(.A(new_n556), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n551), .A2(new_n554), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n605), .A2(new_n582), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n562), .A2(new_n582), .A3(new_n555), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT102), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n562), .A2(new_n610), .A3(new_n582), .A4(new_n555), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n604), .B1(new_n612), .B2(new_n603), .ZN(new_n613));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n614), .B(KEYINPUT103), .Z(new_n615));
  OAI21_X1  g414(.A(KEYINPUT104), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n617));
  INV_X1    g416(.A(new_n615), .ZN(new_n618));
  AOI211_X1 g417(.A(KEYINPUT10), .B(new_n607), .C1(new_n609), .C2(new_n611), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n604), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n612), .A2(new_n618), .ZN(new_n621));
  XOR2_X1   g420(.A(G120gat), .B(G148gat), .Z(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n616), .A2(new_n620), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n624), .B(KEYINPUT105), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n615), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n628), .B1(new_n629), .B2(new_n621), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n602), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n592), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n537), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n541), .A2(new_n592), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n537), .A2(new_n540), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n634), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT18), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n539), .A2(new_n592), .A3(new_n541), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n642), .A2(KEYINPUT18), .A3(new_n634), .A4(new_n636), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n537), .B(new_n635), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n634), .B(KEYINPUT13), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n641), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G113gat), .B(G141gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G169gat), .B(G197gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT92), .Z(new_n654));
  NAND2_X1  g453(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT97), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n641), .A2(new_n643), .A3(new_n646), .A4(new_n653), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT97), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n647), .A2(new_n658), .A3(new_n654), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n633), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n519), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n509), .A2(new_n511), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g466(.A1(new_n663), .A2(new_n430), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT42), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT106), .B1(new_n668), .B2(new_n591), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n668), .A2(KEYINPUT106), .A3(new_n591), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT107), .ZN(G1325gat));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n516), .B2(new_n517), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT36), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n461), .B2(new_n468), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT36), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(KEYINPUT108), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G15gat), .B1(new_n663), .B2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n472), .A2(G15gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n663), .B2(new_n684), .ZN(G1326gat));
  NOR2_X1   g484(.A1(new_n663), .A2(new_n331), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT109), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT43), .B(G22gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  XNOR2_X1  g488(.A(new_n571), .B(new_n574), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n479), .B2(new_n518), .ZN(new_n691));
  INV_X1    g490(.A(new_n601), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n661), .A2(new_n692), .A3(new_n631), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n665), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT45), .Z(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(KEYINPUT44), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n693), .B(KEYINPUT110), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n477), .B1(new_n476), .B2(new_n432), .ZN(new_n699));
  NOR4_X1   g498(.A1(new_n507), .A2(new_n512), .A3(new_n472), .A4(KEYINPUT35), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT112), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT112), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n471), .A2(new_n702), .A3(new_n478), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n505), .A2(new_n513), .A3(new_n682), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n505), .A2(new_n682), .A3(KEYINPUT111), .A4(new_n513), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n690), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n697), .B(new_n698), .C1(new_n711), .C2(KEYINPUT44), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n665), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n713), .ZN(G1328gat));
  OAI21_X1  g513(.A(G36gat), .B1(new_n712), .B2(new_n430), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n694), .A2(G36gat), .A3(new_n430), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(G1329gat));
  INV_X1    g517(.A(new_n694), .ZN(new_n719));
  AOI21_X1  g518(.A(G43gat), .B1(new_n719), .B2(new_n469), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n682), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G43gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n712), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g524(.A(G50gat), .B1(new_n719), .B2(new_n507), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n331), .A2(new_n301), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n712), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n703), .A3(new_n701), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n660), .A2(new_n632), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(new_n601), .A3(new_n575), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n665), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT113), .B(G57gat), .Z(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1332gat));
  NOR2_X1   g538(.A1(new_n736), .A2(new_n430), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n740), .B2(new_n741), .ZN(G1333gat));
  NOR3_X1   g543(.A1(new_n736), .A2(G71gat), .A3(new_n472), .ZN(new_n745));
  INV_X1    g544(.A(new_n736), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n722), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(G71gat), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g548(.A1(new_n736), .A2(new_n331), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n578), .ZN(G1335gat));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n708), .A2(new_n709), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n753), .B(new_n575), .C1(new_n754), .C2(new_n704), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n660), .A2(new_n692), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n753), .B1(new_n732), .B2(new_n575), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n752), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n575), .B1(new_n754), .B2(new_n704), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT115), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n761), .A2(KEYINPUT51), .A3(new_n755), .A4(new_n756), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(new_n543), .A3(new_n664), .A4(new_n631), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n734), .A2(new_n692), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n697), .B(new_n765), .C1(new_n711), .C2(KEYINPUT44), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n766), .A2(KEYINPUT114), .A3(new_n665), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT114), .B1(new_n766), .B2(new_n665), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G85gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n764), .B1(new_n767), .B2(new_n769), .ZN(G1336gat));
  NOR2_X1   g569(.A1(new_n632), .A2(new_n430), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n544), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n759), .B2(new_n762), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  OAI21_X1  g574(.A(G92gat), .B1(new_n766), .B2(new_n430), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n776), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT52), .B1(new_n778), .B2(new_n773), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1337gat));
  NOR2_X1   g579(.A1(new_n472), .A2(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n631), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G99gat), .B1(new_n766), .B2(new_n682), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1338gat));
  XNOR2_X1  g583(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n331), .A2(G106gat), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  AOI211_X1 g587(.A(new_n632), .B(new_n788), .C1(new_n759), .C2(new_n762), .ZN(new_n789));
  OAI21_X1  g588(.A(G106gat), .B1(new_n766), .B2(new_n331), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n786), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n763), .A2(new_n631), .A3(new_n787), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n790), .A3(new_n785), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1339gat));
  INV_X1    g594(.A(G113gat), .ZN(new_n796));
  INV_X1    g595(.A(new_n627), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n613), .A2(new_n615), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n616), .A2(KEYINPUT54), .A3(new_n620), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n624), .B1(new_n629), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n797), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n799), .A2(new_n801), .A3(KEYINPUT55), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n660), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n634), .B1(new_n642), .B2(new_n636), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n644), .A2(new_n645), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n652), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n631), .A2(new_n657), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n575), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n804), .A2(new_n805), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n657), .A2(new_n809), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n812), .A2(new_n690), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n601), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n602), .A2(new_n661), .A3(new_n632), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n507), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n665), .A2(new_n431), .A3(new_n472), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n796), .B1(new_n819), .B2(new_n660), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT118), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n815), .A2(new_n816), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n664), .ZN(new_n823));
  INV_X1    g622(.A(new_n476), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n823), .A2(new_n431), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n796), .A3(new_n660), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n821), .A2(new_n826), .ZN(G1340gat));
  AOI21_X1  g626(.A(G120gat), .B1(new_n825), .B2(new_n631), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n631), .A2(G120gat), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n819), .B2(new_n829), .ZN(G1341gat));
  NAND3_X1  g629(.A1(new_n819), .A2(G127gat), .A3(new_n692), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT119), .ZN(new_n832));
  AOI21_X1  g631(.A(G127gat), .B1(new_n825), .B2(new_n692), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(G1342gat));
  NOR2_X1   g633(.A1(new_n690), .A2(new_n431), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OR4_X1    g635(.A1(G134gat), .A2(new_n823), .A3(new_n824), .A4(new_n836), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n838));
  INV_X1    g637(.A(new_n819), .ZN(new_n839));
  OAI21_X1  g638(.A(G134gat), .B1(new_n839), .B2(new_n690), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(G1343gat));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n682), .A2(new_n664), .A3(new_n430), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n331), .B1(new_n815), .B2(new_n816), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n848), .B1(new_n804), .B2(new_n805), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n804), .A2(new_n848), .A3(new_n805), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n660), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n575), .B1(new_n852), .B2(new_n810), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n601), .B1(new_n853), .B2(new_n814), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n331), .B1(new_n854), .B2(new_n816), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n660), .B(new_n847), .C1(new_n855), .C2(new_n846), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n722), .A2(KEYINPUT121), .A3(new_n331), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n859), .B1(new_n682), .B2(new_n507), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n822), .A3(new_n664), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n661), .A2(G141gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n430), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n843), .B1(new_n857), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n862), .A2(KEYINPUT122), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n861), .A2(new_n822), .A3(new_n870), .A4(new_n664), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n869), .A2(new_n430), .A3(new_n864), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n843), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(G141gat), .B2(new_n856), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT123), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n857), .A2(new_n843), .A3(new_n872), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n856), .A2(G141gat), .B1(new_n863), .B2(new_n866), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n876), .B(new_n877), .C1(new_n843), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(G1344gat));
  OAI21_X1  g679(.A(new_n847), .B1(new_n855), .B2(new_n846), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(new_n632), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n882), .A2(new_n883), .A3(G148gat), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n804), .A2(new_n848), .A3(new_n805), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(new_n849), .A3(new_n661), .ZN(new_n886));
  INV_X1    g685(.A(new_n810), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n690), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n814), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n692), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n816), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n846), .B(new_n507), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n845), .A2(new_n846), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n844), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n631), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n883), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n869), .A2(new_n871), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n430), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n631), .A2(new_n205), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n884), .A2(new_n897), .B1(new_n899), .B2(new_n900), .ZN(G1345gat));
  OAI21_X1  g700(.A(G155gat), .B1(new_n881), .B2(new_n601), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n692), .A2(new_n215), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n899), .B2(new_n903), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n881), .B2(new_n690), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n898), .A2(new_n216), .A3(new_n835), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1347gat));
  AOI21_X1  g706(.A(new_n664), .B1(new_n815), .B2(new_n816), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n476), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n430), .ZN(new_n910));
  AOI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n660), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n664), .A2(new_n430), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n472), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n817), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n660), .A2(G169gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(G1348gat));
  AND2_X1   g716(.A1(new_n915), .A2(new_n631), .ZN(new_n918));
  INV_X1    g717(.A(G176gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n771), .A2(new_n919), .ZN(new_n920));
  OAI22_X1  g719(.A1(new_n918), .A2(new_n919), .B1(new_n909), .B2(new_n920), .ZN(G1349gat));
  AOI21_X1  g720(.A(new_n376), .B1(new_n915), .B2(new_n692), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n922), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n910), .A2(new_n399), .A3(new_n692), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n925), .B(new_n926), .Z(G1350gat));
  AOI21_X1  g726(.A(new_n377), .B1(new_n915), .B2(new_n575), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT61), .Z(new_n929));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n377), .A3(new_n575), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1351gat));
  AND3_X1   g730(.A1(new_n908), .A2(new_n507), .A3(new_n682), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(KEYINPUT125), .A3(new_n431), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT125), .B1(new_n932), .B2(new_n431), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n660), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n722), .A2(new_n913), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n894), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n938), .A2(new_n939), .A3(new_n661), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n936), .A2(new_n940), .ZN(G1352gat));
  INV_X1    g740(.A(G204gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n932), .A2(new_n942), .A3(new_n771), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT62), .Z(new_n944));
  OAI21_X1  g743(.A(KEYINPUT126), .B1(new_n938), .B2(new_n632), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G204gat), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n938), .A2(KEYINPUT126), .A3(new_n632), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1353gat));
  NOR3_X1   g747(.A1(new_n601), .A2(new_n251), .A3(new_n250), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n949), .B1(new_n933), .B2(new_n934), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n892), .A2(new_n692), .A3(new_n893), .A4(new_n937), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n951), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n951), .B2(G211gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n950), .B(new_n956), .C1(new_n952), .C2(new_n953), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1354gat));
  NAND3_X1  g757(.A1(new_n935), .A2(new_n240), .A3(new_n575), .ZN(new_n959));
  OAI21_X1  g758(.A(G218gat), .B1(new_n938), .B2(new_n690), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1355gat));
endmodule


