//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1268, new_n1269,
    new_n1270;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT64), .Z(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT65), .B(G244), .Z(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G107), .A2(G264), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n215), .B1(new_n218), .B2(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  AOI21_X1  g0046(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n247));
  INV_X1    g0047(.A(G274), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n252), .A2(new_n249), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n250), .B1(G226), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G222), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G223), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n259), .B(new_n247), .C1(G77), .C2(new_n255), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G190), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n216), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n268), .A2(new_n269), .B1(new_n202), .B2(new_n265), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT8), .B(G58), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n210), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G150), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI22_X1  g0075(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(G20), .B2(new_n203), .ZN(new_n277));
  INV_X1    g0077(.A(new_n267), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n270), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT9), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(KEYINPUT9), .B(new_n270), .C1(new_n277), .C2(new_n278), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n261), .A2(G200), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n263), .A2(new_n281), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT10), .ZN(new_n285));
  INV_X1    g0085(.A(G179), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n262), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(new_n279), .C1(G169), .C2(new_n262), .ZN(new_n288));
  INV_X1    g0088(.A(new_n271), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n289), .A2(new_n274), .B1(G20), .B2(G77), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT15), .B(G87), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n291), .A2(new_n272), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n267), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n209), .A2(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n268), .A2(G77), .A3(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n294), .B(new_n296), .C1(G77), .C2(new_n264), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n255), .A2(G238), .A3(G1698), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n255), .A2(G232), .A3(new_n257), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n298), .B(new_n299), .C1(new_n206), .C2(new_n255), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n247), .ZN(new_n301));
  INV_X1    g0101(.A(new_n220), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n250), .B1(new_n302), .B2(new_n253), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n297), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n304), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n286), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n297), .B1(new_n304), .B2(G200), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(G190), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n285), .A2(new_n288), .A3(new_n310), .A4(new_n313), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n275), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n272), .A2(new_n221), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n267), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT11), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n264), .A2(G68), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT12), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n321), .A2(KEYINPUT69), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(KEYINPUT69), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n322), .B(new_n323), .C1(new_n320), .C2(new_n319), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n268), .A2(G68), .A3(new_n295), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n318), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n250), .B1(G238), .B2(new_n253), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n257), .A2(G232), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n255), .B(new_n330), .C1(G226), .C2(G1698), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G97), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n252), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n327), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n333), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(new_n328), .A3(KEYINPUT13), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n336), .A3(G169), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(KEYINPUT70), .A3(KEYINPUT14), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n329), .A2(new_n333), .B1(KEYINPUT68), .B2(new_n327), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT68), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n335), .A2(new_n328), .A3(new_n340), .A4(KEYINPUT13), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G179), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n337), .B1(KEYINPUT70), .B2(KEYINPUT14), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n326), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n334), .A2(new_n336), .A3(G200), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT67), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n326), .B1(G190), .B2(new_n342), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n314), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G58), .ZN(new_n353));
  INV_X1    g0153(.A(G68), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(G20), .B1(new_n355), .B2(new_n201), .ZN(new_n356));
  INV_X1    g0156(.A(G159), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(new_n275), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT3), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G33), .ZN(new_n360));
  INV_X1    g0160(.A(G33), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(G20), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(G20), .B1(new_n360), .B2(new_n362), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(KEYINPUT7), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n358), .B1(new_n368), .B2(G68), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n278), .B1(new_n369), .B2(KEYINPUT16), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT71), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n367), .B2(KEYINPUT7), .ZN(new_n372));
  OAI211_X1 g0172(.A(KEYINPUT71), .B(new_n364), .C1(new_n255), .C2(G20), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n361), .B2(KEYINPUT3), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n359), .A2(KEYINPUT72), .A3(G33), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(new_n362), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n365), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT73), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n378), .A2(KEYINPUT73), .A3(new_n365), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n374), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n358), .B1(new_n383), .B2(G68), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n370), .B1(new_n384), .B2(KEYINPUT16), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT74), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n370), .C1(new_n384), .C2(KEYINPUT16), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n268), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n289), .A2(new_n295), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n390), .A2(new_n391), .B1(new_n264), .B2(new_n289), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n250), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n253), .A2(G232), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n257), .A2(G226), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n255), .B(new_n397), .C1(G223), .C2(G1698), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n252), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G190), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G200), .B2(new_n401), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n403), .B(KEYINPUT75), .C1(G200), .C2(new_n401), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND4_X1   g0208(.A1(KEYINPUT17), .A2(new_n389), .A3(new_n393), .A4(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n392), .B1(new_n386), .B2(new_n388), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT17), .B1(new_n410), .B2(new_n408), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  INV_X1    g0213(.A(new_n379), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(KEYINPUT73), .B1(new_n372), .B2(new_n373), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n354), .B1(new_n415), .B2(new_n381), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n413), .B1(new_n416), .B2(new_n358), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n387), .B1(new_n417), .B2(new_n370), .ZN(new_n418));
  INV_X1    g0218(.A(new_n388), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n393), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n401), .A2(new_n305), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(G179), .B2(new_n401), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(KEYINPUT18), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n410), .B2(new_n422), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n352), .A2(new_n412), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n264), .A2(G97), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n361), .A2(G1), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n265), .A2(new_n267), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n429), .B1(new_n431), .B2(G97), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G97), .A2(G107), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT6), .B1(new_n207), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n436), .A2(new_n210), .B1(new_n221), .B2(new_n275), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n383), .B2(G107), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n432), .B1(new_n438), .B2(new_n278), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT76), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT5), .B(G41), .ZN(new_n441));
  INV_X1    g0241(.A(G45), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G1), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n441), .A2(G274), .A3(new_n252), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n247), .B1(new_n443), .B2(new_n441), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n445), .B1(G257), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n360), .A2(new_n362), .A3(G250), .A4(G1698), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n360), .A2(new_n362), .A3(G244), .A4(new_n257), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT4), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT4), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n255), .A2(new_n453), .A3(G244), .A4(new_n257), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n450), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n247), .B1(new_n455), .B2(KEYINPUT77), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n452), .A2(new_n454), .ZN(new_n457));
  INV_X1    g0257(.A(new_n450), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT77), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n402), .B(new_n447), .C1(new_n456), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n447), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n252), .B1(new_n459), .B2(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n455), .A2(KEYINPUT77), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n462), .B1(new_n466), .B2(G200), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT76), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n432), .C1(new_n438), .C2(new_n278), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n440), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(G179), .B(new_n447), .C1(new_n456), .C2(new_n461), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n466), .B2(new_n305), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n439), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n360), .A2(new_n362), .A3(G244), .A4(G1698), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n360), .A2(new_n362), .A3(G238), .A4(new_n257), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n474), .B(new_n475), .C1(new_n361), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n247), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n252), .A2(G274), .A3(new_n443), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n209), .A2(G45), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n252), .A2(G250), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(new_n286), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT78), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n478), .A2(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n305), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n255), .A2(new_n210), .A3(G68), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT19), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n210), .B1(new_n332), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(G87), .B2(new_n207), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n272), .B2(new_n205), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n267), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n291), .A2(new_n265), .ZN(new_n496));
  INV_X1    g0296(.A(new_n431), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(new_n496), .C1(new_n291), .C2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n482), .B1(new_n477), .B2(new_n247), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(KEYINPUT78), .A3(new_n286), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n486), .A2(new_n488), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n431), .A2(G87), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n495), .A2(new_n496), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n487), .A2(G200), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n503), .B(new_n504), .C1(new_n402), .C2(new_n487), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n470), .A2(new_n473), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT79), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT79), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n470), .A2(new_n509), .A3(new_n473), .A4(new_n506), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT25), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n264), .B2(G107), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n264), .A2(new_n512), .A3(G107), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT81), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(KEYINPUT81), .B(new_n512), .C1(new_n264), .C2(G107), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n516), .A2(new_n517), .B1(G107), .B2(new_n431), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n360), .A2(new_n362), .A3(new_n210), .A4(G87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT22), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT22), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n255), .A2(new_n522), .A3(new_n210), .A4(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n361), .A2(new_n476), .A3(G20), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT23), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n210), .B2(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT24), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n524), .A2(new_n532), .A3(new_n529), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n519), .B1(new_n534), .B2(new_n267), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT82), .ZN(new_n536));
  AND2_X1   g0336(.A1(KEYINPUT5), .A2(G41), .ZN(new_n537));
  NOR2_X1   g0337(.A1(KEYINPUT5), .A2(G41), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n443), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n252), .ZN(new_n540));
  INV_X1    g0340(.A(G264), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n539), .A2(KEYINPUT82), .A3(G264), .A4(new_n252), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n360), .A2(new_n362), .A3(G257), .A4(G1698), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n360), .A2(new_n362), .A3(G250), .A4(new_n257), .ZN(new_n545));
  INV_X1    g0345(.A(G294), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n544), .B(new_n545), .C1(new_n361), .C2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n542), .A2(new_n543), .B1(new_n247), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n305), .B1(new_n548), .B2(new_n444), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT83), .ZN(new_n550));
  AOI221_X4 g0350(.A(new_n445), .B1(new_n547), .B2(new_n247), .C1(new_n542), .C2(new_n543), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n549), .A2(new_n550), .B1(new_n551), .B2(G179), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT83), .B1(new_n551), .B2(new_n305), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n535), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT84), .B1(new_n551), .B2(G200), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n542), .A2(new_n543), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n547), .A2(new_n247), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n444), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT84), .ZN(new_n559));
  INV_X1    g0359(.A(G200), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n551), .A2(new_n402), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n555), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n554), .B1(new_n535), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n264), .A2(G116), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT80), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n431), .A2(G116), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n266), .A2(new_n216), .B1(G20), .B2(new_n476), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n449), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT20), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n569), .A2(KEYINPUT20), .A3(new_n570), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n567), .B(new_n568), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n255), .A2(G264), .A3(G1698), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n255), .A2(G257), .A3(new_n257), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n363), .A2(G303), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n247), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n247), .A2(new_n248), .ZN(new_n579));
  INV_X1    g0379(.A(new_n539), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n446), .A2(G270), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n573), .A2(new_n582), .A3(KEYINPUT21), .A4(G169), .ZN(new_n583));
  INV_X1    g0383(.A(G270), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n444), .B1(new_n540), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n247), .B2(new_n577), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(new_n573), .A3(G179), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n573), .B1(new_n582), .B2(G200), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n402), .B2(new_n582), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n573), .A2(new_n582), .A3(G169), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n588), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n428), .A2(new_n511), .A3(new_n564), .A4(new_n594), .ZN(G372));
  INV_X1    g0395(.A(new_n288), .ZN(new_n596));
  INV_X1    g0396(.A(new_n310), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n350), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n598), .A2(new_n346), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n389), .A2(new_n393), .A3(new_n408), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT17), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n410), .A2(KEYINPUT17), .A3(new_n408), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n427), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n596), .B1(new_n605), .B2(new_n285), .ZN(new_n606));
  INV_X1    g0406(.A(new_n535), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n558), .A2(new_n550), .A3(G169), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n548), .A2(G179), .A3(new_n444), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n549), .A2(new_n550), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n593), .A2(new_n587), .A3(new_n583), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n488), .A2(new_n498), .A3(new_n484), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n505), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n563), .B2(new_n535), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n614), .A2(new_n617), .A3(new_n473), .A4(new_n470), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n440), .A2(new_n469), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT26), .ZN(new_n620));
  INV_X1    g0420(.A(new_n616), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n472), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n615), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n506), .A2(new_n439), .A3(new_n472), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n624), .B2(KEYINPUT26), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n618), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n428), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n606), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g0428(.A(new_n628), .B(KEYINPUT85), .Z(G369));
  INV_X1    g0429(.A(KEYINPUT86), .ZN(new_n630));
  INV_X1    g0430(.A(new_n594), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n573), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n630), .B1(new_n631), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n588), .A2(new_n593), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n638), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n630), .A3(new_n638), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT87), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT87), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G330), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n637), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n564), .B1(new_n535), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n612), .B2(new_n650), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n613), .A2(new_n637), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n564), .A2(new_n654), .B1(new_n554), .B2(new_n650), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(G399));
  INV_X1    g0456(.A(new_n213), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(G41), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G1), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n219), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT28), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT30), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n447), .B1(new_n456), .B2(new_n461), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n586), .A2(new_n548), .A3(G179), .A4(new_n499), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT89), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT89), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n669), .B(new_n664), .C1(new_n665), .C2(new_n666), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n556), .A2(new_n499), .A3(new_n557), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n578), .A2(new_n581), .A3(G179), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n466), .A2(new_n673), .A3(KEYINPUT30), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n586), .A2(G179), .A3(new_n499), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n665), .A2(new_n675), .A3(new_n558), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n668), .A2(new_n670), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n637), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT31), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n667), .A2(new_n674), .A3(new_n676), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT88), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT88), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n563), .A2(new_n535), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n594), .A2(new_n686), .A3(new_n612), .A4(new_n650), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n508), .B2(new_n510), .ZN(new_n688));
  OAI21_X1  g0488(.A(G330), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT29), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n619), .A2(new_n472), .A3(new_n621), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT26), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n506), .A2(new_n620), .A3(new_n472), .A4(new_n439), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n615), .B(KEYINPUT90), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT91), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n554), .B2(new_n640), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n612), .A2(KEYINPUT91), .A3(new_n613), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n617), .A2(new_n473), .A3(new_n470), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n693), .B(new_n696), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n691), .B1(new_n702), .B2(new_n650), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n626), .A2(new_n691), .A3(new_n650), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n690), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n663), .B1(new_n705), .B2(G1), .ZN(G364));
  INV_X1    g0506(.A(G13), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G20), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n209), .B1(new_n708), .B2(G45), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n658), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n649), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n647), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G13), .A2(G33), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G20), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n711), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n657), .A2(new_n363), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n722), .A2(G355), .B1(new_n476), .B2(new_n657), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n657), .A2(new_n255), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(G45), .B2(new_n219), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n245), .A2(new_n442), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n216), .B1(G20), .B2(new_n305), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n718), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n721), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  XOR2_X1   g0530(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n210), .A2(G179), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n402), .A3(new_n560), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n732), .B1(new_n735), .B2(G159), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n732), .A2(new_n735), .A3(G159), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n733), .A2(G190), .A3(G200), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT95), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G87), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n210), .A2(new_n286), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n402), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(KEYINPUT92), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n747), .A2(KEYINPUT92), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n736), .B(new_n744), .C1(G58), .C2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n733), .A2(new_n402), .A3(G200), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n745), .A2(new_n402), .A3(new_n560), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n255), .B1(new_n754), .B2(new_n206), .C1(new_n221), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n746), .A2(new_n286), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n745), .A2(new_n402), .A3(G200), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n759), .A2(new_n205), .B1(new_n760), .B2(new_n354), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n745), .A2(G190), .A3(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT93), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n762), .A2(KEYINPUT93), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n756), .B(new_n761), .C1(new_n767), .C2(G50), .ZN(new_n768));
  INV_X1    g0568(.A(G329), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n363), .B1(new_n734), .B2(new_n769), .C1(new_n770), .C2(new_n755), .ZN(new_n771));
  INV_X1    g0571(.A(G303), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n742), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n771), .B(new_n773), .C1(G322), .C2(new_n752), .ZN(new_n774));
  INV_X1    g0574(.A(new_n760), .ZN(new_n775));
  NOR2_X1   g0575(.A1(KEYINPUT33), .A2(G317), .ZN(new_n776));
  AND2_X1   g0576(.A1(KEYINPUT33), .A2(G317), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G283), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n778), .B1(new_n779), .B2(new_n754), .C1(new_n546), .C2(new_n759), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT96), .B(G326), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(new_n767), .B2(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n753), .A2(new_n768), .B1(new_n774), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n728), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n730), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n713), .A2(new_n715), .B1(new_n720), .B2(new_n786), .ZN(G396));
  NAND2_X1  g0587(.A1(new_n297), .A2(new_n637), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n313), .A2(new_n310), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT99), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(KEYINPUT99), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n626), .A2(new_n792), .A3(new_n650), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n626), .A2(new_n650), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n790), .B(new_n791), .C1(new_n310), .C2(new_n650), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n721), .B1(new_n796), .B2(new_n689), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n689), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(KEYINPUT100), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(KEYINPUT100), .B2(new_n798), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n728), .A2(new_n716), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT97), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n711), .B1(new_n802), .B2(G77), .ZN(new_n803));
  INV_X1    g0603(.A(new_n755), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G150), .A2(new_n775), .B1(new_n804), .B2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G143), .ZN(new_n806));
  INV_X1    g0606(.A(G137), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(new_n751), .B2(new_n806), .C1(new_n807), .C2(new_n766), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT34), .Z(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n759), .A2(new_n353), .B1(new_n734), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n255), .B1(new_n754), .B2(new_n354), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n202), .B2(new_n742), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n759), .A2(new_n205), .B1(new_n755), .B2(new_n476), .ZN(new_n815));
  INV_X1    g0615(.A(new_n754), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G283), .A2(new_n775), .B1(new_n816), .B2(G87), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n770), .B2(new_n734), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n815), .B(new_n818), .C1(G294), .C2(new_n752), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n772), .B2(new_n766), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n363), .B1(new_n742), .B2(new_n206), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT98), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n809), .A2(new_n814), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n803), .B1(new_n823), .B2(new_n728), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n795), .B2(new_n717), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n800), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G384));
  INV_X1    g0627(.A(new_n436), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n828), .A2(KEYINPUT35), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(KEYINPUT35), .ZN(new_n830));
  NOR4_X1   g0630(.A1(new_n829), .A2(new_n830), .A3(new_n476), .A4(new_n218), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT36), .ZN(new_n832));
  OR3_X1    g0632(.A1(new_n355), .A2(new_n219), .A3(new_n221), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n202), .A2(G68), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n209), .B(G13), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n351), .B1(new_n326), .B2(new_n637), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n326), .A2(new_n637), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n346), .B2(new_n350), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n310), .A2(new_n637), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n793), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n370), .B1(KEYINPUT16), .B2(new_n369), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n393), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n635), .B(new_n848), .C1(new_n412), .C2(new_n427), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n422), .A2(new_n635), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n847), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n600), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n420), .A2(new_n850), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n600), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(KEYINPUT37), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n845), .B1(new_n849), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n635), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n424), .A2(new_n426), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n859), .B(new_n847), .C1(new_n860), .C2(new_n604), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n856), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n844), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n860), .B2(new_n635), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT39), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n856), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n420), .B(new_n859), .C1(new_n860), .C2(new_n604), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n854), .A2(KEYINPUT101), .A3(KEYINPUT37), .A4(new_n600), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT101), .ZN(new_n870));
  INV_X1    g0670(.A(new_n850), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n410), .B2(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .B1(new_n854), .B2(new_n600), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n867), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n865), .B1(new_n866), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n858), .A2(KEYINPUT39), .A3(new_n862), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n346), .A2(new_n637), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n864), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n428), .B1(new_n703), .B2(new_n704), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n606), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n880), .B(new_n882), .Z(new_n883));
  OAI21_X1  g0683(.A(new_n795), .B1(new_n837), .B2(new_n839), .ZN(new_n884));
  INV_X1    g0684(.A(new_n687), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n511), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(KEYINPUT102), .A3(new_n680), .A4(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n680), .A2(new_n887), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n889), .B1(new_n890), .B2(new_n688), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n884), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n866), .B2(new_n875), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT40), .B1(new_n858), .B2(new_n862), .ZN(new_n894));
  AOI22_X1  g0694(.A1(KEYINPUT40), .A2(new_n893), .B1(new_n894), .B2(new_n892), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n352), .A2(new_n412), .A3(new_n427), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n888), .B2(new_n891), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n648), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n898), .B2(new_n896), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n883), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n708), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(G1), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT103), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n883), .A2(new_n900), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n836), .B1(new_n906), .B2(new_n908), .ZN(G367));
  NAND2_X1  g0709(.A1(new_n619), .A2(new_n637), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n473), .A3(new_n470), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n619), .A2(new_n472), .A3(new_n637), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n564), .A2(new_n654), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT42), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n473), .B1(new_n914), .B2(new_n612), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n650), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n503), .A2(new_n650), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n615), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n621), .B2(new_n921), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT104), .Z(new_n924));
  INV_X1    g0724(.A(KEYINPUT43), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n917), .A2(new_n925), .A3(new_n924), .A4(new_n919), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n927), .B1(KEYINPUT105), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(KEYINPUT105), .B2(new_n928), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n653), .A2(new_n914), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n658), .B(KEYINPUT41), .Z(new_n933));
  NAND2_X1  g0733(.A1(new_n655), .A2(new_n913), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT106), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT45), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n655), .A2(new_n913), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT44), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(new_n653), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n915), .B1(new_n652), .B2(new_n654), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n649), .B(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n705), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n933), .B1(new_n945), .B2(new_n705), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n932), .B1(new_n946), .B2(new_n710), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n924), .A2(new_n718), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n724), .A2(new_n237), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n213), .A2(new_n291), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n950), .A2(new_n718), .A3(new_n728), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n721), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n751), .A2(new_n772), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n754), .A2(new_n205), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n759), .A2(new_n206), .B1(new_n760), .B2(new_n546), .ZN(new_n955));
  XOR2_X1   g0755(.A(KEYINPUT107), .B(G317), .Z(new_n956));
  OAI221_X1 g0756(.A(new_n363), .B1(new_n755), .B2(new_n779), .C1(new_n734), .C2(new_n956), .ZN(new_n957));
  NOR4_X1   g0757(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT46), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n742), .B2(new_n476), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n767), .A2(G311), .ZN(new_n961));
  INV_X1    g0761(.A(new_n742), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(KEYINPUT46), .A3(G116), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n958), .A2(new_n960), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT108), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT109), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n255), .B1(new_n754), .B2(new_n221), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n767), .A2(G143), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G150), .A2(new_n752), .B1(new_n962), .B2(G58), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n759), .A2(new_n354), .B1(new_n760), .B2(new_n357), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n755), .A2(new_n202), .B1(new_n734), .B2(new_n807), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n967), .A2(new_n966), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n968), .A2(new_n969), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n965), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT110), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT47), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n948), .B(new_n952), .C1(new_n977), .C2(new_n785), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT111), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n947), .A2(new_n979), .ZN(G387));
  OR2_X1    g0780(.A1(new_n652), .A2(new_n719), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n289), .A2(new_n202), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT50), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n660), .B(new_n442), .C1(new_n354), .C2(new_n221), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n724), .B1(new_n983), .B2(new_n984), .C1(new_n234), .C2(new_n442), .ZN(new_n985));
  INV_X1    g0785(.A(new_n660), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n722), .A2(new_n986), .B1(new_n206), .B2(new_n657), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n985), .A2(KEYINPUT112), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n729), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT112), .B1(new_n985), .B2(new_n987), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n711), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n759), .A2(new_n291), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n760), .A2(new_n271), .B1(new_n734), .B2(new_n273), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n767), .C2(G159), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n752), .A2(G50), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n962), .A2(G77), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n363), .B(new_n954), .C1(G68), .C2(new_n804), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT113), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n255), .B1(new_n816), .B2(G116), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n742), .A2(new_n546), .B1(new_n779), .B2(new_n759), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT114), .Z(new_n1002));
  INV_X1    g0802(.A(KEYINPUT48), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G303), .A2(new_n804), .B1(new_n775), .B2(G311), .ZN(new_n1004));
  INV_X1    g0804(.A(G322), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1004), .B1(new_n751), .B2(new_n956), .C1(new_n766), .C2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1002), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1000), .B1(new_n734), .B2(new_n781), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n999), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n991), .B1(new_n1012), .B2(new_n728), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n944), .A2(new_n710), .B1(new_n981), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n944), .A2(new_n705), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n658), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n944), .A2(new_n705), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT115), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(G393));
  NAND2_X1  g0822(.A1(new_n942), .A2(new_n710), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n767), .A2(G317), .B1(new_n752), .B2(G311), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT52), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n363), .B1(new_n755), .B2(new_n546), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G107), .B2(new_n816), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n1005), .B2(new_n734), .C1(new_n779), .C2(new_n742), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G303), .A2(new_n775), .B1(new_n758), .B2(G116), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT116), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1025), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n766), .A2(new_n273), .B1(new_n751), .B2(new_n357), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT51), .Z(new_n1033));
  NAND2_X1  g0833(.A1(new_n758), .A2(G77), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n806), .B2(new_n734), .C1(new_n202), .C2(new_n760), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n363), .B1(new_n804), .B2(new_n289), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n743), .B2(new_n754), .C1(new_n742), .C2(new_n354), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1033), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n728), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n729), .B1(new_n205), .B2(new_n213), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n242), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1040), .B1(new_n1041), .B2(new_n724), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(new_n721), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1039), .B(new_n1043), .C1(new_n913), .C2(new_n719), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n945), .A2(new_n658), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n942), .B1(new_n705), .B2(new_n944), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1023), .B(new_n1044), .C1(new_n1045), .C2(new_n1046), .ZN(G390));
  AOI21_X1  g0847(.A(new_n878), .B1(new_n840), .B2(new_n843), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT38), .B1(new_n861), .B2(new_n856), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n866), .A2(new_n1050), .A3(new_n865), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n410), .B(new_n635), .C1(new_n412), .C2(new_n427), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n873), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n868), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n845), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT39), .B1(new_n1055), .B2(new_n862), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1049), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(G330), .B(new_n795), .C1(new_n685), .C2(new_n688), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n837), .A2(new_n839), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1055), .A2(new_n862), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n702), .A2(new_n650), .A3(new_n792), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n842), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n878), .B1(new_n1063), .B2(new_n840), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1057), .A2(new_n1060), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n648), .B1(new_n888), .B2(new_n891), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n884), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1048), .B1(new_n876), .B2(new_n877), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1066), .A2(new_n1073), .A3(new_n710), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n716), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n711), .B1(new_n802), .B2(new_n289), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1034), .B1(new_n546), .B2(new_n734), .C1(new_n206), .C2(new_n760), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G283), .B2(new_n767), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n363), .B1(new_n754), .B2(new_n354), .C1(new_n205), .C2(new_n755), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n962), .B2(G87), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(new_n476), .C2(new_n751), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n742), .A2(new_n273), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT53), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n767), .A2(G128), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n759), .A2(new_n357), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT54), .B(G143), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n807), .A2(new_n760), .B1(new_n755), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1085), .B(new_n1087), .C1(new_n752), .C2(G132), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1083), .A2(new_n1084), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(G125), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n255), .B1(new_n734), .B2(new_n1090), .C1(new_n202), .C2(new_n754), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT118), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1081), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1076), .B1(new_n1093), .B2(new_n728), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1075), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1074), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT119), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT119), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1074), .A2(new_n1098), .A3(new_n1095), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1066), .A2(new_n1073), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n888), .A2(new_n891), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(G330), .A3(new_n428), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT117), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n606), .A4(new_n881), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n648), .B(new_n897), .C1(new_n888), .C2(new_n891), .ZN(new_n1107));
  OAI21_X1  g0907(.A(KEYINPUT117), .B1(new_n1107), .B2(new_n882), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1069), .A2(new_n1109), .B1(new_n793), .B2(new_n842), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n842), .B(new_n1062), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1067), .A2(new_n795), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n1059), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1106), .B(new_n1108), .C1(new_n1110), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n659), .B1(new_n1102), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1101), .A2(new_n1114), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1100), .A2(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(KEYINPUT123), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1108), .A2(new_n1106), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n1108), .B2(new_n1106), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1101), .B2(new_n1114), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n285), .A2(new_n288), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n279), .A2(new_n859), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1125), .B(new_n1126), .Z(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1127), .B(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n895), .B2(new_n648), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1129), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT40), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n892), .B(new_n1132), .C1(new_n866), .C2(new_n1050), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1132), .B1(new_n1061), .B2(new_n892), .ZN(new_n1135));
  OAI211_X1 g0935(.A(G330), .B(new_n1131), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1130), .A2(new_n880), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n880), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1124), .B(KEYINPUT57), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n658), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1130), .A2(new_n1136), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n880), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1130), .A2(new_n880), .A3(new_n1136), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT57), .B1(new_n1145), .B2(new_n1124), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n710), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n721), .B1(new_n202), .B2(new_n801), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n760), .A2(new_n810), .B1(new_n755), .B2(new_n807), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n752), .A2(G128), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1086), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n962), .A2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1150), .B(new_n1151), .C1(KEYINPUT121), .C2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(KEYINPUT121), .B2(new_n1153), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n766), .A2(new_n1090), .B1(new_n273), .B2(new_n759), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT122), .Z(new_n1157));
  NOR2_X1   g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n735), .A2(G124), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G33), .B(G41), .C1(new_n816), .C2(G159), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n255), .A2(G41), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n291), .B2(new_n755), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G68), .B2(new_n758), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n996), .B(new_n1167), .C1(new_n206), .C2(new_n751), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n766), .A2(new_n476), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n754), .A2(new_n353), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n760), .A2(new_n205), .B1(new_n734), .B2(new_n779), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT120), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT58), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1173), .A2(KEYINPUT58), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1165), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1176), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1177));
  AND4_X1   g0977(.A1(new_n1164), .A2(new_n1174), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1149), .B1(new_n785), .B2(new_n1178), .C1(new_n1131), .C2(new_n717), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1148), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1147), .A2(new_n1180), .ZN(G375));
  NOR2_X1   g0981(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT124), .B1(new_n1183), .B2(new_n710), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(KEYINPUT124), .A3(new_n710), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1059), .A2(new_n716), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n711), .B1(new_n802), .B2(G68), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n992), .B1(G116), .B2(new_n775), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n772), .B2(new_n734), .C1(new_n766), .C2(new_n546), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n363), .B1(new_n755), .B2(new_n206), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G77), .B2(new_n816), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n742), .B2(new_n205), .C1(new_n779), .C2(new_n751), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n363), .B(new_n1170), .C1(G150), .C2(new_n804), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n807), .B2(new_n751), .C1(new_n357), .C2(new_n742), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n735), .A2(G128), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n775), .A2(new_n1152), .B1(new_n758), .B2(G50), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n766), .C2(new_n810), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n1190), .A2(new_n1193), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1188), .B1(new_n1199), .B2(new_n728), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1184), .B(new_n1186), .C1(new_n1187), .C2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1108), .A2(new_n1106), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1182), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n933), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n1204), .A3(new_n1114), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n1205), .ZN(G381));
  AOI22_X1  g1006(.A1(new_n1097), .A2(new_n1099), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1147), .A2(new_n1207), .A3(new_n1180), .ZN(new_n1208));
  INV_X1    g1008(.A(G396), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1020), .A2(new_n1209), .A3(new_n1021), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(G390), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n826), .A3(new_n1212), .ZN(new_n1213));
  OR4_X1    g1013(.A1(G387), .A2(new_n1208), .A3(new_n1213), .A4(G381), .ZN(G407));
  OAI211_X1 g1014(.A(G407), .B(G213), .C1(G343), .C2(new_n1208), .ZN(G409));
  OAI211_X1 g1015(.A(new_n1124), .B(new_n1204), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n1148), .A3(new_n1179), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1207), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT125), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1180), .B(G378), .C1(new_n1140), .C2(new_n1146), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1217), .A2(new_n1207), .A3(KEYINPUT125), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n636), .A2(G213), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT127), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1114), .A2(KEYINPUT60), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1203), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n659), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1228), .B2(new_n1227), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1201), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(new_n826), .ZN(new_n1232));
  AOI21_X1  g1032(.A(G384), .B1(new_n1201), .B2(new_n1230), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT127), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1223), .A2(new_n1235), .A3(new_n1224), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1226), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT62), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT61), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1231), .B(new_n826), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT126), .B1(new_n1225), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT62), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT126), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1234), .A2(new_n1223), .A3(new_n1243), .A4(new_n1224), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n636), .A2(G213), .A3(G2897), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1240), .A2(new_n1246), .ZN(new_n1247));
  OR3_X1    g1047(.A1(new_n1232), .A2(new_n1233), .A3(new_n1246), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1236), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1235), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1238), .A2(new_n1239), .A3(new_n1245), .A4(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G393), .B(G396), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(G387), .A2(new_n1212), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G390), .B1(new_n947), .B2(new_n979), .ZN(new_n1256));
  OR3_X1    g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1253), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1257), .A2(new_n1239), .A3(new_n1258), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1225), .B2(new_n1249), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1262), .B(new_n1265), .C1(new_n1264), .C2(new_n1237), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1260), .A2(new_n1266), .ZN(G405));
  NAND2_X1  g1067(.A1(G375), .A2(new_n1207), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1221), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(new_n1240), .ZN(new_n1270));
  XOR2_X1   g1070(.A(new_n1270), .B(new_n1259), .Z(G402));
endmodule


