//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(G20), .A3(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT64), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT5), .B(G41), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  OAI211_X1 g0049(.A(G1), .B(G13), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G45), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n247), .A2(new_n250), .A3(G274), .A4(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(new_n252), .B2(new_n247), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n254), .B1(G270), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT75), .B1(new_n248), .B2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT75), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n225), .A2(G1698), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G257), .B2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G303), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n263), .A2(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n255), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n257), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT86), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT86), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n257), .A2(new_n272), .A3(new_n269), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G283), .ZN(new_n275));
  INV_X1    g0075(.A(G20), .ZN(new_n276));
  INV_X1    g0076(.A(G97), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n275), .B(new_n276), .C1(G33), .C2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n212), .B1(new_n206), .B2(new_n248), .ZN(new_n279));
  INV_X1    g0079(.A(G116), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G20), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT88), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n282), .A2(KEYINPUT88), .A3(new_n283), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT20), .A4(new_n281), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT87), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n289), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n286), .A2(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G13), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G1), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n293), .A2(new_n276), .A3(G1), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT69), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n279), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G1), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n280), .B1(new_n301), .B2(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n296), .A2(new_n299), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(G116), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(G169), .B1(new_n292), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n274), .A2(new_n307), .A3(KEYINPUT21), .ZN(new_n308));
  INV_X1    g0108(.A(new_n292), .ZN(new_n309));
  INV_X1    g0109(.A(new_n305), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n270), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT21), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n271), .A2(new_n273), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n306), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n311), .B1(new_n317), .B2(G190), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n317), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n315), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(G222), .A2(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(G1698), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(G223), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n267), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n326), .B(new_n255), .C1(G77), .C2(new_n267), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n301), .B1(G41), .B2(G45), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(new_n250), .A3(G274), .ZN(new_n330));
  INV_X1    g0130(.A(G226), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n250), .A2(new_n328), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n327), .B(new_n330), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n333), .B(KEYINPUT65), .Z(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G200), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n276), .A2(G1), .ZN(new_n336));
  OR3_X1    g0136(.A1(new_n336), .A2(KEYINPUT66), .A3(new_n202), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n297), .A2(new_n279), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT66), .B1(new_n336), .B2(new_n202), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n276), .B1(new_n201), .B2(new_n202), .ZN(new_n341));
  NOR2_X1   g0141(.A1(G20), .A2(G33), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G150), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n276), .A2(G33), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  XOR2_X1   g0147(.A(KEYINPUT8), .B(G58), .Z(new_n348));
  AOI211_X1 g0148(.A(new_n341), .B(new_n345), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n279), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n340), .B1(G50), .B2(new_n295), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT9), .ZN(new_n352));
  INV_X1    g0152(.A(G190), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n335), .B(new_n352), .C1(new_n353), .C2(new_n334), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT10), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n334), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n351), .C1(G179), .C2(new_n334), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n231), .A2(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n267), .B(new_n360), .C1(G226), .C2(G1698), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n255), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n330), .B1(new_n332), .B2(new_n217), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n250), .B1(new_n361), .B2(new_n362), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT13), .B1(new_n369), .B2(new_n365), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n320), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n216), .A2(G20), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n373), .B1(new_n346), .B2(new_n222), .C1(new_n343), .C2(new_n202), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT73), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(new_n279), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n375), .B1(new_n374), .B2(new_n279), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT11), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT12), .B1(new_n304), .B2(G68), .ZN(new_n380));
  OR4_X1    g0180(.A1(KEYINPUT12), .A2(new_n373), .A3(G1), .A4(new_n293), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n336), .A2(new_n216), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n380), .A2(new_n381), .B1(new_n300), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n378), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT11), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n376), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n379), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n368), .A2(KEYINPUT72), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT72), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n364), .A2(new_n366), .A3(new_n389), .A4(new_n367), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n370), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n387), .B1(new_n391), .B2(new_n353), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n372), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n356), .B1(new_n368), .B2(new_n370), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT14), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n390), .A2(new_n370), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n369), .A2(new_n365), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n389), .B1(new_n397), .B2(new_n367), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT74), .B1(new_n399), .B2(G179), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n388), .A2(G179), .A3(new_n370), .A4(new_n390), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT74), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n395), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n387), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n393), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n330), .B1(new_n332), .B2(new_n223), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n267), .A2(G238), .A3(G1698), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n267), .A2(G232), .A3(new_n324), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n408), .B(new_n409), .C1(new_n224), .C2(new_n267), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n410), .A2(KEYINPUT67), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n250), .B1(new_n410), .B2(KEYINPUT67), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n312), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT70), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(KEYINPUT70), .A3(new_n312), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT15), .B(G87), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n347), .B1(G20), .B2(G77), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT68), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n348), .B(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n423), .B2(new_n343), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n279), .ZN(new_n425));
  INV_X1    g0225(.A(new_n304), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n336), .A2(new_n222), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n426), .A2(new_n222), .B1(new_n300), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n413), .B2(G169), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n418), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n413), .A2(G190), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n433), .B(new_n434), .C1(new_n320), .C2(new_n413), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n359), .A2(new_n406), .A3(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n338), .B(new_n348), .C1(G1), .C2(new_n276), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n295), .B2(new_n348), .ZN(new_n439));
  XOR2_X1   g0239(.A(new_n439), .B(KEYINPUT79), .Z(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(G58), .A2(G68), .ZN(new_n442));
  OAI21_X1  g0242(.A(G20), .B1(new_n442), .B2(new_n201), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n342), .A2(G159), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(G20), .C1(new_n442), .C2(new_n201), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n263), .A2(new_n276), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n216), .B1(new_n449), .B2(KEYINPUT7), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT7), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n263), .A2(new_n451), .A3(new_n276), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n448), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT16), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n260), .A2(G33), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n262), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT7), .B1(new_n456), .B2(new_n276), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n451), .B(G20), .C1(new_n455), .C2(new_n262), .ZN(new_n458));
  OAI21_X1  g0258(.A(G68), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT16), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT77), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n451), .B1(new_n267), .B2(G20), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n260), .A2(G33), .ZN(new_n466));
  OAI211_X1 g0266(.A(KEYINPUT7), .B(new_n276), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n216), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(KEYINPUT77), .B(new_n462), .C1(new_n468), .C2(new_n448), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n279), .B(new_n454), .C1(new_n463), .C2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT78), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n462), .B1(new_n468), .B2(new_n448), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT77), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n350), .B1(new_n476), .B2(new_n469), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(KEYINPUT78), .A3(new_n454), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n441), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n330), .B1(new_n332), .B2(new_n231), .ZN(new_n480));
  XOR2_X1   g0280(.A(new_n480), .B(KEYINPUT80), .Z(new_n481));
  OR2_X1    g0281(.A1(G223), .A2(G1698), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(G226), .B2(new_n324), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n263), .A2(new_n483), .B1(new_n248), .B2(new_n218), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n255), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n312), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n480), .B1(new_n255), .B2(new_n484), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n481), .A2(new_n486), .B1(G169), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT18), .B1(new_n479), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n476), .A2(new_n469), .ZN(new_n490));
  AND4_X1   g0290(.A1(KEYINPUT78), .A2(new_n490), .A3(new_n279), .A4(new_n454), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT78), .B1(new_n477), .B2(new_n454), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n440), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT18), .ZN(new_n494));
  INV_X1    g0294(.A(new_n488), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n485), .A2(new_n353), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n481), .A2(new_n498), .B1(G200), .B2(new_n487), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n440), .B(new_n499), .C1(new_n491), .C2(new_n492), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT17), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT17), .B1(new_n479), .B2(new_n499), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n437), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(G250), .A2(G1698), .ZN(new_n507));
  INV_X1    g0307(.A(G257), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(G1698), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n509), .A2(new_n262), .A3(new_n258), .A4(new_n261), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n250), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  NOR2_X1   g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n252), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n515), .A2(G264), .A3(new_n250), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT89), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n508), .A2(G1698), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(G250), .B2(G1698), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n511), .B1(new_n263), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n255), .ZN(new_n521));
  INV_X1    g0321(.A(new_n516), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT89), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n517), .A2(new_n524), .A3(new_n253), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n320), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n512), .A2(new_n254), .A3(new_n516), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n353), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n267), .A2(new_n276), .A3(G87), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT22), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n276), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n224), .A2(KEYINPUT23), .A3(G20), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n276), .A2(G33), .A3(G116), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n532), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n258), .A2(new_n261), .A3(new_n276), .A4(new_n262), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n541), .A2(new_n531), .A3(new_n218), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT24), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n538), .B1(new_n531), .B2(new_n530), .ZN(new_n544));
  INV_X1    g0344(.A(new_n263), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n545), .A2(KEYINPUT22), .A3(new_n276), .A4(G87), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n350), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n338), .B1(G1), .B2(new_n248), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n224), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n297), .A2(new_n224), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT25), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n529), .A2(new_n554), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n525), .A2(new_n312), .B1(new_n527), .B2(new_n356), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n540), .A2(new_n542), .A3(KEYINPUT24), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n547), .B1(new_n544), .B2(new_n546), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n279), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n551), .A2(new_n553), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n455), .A2(new_n262), .A3(G250), .A4(G1698), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n275), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT4), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n223), .A2(G1698), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n258), .A2(new_n261), .A3(new_n262), .A4(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(KEYINPUT4), .A2(G244), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n455), .A2(new_n262), .A3(new_n570), .A4(new_n324), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT82), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT82), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n267), .A2(new_n573), .A3(new_n324), .A4(new_n570), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n250), .B1(new_n569), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n515), .A2(G257), .A3(new_n250), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n253), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT83), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n253), .A3(KEYINPUT83), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(G200), .B1(new_n576), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n568), .A2(new_n566), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n575), .A2(new_n275), .A3(new_n584), .A4(new_n564), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n255), .ZN(new_n586));
  INV_X1    g0386(.A(new_n578), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(G190), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n295), .A2(G97), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n550), .B2(new_n277), .ZN(new_n591));
  OAI21_X1  g0391(.A(G107), .B1(new_n457), .B2(new_n458), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n342), .A2(G77), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT6), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n594), .A2(G97), .A3(G107), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n277), .A2(KEYINPUT6), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n224), .A2(KEYINPUT81), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n224), .A2(KEYINPUT81), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n595), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g0399(.A(KEYINPUT81), .B(G107), .ZN(new_n600));
  INV_X1    g0400(.A(new_n596), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n277), .A2(new_n224), .A3(KEYINPUT6), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(new_n603), .A3(G20), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n592), .A2(new_n593), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n591), .B1(new_n605), .B2(new_n279), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n583), .A2(new_n588), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n356), .B1(new_n576), .B2(new_n578), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n577), .A2(new_n253), .A3(KEYINPUT83), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT83), .B1(new_n577), .B2(new_n253), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n586), .A2(new_n312), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n604), .A2(new_n593), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n224), .B1(new_n464), .B2(new_n467), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n279), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n591), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n608), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n607), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n252), .A2(new_n219), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n250), .ZN(new_n621));
  INV_X1    g0421(.A(new_n252), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n250), .A2(G274), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n223), .A2(G1698), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(G238), .B2(G1698), .ZN(new_n626));
  OAI22_X1  g0426(.A1(new_n263), .A2(new_n626), .B1(new_n248), .B2(new_n280), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n624), .B1(new_n255), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT85), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(G190), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n255), .ZN(new_n631));
  INV_X1    g0431(.A(G274), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n255), .A2(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n633), .A2(new_n252), .B1(new_n250), .B2(new_n620), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(G190), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT85), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT19), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n346), .B2(new_n277), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n541), .B2(new_n216), .ZN(new_n641));
  NAND3_X1  g0441(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT84), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n643), .A3(new_n276), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n218), .A2(new_n277), .A3(new_n224), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n642), .B2(new_n276), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n279), .B1(new_n641), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n426), .A2(new_n419), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n338), .B(G87), .C1(G1), .C2(new_n248), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n631), .A2(new_n634), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(G200), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n628), .A2(new_n312), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n356), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n649), .B(new_n650), .C1(new_n550), .C2(new_n419), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n638), .A2(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n619), .A2(new_n659), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n322), .A2(new_n506), .A3(new_n563), .A4(new_n660), .ZN(G372));
  AOI22_X1  g0461(.A1(new_n525), .A2(new_n320), .B1(new_n527), .B2(new_n353), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n618), .B(new_n607), .C1(new_n662), .C2(new_n561), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n649), .A2(new_n650), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n653), .A2(G200), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(new_n651), .A4(new_n635), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n658), .A2(new_n655), .A3(new_n656), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT90), .B1(new_n663), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  INV_X1    g0470(.A(new_n668), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n619), .A2(new_n670), .A3(new_n555), .A4(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n308), .A2(new_n562), .A3(new_n318), .A4(new_n314), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n667), .B(KEYINPUT91), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n664), .A2(new_n665), .A3(new_n651), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n667), .B1(new_n677), .B2(new_n637), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT26), .B1(new_n678), .B2(new_n618), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  INV_X1    g0480(.A(new_n618), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n671), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n676), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n506), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g0485(.A(new_n685), .B(KEYINPUT92), .Z(new_n686));
  NAND2_X1  g0486(.A1(new_n500), .A2(new_n501), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n479), .A2(KEYINPUT17), .A3(new_n499), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n404), .A2(new_n405), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n372), .A2(new_n392), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n430), .B1(new_n416), .B2(new_n417), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n689), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n489), .A2(new_n496), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n355), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(new_n358), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n686), .A2(new_n697), .ZN(G369));
  NAND2_X1  g0498(.A1(new_n315), .A2(new_n318), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n294), .A2(new_n276), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n311), .A2(new_n705), .ZN(new_n706));
  MUX2_X1   g0506(.A(new_n699), .B(new_n322), .S(new_n706), .Z(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n705), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n563), .B1(new_n554), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n562), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n562), .A2(new_n705), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n705), .B1(new_n315), .B2(new_n318), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n563), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(new_n716), .ZN(G399));
  NOR2_X1   g0517(.A1(new_n645), .A2(G116), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n207), .A2(new_n249), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(G1), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n210), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n313), .A2(new_n586), .A3(new_n587), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n517), .A2(new_n524), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n628), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT93), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(KEYINPUT93), .A3(new_n628), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n586), .A2(new_n611), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n628), .A2(G179), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n274), .A2(new_n525), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n729), .B2(KEYINPUT30), .ZN(new_n734));
  OAI211_X1 g0534(.A(KEYINPUT31), .B(new_n705), .C1(new_n730), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(KEYINPUT94), .ZN(new_n736));
  INV_X1    g0536(.A(G330), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n705), .B1(new_n730), .B2(new_n734), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n322), .A2(new_n563), .A3(new_n660), .A4(new_n710), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(KEYINPUT94), .A3(new_n742), .A4(new_n735), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n659), .A2(new_n680), .A3(new_n681), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT95), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT26), .B1(new_n668), .B2(new_n618), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n745), .A2(new_n676), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n673), .A2(new_n555), .A3(new_n619), .A4(new_n671), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n678), .A2(new_n618), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n675), .B1(new_n751), .B2(new_n680), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n746), .B1(new_n752), .B2(new_n747), .ZN(new_n753));
  OAI211_X1 g0553(.A(KEYINPUT29), .B(new_n710), .C1(new_n750), .C2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n705), .B1(new_n674), .B2(new_n683), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n754), .B1(KEYINPUT29), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n744), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT96), .Z(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n722), .B1(new_n759), .B2(G1), .ZN(G364));
  NOR2_X1   g0560(.A1(new_n293), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n301), .B1(new_n761), .B2(G45), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n719), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT97), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n709), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G330), .B2(new_n707), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n267), .A2(new_n207), .ZN(new_n768));
  INV_X1    g0568(.A(G355), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n768), .A2(new_n769), .B1(G116), .B2(new_n207), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n245), .A2(new_n251), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n263), .A2(new_n207), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n251), .B2(new_n211), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n213), .B1(new_n276), .B2(G169), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT98), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT98), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n765), .B1(new_n774), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n276), .A2(G179), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(new_n353), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n224), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n276), .A2(new_n312), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n353), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n785), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G159), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n791), .A2(new_n202), .B1(new_n795), .B2(KEYINPUT32), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n787), .B(new_n796), .C1(KEYINPUT32), .C2(new_n795), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n789), .A2(G190), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n353), .A2(G179), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n276), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n799), .A2(new_n216), .B1(new_n277), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT100), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n218), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n788), .A2(new_n792), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n267), .B1(new_n806), .B2(new_n222), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n788), .A2(G190), .A3(new_n320), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT99), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n805), .B(new_n807), .C1(new_n809), .C2(G58), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n797), .A2(new_n803), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  INV_X1    g0612(.A(G329), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n806), .A2(new_n812), .B1(new_n793), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n808), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n267), .B(new_n814), .C1(G322), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G317), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n798), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n801), .ZN(new_n821));
  INV_X1    g0621(.A(new_n804), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n821), .A2(G294), .B1(new_n822), .B2(G303), .ZN(new_n823));
  INV_X1    g0623(.A(new_n786), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n790), .A2(G326), .B1(new_n824), .B2(G283), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n816), .A2(new_n820), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n811), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n784), .B1(new_n827), .B2(new_n778), .ZN(new_n828));
  INV_X1    g0628(.A(new_n781), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n707), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n767), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  NOR2_X1   g0632(.A1(new_n433), .A2(new_n710), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n692), .A2(new_n834), .A3(KEYINPUT104), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT104), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n432), .A2(new_n836), .A3(new_n435), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n835), .B1(new_n837), .B2(new_n834), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT105), .ZN(new_n839));
  MUX2_X1   g0639(.A(new_n839), .B(new_n838), .S(new_n755), .Z(new_n840));
  AOI21_X1  g0640(.A(new_n765), .B1(new_n840), .B2(new_n744), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n744), .B2(new_n840), .ZN(new_n842));
  INV_X1    g0642(.A(new_n778), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n780), .ZN(new_n844));
  INV_X1    g0644(.A(new_n806), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G116), .A2(new_n845), .B1(new_n794), .B2(G311), .ZN(new_n846));
  INV_X1    g0646(.A(G294), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n846), .B(new_n456), .C1(new_n847), .C2(new_n808), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n791), .A2(new_n266), .B1(new_n804), .B2(new_n224), .ZN(new_n849));
  INV_X1    g0649(.A(G283), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n799), .A2(new_n850), .B1(new_n277), .B2(new_n801), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n786), .A2(new_n218), .ZN(new_n852));
  NOR4_X1   g0652(.A1(new_n848), .A2(new_n849), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n790), .A2(G137), .B1(new_n845), .B2(G159), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n344), .B2(new_n799), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G143), .B2(new_n809), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT34), .Z(new_n857));
  OAI22_X1  g0657(.A1(new_n202), .A2(new_n804), .B1(new_n786), .B2(new_n216), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n858), .A2(KEYINPUT101), .B1(G58), .B2(new_n821), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(KEYINPUT101), .B2(new_n858), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n263), .B1(new_n794), .B2(G132), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT102), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n853), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n765), .B1(G77), .B2(new_n844), .C1(new_n864), .C2(new_n843), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT103), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n780), .B2(new_n838), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n842), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(G384));
  NOR3_X1   g0669(.A1(new_n212), .A2(new_n276), .A3(new_n280), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n599), .A2(new_n603), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT35), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n872), .B2(new_n871), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT36), .ZN(new_n875));
  INV_X1    g0675(.A(G58), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n211), .B(G77), .C1(new_n876), .C2(new_n216), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n202), .A2(G68), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n301), .B(G13), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n761), .A2(new_n301), .ZN(new_n881));
  INV_X1    g0681(.A(new_n703), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n497), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n684), .A2(new_n838), .A3(new_n710), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n692), .A2(new_n710), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n405), .A2(new_n705), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n368), .A2(new_n370), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(G169), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT14), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT14), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n394), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n401), .A2(new_n402), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n399), .A2(KEYINPUT74), .A3(G179), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n691), .B(new_n887), .C1(new_n896), .C2(new_n387), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n405), .B(new_n705), .C1(new_n404), .C2(new_n393), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT106), .B1(new_n886), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT106), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n902), .B(new_n899), .C1(new_n884), .C2(new_n885), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT108), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n462), .B1(new_n453), .B2(KEYINPUT107), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT107), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n907), .B(new_n448), .C1(new_n450), .C2(new_n452), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n905), .B(new_n279), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n454), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n449), .A2(KEYINPUT7), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(G68), .A3(new_n452), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n460), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n907), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n453), .A2(KEYINPUT107), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n462), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n905), .B1(new_n916), .B2(new_n279), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n440), .B1(new_n910), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n918), .A2(KEYINPUT109), .A3(new_n882), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT109), .B1(new_n918), .B2(new_n882), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n695), .A2(new_n689), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT37), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n919), .A2(new_n920), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n918), .A2(new_n495), .B1(new_n479), .B2(new_n499), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n500), .B1(new_n479), .B2(new_n488), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n479), .A2(new_n703), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n926), .A2(KEYINPUT37), .A3(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(KEYINPUT38), .B(new_n921), .C1(new_n925), .C2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT38), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT109), .ZN(new_n931));
  INV_X1    g0731(.A(new_n454), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT16), .B1(new_n913), .B2(new_n907), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n350), .B1(new_n933), .B2(new_n915), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n934), .B2(new_n905), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n916), .A2(new_n279), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT108), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n441), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n931), .B1(new_n938), .B2(new_n703), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n918), .A2(KEYINPUT109), .A3(new_n882), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(new_n940), .A3(new_n924), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n928), .B1(new_n941), .B2(KEYINPUT37), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n497), .A2(new_n504), .B1(new_n939), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n930), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n929), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n883), .B1(new_n904), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n942), .A2(new_n930), .A3(new_n943), .ZN(new_n948));
  XOR2_X1   g0748(.A(KEYINPUT110), .B(KEYINPUT38), .Z(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT37), .B1(new_n926), .B2(new_n927), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n493), .A2(new_n495), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n493), .A2(new_n882), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(new_n922), .A4(new_n500), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n927), .B1(new_n695), .B2(new_n689), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n947), .B1(new_n948), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n690), .A2(new_n705), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n929), .A2(new_n944), .A3(KEYINPUT39), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n946), .A2(new_n961), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n756), .A2(new_n437), .A3(new_n505), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n963), .A2(new_n697), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n962), .B(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n741), .A2(new_n735), .A3(new_n742), .ZN(new_n966));
  INV_X1    g0766(.A(new_n838), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n899), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n948), .B2(new_n957), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT40), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n966), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n970), .A2(KEYINPUT40), .B1(new_n945), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n506), .A2(new_n966), .ZN(new_n974));
  OAI21_X1  g0774(.A(G330), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n974), .B2(new_n973), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n881), .B1(new_n965), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT111), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n977), .A2(new_n978), .B1(new_n965), .B2(new_n976), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n880), .B1(new_n979), .B2(new_n980), .ZN(G367));
  OAI21_X1  g0781(.A(new_n619), .B1(new_n606), .B2(new_n710), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n681), .A2(new_n705), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n716), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT45), .Z(new_n987));
  NOR2_X1   g0787(.A1(new_n716), .A2(new_n985), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(new_n713), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n715), .A2(new_n563), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n712), .B2(new_n715), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n708), .B(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n758), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n719), .B(KEYINPUT41), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n762), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n982), .A2(new_n562), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n705), .B1(new_n999), .B2(new_n618), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n985), .A2(new_n563), .A3(new_n715), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(KEYINPUT42), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT42), .B2(new_n1001), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT43), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n652), .A2(new_n705), .ZN(new_n1005));
  MUX2_X1   g0805(.A(new_n676), .B(new_n668), .S(new_n1005), .Z(new_n1006));
  OAI21_X1  g0806(.A(new_n1003), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1004), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1007), .B(new_n1008), .Z(new_n1009));
  NOR2_X1   g0809(.A1(new_n713), .A2(new_n984), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n998), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n782), .B1(new_n207), .B2(new_n419), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n237), .A2(new_n772), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n765), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n786), .A2(new_n222), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n456), .B(new_n1016), .C1(G50), .C2(new_n845), .ZN(new_n1017));
  INV_X1    g0817(.A(G137), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n804), .A2(new_n876), .B1(new_n793), .B2(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT113), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G143), .A2(new_n790), .B1(new_n798), .B2(G159), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n801), .A2(new_n216), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G150), .B2(new_n815), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT112), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1022), .B(new_n1025), .C1(KEYINPUT113), .C2(new_n1019), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n799), .A2(new_n847), .B1(new_n224), .B2(new_n801), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n791), .A2(new_n812), .B1(new_n786), .B2(new_n277), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n263), .B1(new_n793), .B2(new_n817), .C1(new_n850), .C2(new_n806), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n804), .A2(new_n280), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT46), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(G303), .C2(new_n809), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1026), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT47), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n843), .B1(new_n1034), .B2(KEYINPUT47), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1015), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1006), .A2(new_n781), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1012), .A2(new_n1039), .ZN(G387));
  NOR2_X1   g0840(.A1(new_n758), .A2(new_n994), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(new_n719), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n759), .B2(new_n995), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n762), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n712), .A2(new_n829), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n768), .A2(new_n718), .B1(G107), .B2(new_n207), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n423), .A2(G50), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT50), .ZN(new_n1048));
  AOI21_X1  g0848(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n718), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n772), .B1(new_n234), .B2(G45), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT114), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n782), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n765), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n808), .A2(new_n202), .B1(new_n806), .B2(new_n216), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G150), .B2(new_n794), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n420), .A2(new_n821), .B1(new_n790), .B2(G159), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n798), .A2(new_n348), .B1(new_n822), .B2(G77), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n263), .B1(new_n824), .B2(G97), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n801), .A2(new_n850), .B1(new_n804), .B2(new_n847), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n798), .A2(G311), .B1(new_n845), .B2(G303), .ZN(new_n1064));
  INV_X1    g0864(.A(G322), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n791), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G317), .B2(new_n809), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1063), .B1(new_n1067), .B2(KEYINPUT48), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT115), .Z(new_n1069));
  OR2_X1    g0869(.A1(new_n1067), .A2(KEYINPUT48), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(KEYINPUT49), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n545), .B1(G326), .B2(new_n794), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n280), .C2(new_n786), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT49), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1062), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1056), .B1(new_n1075), .B2(new_n778), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n995), .A2(new_n1044), .B1(new_n1045), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1043), .A2(new_n1077), .ZN(G393));
  NAND2_X1  g0878(.A1(new_n1041), .A2(new_n991), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n719), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1041), .A2(new_n991), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n991), .A2(new_n1044), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n782), .B1(new_n277), .B2(new_n207), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n241), .A2(new_n772), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n765), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n799), .A2(new_n202), .B1(new_n804), .B2(new_n216), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n801), .A2(new_n222), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1088), .A2(new_n852), .A3(new_n1089), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n423), .A2(new_n806), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n263), .B1(new_n794), .B2(G143), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(G159), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n791), .A2(new_n344), .B1(new_n1094), .B2(new_n808), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT51), .Z(new_n1096));
  AOI22_X1  g0896(.A1(G317), .A2(new_n790), .B1(new_n815), .B2(G311), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n799), .A2(new_n266), .B1(new_n280), .B2(new_n801), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n456), .B1(new_n806), .B2(new_n847), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1099), .A2(new_n787), .A3(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n804), .A2(new_n850), .B1(new_n793), .B2(new_n1065), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT116), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1093), .A2(new_n1096), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1087), .B1(new_n1107), .B2(new_n778), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n985), .B2(new_n829), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1084), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1083), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(G390));
  OAI22_X1  g0912(.A1(new_n799), .A2(new_n224), .B1(new_n791), .B2(new_n850), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n456), .B1(new_n806), .B2(new_n277), .C1(new_n280), .C2(new_n808), .ZN(new_n1114));
  NOR4_X1   g0914(.A1(new_n1113), .A2(new_n805), .A3(new_n1089), .A4(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n786), .A2(new_n216), .B1(new_n793), .B2(new_n847), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT118), .Z(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n456), .B1(new_n845), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G159), .A2(new_n821), .B1(new_n798), .B2(G137), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n815), .A2(G132), .B1(new_n794), .B2(G125), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n790), .A2(G128), .B1(new_n824), .B2(G50), .ZN(new_n1123));
  AND4_X1   g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n804), .A2(new_n344), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT53), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1115), .A2(new_n1117), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n765), .B1(new_n348), .B2(new_n844), .C1(new_n1127), .C2(new_n843), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT119), .Z(new_n1129));
  NAND2_X1  g0929(.A1(new_n958), .A2(new_n960), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n779), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n959), .B1(new_n886), .B2(new_n900), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n929), .A2(new_n944), .A3(KEYINPUT39), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n957), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT39), .B1(new_n929), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1133), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n738), .A2(new_n743), .A3(new_n838), .A4(new_n900), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n929), .A2(new_n1135), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n710), .B(new_n838), .C1(new_n750), .C2(new_n753), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n885), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n959), .B1(new_n1142), .B2(new_n900), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1139), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1137), .A2(new_n1144), .A3(KEYINPUT117), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT117), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1132), .B1(new_n958), .B2(new_n960), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n948), .A2(new_n957), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n959), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1141), .A2(new_n885), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n899), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1138), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1146), .B1(new_n1147), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1137), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n966), .A2(G330), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n968), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1145), .A2(new_n1153), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1131), .B1(new_n1160), .B2(new_n1044), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1157), .A2(new_n506), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n963), .A2(new_n1162), .A3(new_n697), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n899), .B1(new_n744), .B2(new_n967), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1158), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n886), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n899), .B1(new_n1156), .B2(new_n839), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n1150), .A3(new_n1138), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1163), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1080), .B1(new_n1160), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1154), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1159), .B1(new_n1147), .B2(new_n1171), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1147), .A2(new_n1152), .A3(new_n1146), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT117), .B1(new_n1137), .B2(new_n1144), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1172), .B(new_n1169), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1161), .B1(new_n1170), .B2(new_n1176), .ZN(G378));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1163), .B1(new_n1160), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n351), .A2(new_n882), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT55), .Z(new_n1183));
  XNOR2_X1  g0983(.A(new_n359), .B(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1184), .B(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n973), .B2(new_n737), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n946), .A2(new_n961), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n941), .A2(KEYINPUT37), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n954), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT38), .B1(new_n1191), .B2(new_n921), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n972), .B1(new_n1192), .B2(new_n948), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n966), .A2(new_n968), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n929), .B2(new_n1135), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n971), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1184), .B(new_n1185), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(G330), .A3(new_n1197), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1188), .A2(new_n1189), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1189), .B1(new_n1188), .B2(new_n1198), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1178), .B1(new_n1181), .B2(new_n1201), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n973), .A2(new_n1187), .A3(new_n737), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1197), .B1(new_n1196), .B2(G330), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n962), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1188), .A2(new_n1189), .A3(new_n1198), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1178), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1163), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1175), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n719), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1202), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1187), .A2(new_n779), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n765), .B1(new_n844), .B2(G50), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n545), .A2(G41), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G50), .B(new_n1215), .C1(new_n248), .C2(new_n249), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n815), .A2(G107), .B1(new_n794), .B2(G283), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n419), .B2(new_n806), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1023), .B(new_n1218), .C1(G77), .C2(new_n822), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n791), .A2(new_n280), .B1(new_n786), .B2(new_n876), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G97), .B2(new_n798), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1221), .A3(new_n1215), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1216), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n815), .A2(G128), .B1(new_n845), .B2(G137), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n804), .B2(new_n1118), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G150), .A2(new_n821), .B1(new_n790), .B2(G125), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT120), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(G132), .C2(new_n798), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT59), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI211_X1 g1031(.A(G33), .B(G41), .C1(new_n794), .C2(G124), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1094), .B2(new_n786), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT121), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1224), .B1(new_n1223), .B2(new_n1222), .C1(new_n1231), .C2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1214), .B1(new_n1236), .B2(new_n778), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1212), .A2(new_n1044), .B1(new_n1213), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1211), .A2(new_n1238), .ZN(G375));
  NAND2_X1  g1039(.A1(new_n899), .A2(new_n779), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n765), .B1(new_n844), .B2(G68), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n799), .A2(new_n280), .B1(new_n791), .B2(new_n847), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G97), .B2(new_n822), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n808), .A2(new_n850), .B1(new_n806), .B2(new_n224), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n267), .B(new_n1244), .C1(G303), .C2(new_n794), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1016), .B1(new_n420), .B2(new_n821), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n806), .A2(new_n344), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n263), .B(new_n1248), .C1(G128), .C2(new_n794), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n801), .A2(new_n202), .B1(new_n804), .B2(new_n1094), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G132), .B2(new_n790), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n809), .A2(G137), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n798), .A2(new_n1119), .B1(new_n824), .B2(G58), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1249), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1247), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1241), .B1(new_n1255), .B2(new_n778), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1180), .A2(new_n1044), .B1(new_n1240), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1179), .A2(new_n1163), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1169), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n997), .B(KEYINPUT123), .Z(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1257), .A2(new_n1261), .ZN(G381));
  NOR2_X1   g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1111), .A2(new_n868), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1264), .A2(new_n1265), .A3(G387), .A4(G381), .ZN(new_n1266));
  INV_X1    g1066(.A(G378), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1211), .A4(new_n1238), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(KEYINPUT124), .ZN(G407));
  NAND2_X1  g1069(.A1(new_n704), .A2(G213), .ZN(new_n1270));
  XOR2_X1   g1070(.A(new_n1270), .B(KEYINPUT125), .Z(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G375), .C2(new_n1272), .ZN(G409));
  INV_X1    g1073(.A(G387), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(G390), .A2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1111), .A2(G387), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1279), .B1(new_n1281), .B2(new_n1263), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1264), .A2(KEYINPUT127), .A3(new_n1280), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1278), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1277), .A2(new_n1282), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1258), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(KEYINPUT60), .B2(new_n1259), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1179), .A2(KEYINPUT60), .A3(new_n1163), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1080), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1257), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n868), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G384), .B(new_n1257), .C1(new_n1291), .C2(new_n1293), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1271), .A2(G2897), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1209), .A2(new_n1212), .A3(new_n1260), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G378), .B1(new_n1301), .B2(new_n1238), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT57), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1080), .B1(new_n1303), .B2(new_n1181), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G378), .B(new_n1238), .C1(new_n1304), .C2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT126), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT126), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1211), .A2(new_n1308), .A3(G378), .A4(new_n1238), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1302), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1300), .B1(new_n1310), .B2(new_n1271), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1310), .A2(new_n1271), .A3(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1289), .B(new_n1311), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1302), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1271), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1320), .A2(KEYINPUT62), .A3(new_n1312), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1288), .B1(new_n1315), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1323), .B1(new_n1320), .B2(new_n1312), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT61), .B1(new_n1320), .B2(new_n1300), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1313), .A2(KEYINPUT63), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1287), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1322), .A2(new_n1327), .ZN(G405));
  NAND2_X1  g1128(.A1(G375), .A2(new_n1267), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1316), .A2(new_n1329), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1330), .B(new_n1312), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(new_n1287), .ZN(G402));
endmodule


