//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  XNOR2_X1  g000(.A(KEYINPUT2), .B(G113), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n192), .A2(KEYINPUT67), .A3(G116), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n194), .B1(new_n189), .B2(G119), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n188), .B(new_n191), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n191), .B1(new_n195), .B2(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(new_n187), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G134), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n202), .A2(new_n203), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n205), .A2(G137), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n209), .B2(new_n201), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n215), .B2(KEYINPUT1), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT65), .A2(G143), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT65), .A2(G143), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n218), .B1(new_n221), .B2(KEYINPUT66), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n223), .B(new_n217), .C1(new_n219), .C2(new_n220), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n216), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT65), .B(G143), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n215), .B1(new_n226), .B2(new_n217), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n227), .A2(KEYINPUT1), .A3(new_n212), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n211), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT64), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT64), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(KEYINPUT0), .B2(G128), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n231), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n218), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n213), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT65), .A2(G143), .ZN(new_n238));
  AOI21_X1  g052(.A(G146), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n235), .B1(new_n239), .B2(new_n223), .ZN(new_n240));
  INV_X1    g054(.A(new_n224), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n234), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n202), .A2(new_n206), .A3(new_n207), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n208), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n219), .A2(new_n220), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n214), .B1(new_n246), .B2(G146), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT0), .A3(G128), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n242), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT30), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n229), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n250), .B1(new_n229), .B2(new_n249), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n199), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G237), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G210), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n256), .B(KEYINPUT27), .Z(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n199), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n229), .A2(new_n249), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n253), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT31), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n229), .A2(new_n249), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n199), .B1(new_n265), .B2(KEYINPUT68), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n229), .A2(new_n249), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT28), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(new_n199), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(new_n262), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n259), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n253), .A2(new_n274), .A3(new_n260), .A4(new_n262), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n264), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(G472), .A2(G902), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n269), .A2(new_n272), .A3(new_n259), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n280), .B2(KEYINPUT29), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT29), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n253), .A2(new_n262), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(new_n260), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n281), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(KEYINPUT32), .A2(new_n279), .B1(new_n285), .B2(G472), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n276), .A2(new_n287), .A3(new_n277), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n276), .B2(new_n277), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT32), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT70), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n276), .A2(new_n287), .A3(new_n277), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n293), .A2(KEYINPUT70), .A3(new_n291), .A4(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n286), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  XOR2_X1   g112(.A(new_n298), .B(KEYINPUT88), .Z(new_n299));
  INV_X1    g113(.A(KEYINPUT5), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT82), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT5), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT83), .B1(new_n304), .B2(new_n191), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n190), .A2(new_n301), .A3(new_n303), .A4(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(G113), .A3(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n304), .B(new_n191), .C1(new_n193), .C2(new_n195), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT84), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n307), .A2(G113), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n309), .A4(new_n305), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G104), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT3), .B1(new_n316), .B2(G107), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n318));
  INV_X1    g132(.A(G107), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G104), .ZN(new_n320));
  INV_X1    g134(.A(G101), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(G107), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n317), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n316), .A2(G107), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n319), .A2(G104), .ZN(new_n325));
  OAI21_X1  g139(.A(G101), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n196), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n315), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G110), .B(G122), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n332), .B(KEYINPUT85), .Z(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n317), .A2(new_n320), .A3(new_n322), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(G101), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(G101), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT4), .A3(new_n323), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n199), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n331), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G224), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(G953), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT7), .ZN(new_n345));
  INV_X1    g159(.A(new_n216), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n240), .B2(new_n241), .ZN(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT1), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n247), .A2(new_n349), .A3(G128), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n348), .B1(new_n242), .B2(new_n248), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n345), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n353), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n355), .A2(KEYINPUT7), .A3(new_n344), .A4(new_n351), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n341), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n315), .A2(new_n196), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n327), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n197), .A2(new_n300), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n330), .B1(new_n308), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n333), .B(KEYINPUT8), .Z(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n344), .B1(new_n355), .B2(new_n351), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n352), .A2(new_n343), .A3(new_n353), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT86), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT6), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n334), .B1(new_n331), .B2(new_n340), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n329), .B1(new_n311), .B2(new_n314), .ZN(new_n373));
  INV_X1    g187(.A(new_n340), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n373), .A2(new_n374), .A3(new_n333), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n371), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n333), .B1(new_n373), .B2(new_n374), .ZN(new_n377));
  INV_X1    g191(.A(new_n371), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n368), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT87), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n365), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n368), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n378), .B1(new_n341), .B2(new_n377), .ZN(new_n384));
  INV_X1    g198(.A(new_n379), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n381), .B(new_n383), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n299), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G902), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n341), .A2(new_n354), .A3(new_n356), .ZN(new_n390));
  INV_X1    g204(.A(new_n363), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n359), .B2(new_n361), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n389), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(KEYINPUT87), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n298), .A3(new_n386), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n212), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT77), .B1(new_n398), .B2(new_n247), .ZN(new_n399));
  OAI21_X1  g213(.A(G128), .B1(new_n239), .B2(new_n349), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT77), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n401), .A3(new_n227), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n402), .A3(new_n350), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n328), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT10), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n242), .A2(new_n337), .A3(new_n248), .A4(new_n339), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n327), .A2(new_n405), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n225), .B2(new_n228), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n245), .B(KEYINPUT78), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT10), .B1(new_n403), .B2(new_n328), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n407), .A2(new_n409), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n245), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G110), .B(G140), .ZN(new_n417));
  INV_X1    g231(.A(G227), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G953), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n417), .B(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT81), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n420), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n347), .A2(new_n350), .A3(new_n327), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT79), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n347), .A2(new_n428), .A3(new_n350), .A4(new_n327), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n404), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT12), .ZN(new_n431));
  INV_X1    g245(.A(new_n245), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(KEYINPUT80), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n430), .A2(new_n245), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(new_n430), .B2(new_n245), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n425), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n416), .A2(KEYINPUT81), .A3(new_n420), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n423), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G469), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n389), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n425), .A2(new_n415), .ZN(new_n441));
  INV_X1    g255(.A(new_n412), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n430), .A2(new_n245), .ZN(new_n443));
  INV_X1    g257(.A(new_n433), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n430), .A2(new_n245), .A3(new_n433), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n441), .B(G469), .C1(new_n447), .C2(new_n424), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n439), .A2(new_n389), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT9), .B(G234), .ZN(new_n452));
  OAI21_X1  g266(.A(G221), .B1(new_n452), .B2(G902), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n453), .B(KEYINPUT76), .Z(new_n454));
  OAI21_X1  g268(.A(G214), .B1(G237), .B2(G902), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n397), .A2(new_n451), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(G475), .A2(G902), .ZN(new_n457));
  INV_X1    g271(.A(G140), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G125), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n348), .A2(G140), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT16), .ZN(new_n461));
  OR3_X1    g275(.A1(new_n348), .A2(KEYINPUT16), .A3(G140), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(G146), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(G146), .B1(new_n461), .B2(new_n462), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n254), .A2(new_n255), .A3(G214), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n468), .B(new_n213), .C1(new_n236), .C2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n467), .B1(new_n226), .B2(KEYINPUT89), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT17), .A4(G131), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n471), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n203), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n470), .A2(new_n471), .A3(G131), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G113), .B(G122), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(G104), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(KEYINPUT18), .A2(G131), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n474), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n459), .A2(new_n460), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(new_n217), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT18), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n484), .B(new_n486), .C1(new_n487), .C2(new_n477), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n479), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n475), .A2(new_n477), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT71), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n463), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT71), .A4(G146), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n485), .A2(KEYINPUT19), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n485), .A2(KEYINPUT19), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n217), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n482), .B1(new_n498), .B2(new_n488), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n457), .B1(new_n489), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT20), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(new_n488), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n481), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n479), .A2(new_n482), .A3(new_n488), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n457), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n482), .B1(new_n479), .B2(new_n488), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n389), .B1(new_n489), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G475), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G217), .ZN(new_n513));
  OR3_X1    g327(.A1(new_n452), .A2(new_n513), .A3(G953), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G122), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G116), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n189), .A2(G122), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT90), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G107), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n237), .A2(G128), .A3(new_n238), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n212), .A2(G143), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n205), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n521), .A2(new_n522), .A3(new_n319), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(KEYINPUT13), .A3(new_n526), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT13), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n246), .A2(new_n531), .A3(G128), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(G134), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n530), .A2(new_n532), .A3(KEYINPUT91), .A4(G134), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n529), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n517), .A2(KEYINPUT14), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n519), .A2(new_n539), .A3(G107), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n517), .B(new_n518), .C1(KEYINPUT14), .C2(new_n319), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n525), .A2(new_n526), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G134), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n544), .B2(new_n527), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n515), .B1(new_n538), .B2(new_n546), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n514), .B(new_n545), .C1(new_n529), .C2(new_n537), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n389), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G478), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI221_X1 g366(.A(new_n389), .B1(KEYINPUT15), .B2(new_n550), .C1(new_n547), .C2(new_n548), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(G234), .A2(G237), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(G952), .A3(new_n255), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT21), .B(G898), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT92), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n555), .A2(G902), .A3(G953), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n512), .A2(new_n554), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n456), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n513), .B1(G234), .B2(new_n389), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT22), .B(G137), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n255), .A2(G221), .A3(G234), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G110), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT24), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT24), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G110), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n212), .A2(G119), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n192), .A2(G128), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n571), .B(new_n573), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT23), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n192), .B2(G128), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n212), .A2(KEYINPUT23), .A3(G119), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n192), .A2(G128), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n570), .A4(new_n580), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n576), .A2(new_n581), .B1(new_n217), .B2(new_n485), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n492), .A3(new_n493), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n578), .A2(new_n580), .A3(new_n579), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n574), .A2(new_n575), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n571), .A2(new_n573), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n584), .A2(G110), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n464), .B2(new_n465), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n583), .A2(new_n588), .A3(KEYINPUT72), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT72), .B1(new_n583), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n569), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n583), .A2(new_n588), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n568), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT25), .B1(new_n594), .B2(new_n389), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT25), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n596), .B(G902), .C1(new_n591), .C2(new_n593), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n565), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT73), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(KEYINPUT73), .B(new_n565), .C1(new_n595), .C2(new_n597), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n565), .A2(G902), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT74), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT75), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n600), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n297), .A2(new_n564), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NAND2_X1  g423(.A1(new_n451), .A2(new_n454), .ZN(new_n610));
  INV_X1    g424(.A(new_n607), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n276), .A2(new_n389), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G472), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n293), .A2(new_n613), .A3(new_n294), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n610), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n455), .ZN(new_n616));
  INV_X1    g430(.A(new_n298), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n382), .B2(new_n387), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n616), .B1(new_n618), .B2(new_n396), .ZN(new_n619));
  INV_X1    g433(.A(new_n561), .ZN(new_n620));
  INV_X1    g434(.A(new_n547), .ZN(new_n621));
  INV_X1    g435(.A(new_n548), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n621), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g440(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n626), .B(new_n627), .C1(new_n547), .C2(new_n548), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n550), .B(G902), .C1(new_n625), .C2(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n549), .A2(new_n550), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n512), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n619), .A2(new_n620), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n615), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NOR3_X1   g451(.A1(new_n382), .A2(new_n387), .A3(new_n617), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n298), .B1(new_n395), .B2(new_n386), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n455), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n501), .A2(new_n507), .B1(G475), .B2(new_n510), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n554), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n640), .A2(new_n561), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n615), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  INV_X1    g460(.A(new_n456), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n569), .A2(KEYINPUT36), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT94), .Z(new_n649));
  OR2_X1    g463(.A1(new_n589), .A2(new_n590), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n603), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n600), .A2(new_n601), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n562), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n614), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT95), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT37), .B(G110), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  NOR2_X1   g473(.A1(new_n255), .A2(G900), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(G902), .A3(new_n555), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n557), .B1(new_n662), .B2(KEYINPUT96), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(KEYINPUT96), .B2(new_n662), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n508), .A2(new_n554), .A3(new_n511), .A4(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT97), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n641), .A2(KEYINPUT97), .A3(new_n554), .A4(new_n664), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n653), .A3(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n610), .A2(new_n640), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n297), .A2(new_n670), .A3(KEYINPUT98), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n285), .A2(G472), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n673), .B1(new_n291), .B2(new_n278), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n293), .A2(new_n291), .A3(new_n294), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT70), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n674), .B1(new_n677), .B2(new_n295), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n667), .A2(new_n653), .A3(new_n668), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(new_n619), .A3(new_n451), .A4(new_n454), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n672), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n671), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NOR2_X1   g497(.A1(new_n283), .A2(new_n259), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n271), .A2(new_n262), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n685), .B(new_n389), .C1(new_n260), .C2(new_n686), .ZN(new_n687));
  AOI22_X1  g501(.A1(KEYINPUT32), .A2(new_n279), .B1(new_n687), .B2(G472), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n688), .B1(new_n292), .B2(new_n296), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT99), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n397), .B(KEYINPUT38), .Z(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n512), .A2(new_n554), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n653), .A2(new_n693), .A3(new_n616), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n451), .A2(new_n454), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n664), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n695), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n246), .ZN(G45));
  NAND2_X1  g519(.A1(new_n696), .A2(new_n653), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n678), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n632), .A2(new_n664), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n640), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  NAND2_X1  g526(.A1(new_n412), .A2(new_n424), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n445), .B2(new_n446), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT81), .B1(new_n416), .B2(new_n420), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n422), .B(new_n424), .C1(new_n412), .C2(new_n415), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(G469), .B1(new_n717), .B2(G902), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n440), .A3(new_n453), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n611), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n297), .A2(new_n634), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G15));
  NAND3_X1  g537(.A1(new_n297), .A2(new_n643), .A3(new_n720), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NOR3_X1   g539(.A1(new_n640), .A2(new_n719), .A3(new_n654), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n297), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  INV_X1    g542(.A(new_n693), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n729), .B(new_n455), .C1(new_n638), .C2(new_n639), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n718), .A2(new_n440), .A3(new_n453), .A4(new_n620), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n612), .A2(G472), .B1(new_n276), .B2(new_n277), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n607), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n516), .ZN(G24));
  INV_X1    g549(.A(new_n719), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n619), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n732), .ZN(new_n739));
  INV_X1    g553(.A(new_n653), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(new_n708), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  NAND2_X1  g557(.A1(new_n448), .A2(KEYINPUT102), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n412), .B1(new_n434), .B2(new_n435), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n745), .A2(new_n420), .B1(new_n425), .B2(new_n415), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT102), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(G469), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT103), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n440), .A4(new_n450), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n440), .A2(new_n744), .A3(new_n748), .A4(new_n450), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT103), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n278), .A2(new_n291), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n611), .B1(new_n286), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n388), .A2(new_n396), .A3(new_n453), .A4(new_n455), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n754), .A2(new_n708), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT42), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n709), .A2(KEYINPUT42), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n757), .B1(new_n751), .B2(new_n753), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n297), .A4(new_n607), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n203), .ZN(G33));
  AND2_X1   g579(.A1(new_n667), .A2(new_n668), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n762), .A2(new_n297), .A3(new_n607), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n678), .A2(new_n611), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(KEYINPUT104), .A3(new_n766), .A4(new_n762), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NAND2_X1  g587(.A1(new_n614), .A2(new_n653), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT106), .Z(new_n775));
  NOR2_X1   g589(.A1(new_n629), .A2(new_n630), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n512), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT43), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT44), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(G469), .B1(new_n746), .B2(KEYINPUT45), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n745), .A2(new_n420), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n781), .A2(KEYINPUT45), .A3(new_n441), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT105), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n783), .B1(new_n780), .B2(new_n782), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n449), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n786), .A2(KEYINPUT46), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n440), .B1(new_n786), .B2(KEYINPUT46), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n453), .B(new_n698), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n388), .A2(new_n455), .A3(new_n396), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n779), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n775), .A2(KEYINPUT44), .A3(new_n778), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(KEYINPUT107), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n792), .A2(KEYINPUT107), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT108), .B(G137), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G39));
  OAI21_X1  g611(.A(new_n453), .B1(new_n787), .B2(new_n788), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(KEYINPUT47), .B(new_n453), .C1(new_n787), .C2(new_n788), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n709), .A2(new_n607), .A3(new_n790), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n678), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  NOR2_X1   g619(.A1(G952), .A2(G953), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT114), .ZN(new_n807));
  INV_X1    g621(.A(new_n790), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n607), .A2(new_n778), .A3(new_n557), .A4(new_n732), .ZN(new_n809));
  INV_X1    g623(.A(new_n440), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n439), .B1(new_n438), .B2(new_n389), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n454), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n808), .B(new_n809), .C1(new_n802), .C2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n690), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n719), .A2(new_n790), .A3(new_n611), .A4(new_n556), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n641), .A3(new_n776), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n778), .A2(new_n557), .A3(new_n736), .A4(new_n808), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n819), .A2(new_n740), .A3(new_n739), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n455), .B1(KEYINPUT111), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n809), .A2(new_n691), .A3(new_n736), .A4(new_n822), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n821), .A2(KEYINPUT111), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n815), .A2(new_n818), .A3(new_n820), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n825), .A2(new_n818), .A3(new_n820), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(KEYINPUT51), .A3(new_n815), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n816), .A2(new_n632), .A3(new_n817), .ZN(new_n831));
  INV_X1    g645(.A(new_n756), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n819), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g647(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n834));
  OR2_X1    g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n255), .A2(G952), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n809), .B2(new_n738), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n831), .A2(new_n835), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n828), .A2(new_n830), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT98), .B1(new_n297), .B2(new_n670), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n678), .A2(new_n680), .A3(new_n672), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n742), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n664), .A2(new_n453), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n619), .A2(new_n740), .A3(new_n729), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n751), .B2(new_n753), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n689), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n711), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT52), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n741), .A2(new_n708), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n671), .A2(new_n681), .B1(new_n738), .B2(new_n853), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n707), .A2(new_n710), .B1(new_n849), .B2(new_n689), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n734), .B1(new_n297), .B2(new_n726), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n721), .A3(new_n724), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n561), .B1(new_n631), .B2(new_n642), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n397), .A3(new_n455), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n615), .A2(new_n863), .B1(new_n647), .B2(new_n655), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n608), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n760), .A2(new_n763), .ZN(new_n867));
  INV_X1    g681(.A(new_n664), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n790), .A2(new_n554), .A3(new_n512), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n707), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n762), .A2(new_n708), .A3(new_n741), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n866), .A2(new_n867), .A3(new_n772), .A4(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n843), .B1(new_n858), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT109), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n764), .B1(new_n769), .B2(new_n771), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n870), .A2(new_n871), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n879), .A2(new_n860), .A3(new_n865), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n878), .A2(new_n880), .A3(new_n852), .A4(new_n857), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(KEYINPUT109), .A3(new_n843), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT110), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n860), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n865), .A2(new_n843), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n859), .A2(new_n721), .A3(new_n724), .A4(KEYINPUT110), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n872), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n772), .A2(new_n867), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n852), .A2(new_n857), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n876), .A2(new_n877), .A3(new_n882), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n874), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n881), .A2(new_n843), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT54), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n807), .B1(new_n842), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n777), .A2(new_n454), .A3(new_n455), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT49), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n899), .B(new_n607), .C1(new_n812), .C2(new_n900), .ZN(new_n901));
  OR3_X1    g715(.A1(new_n692), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n897), .B1(new_n690), .B2(new_n902), .ZN(G75));
  AOI22_X1  g717(.A1(new_n874), .A2(new_n875), .B1(new_n890), .B2(new_n889), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n389), .B1(new_n904), .B2(new_n882), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n299), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n384), .A2(new_n385), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n368), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n394), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n255), .A2(G952), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT56), .B1(new_n905), .B2(G210), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT116), .ZN(new_n918));
  OR3_X1    g732(.A1(new_n917), .A2(new_n918), .A3(new_n912), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n917), .B2(new_n912), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(G51));
  XNOR2_X1  g735(.A(new_n449), .B(KEYINPUT57), .ZN(new_n922));
  INV_X1    g736(.A(new_n892), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n877), .B1(new_n904), .B2(new_n882), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n438), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n905), .A2(new_n785), .A3(new_n784), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n914), .B1(new_n926), .B2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n929), .A2(new_n504), .A3(new_n503), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n504), .B2(new_n503), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n914), .ZN(G60));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT59), .Z(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n625), .B2(new_n628), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n923), .B2(new_n924), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n915), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n625), .A2(new_n628), .ZN(new_n938));
  INV_X1    g752(.A(new_n934), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n896), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT117), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT117), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n942), .A2(new_n943), .A3(new_n915), .A4(new_n936), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n941), .A2(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n904), .B2(new_n882), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n948), .A2(new_n594), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n651), .B(KEYINPUT118), .Z(new_n950));
  AOI21_X1  g764(.A(new_n914), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT119), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n948), .B2(new_n950), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n949), .B(new_n951), .C1(new_n954), .C2(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  INV_X1    g772(.A(new_n866), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n255), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n559), .B2(new_n342), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(KEYINPUT120), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(KEYINPUT120), .B2(new_n960), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n908), .B1(G898), .B2(new_n255), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n963), .B(new_n964), .Z(G69));
  INV_X1    g779(.A(G900), .ZN(new_n966));
  OAI21_X1  g780(.A(G953), .B1(new_n418), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n790), .B1(new_n631), .B2(new_n642), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n770), .A2(new_n696), .A3(new_n698), .A4(new_n971), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n795), .A2(new_n804), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n854), .A2(new_n711), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n702), .A2(new_n703), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n974), .B(new_n976), .C1(new_n977), .C2(new_n695), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT62), .B1(new_n704), .B2(new_n975), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT122), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n251), .A2(new_n252), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n495), .A2(new_n496), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT121), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n985), .B(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n988), .A2(G953), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n988), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n795), .A2(new_n804), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n878), .A2(KEYINPUT124), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n832), .A2(new_n730), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OR3_X1    g810(.A1(new_n789), .A2(KEYINPUT123), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT123), .B1(new_n789), .B2(new_n996), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT124), .ZN(new_n999));
  AOI22_X1  g813(.A1(new_n997), .A2(new_n998), .B1(new_n888), .B2(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n993), .A2(new_n976), .A3(new_n994), .A4(new_n1000), .ZN(new_n1001));
  AOI211_X1 g815(.A(new_n660), .B(new_n992), .C1(new_n1001), .C2(new_n255), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n969), .B(new_n970), .C1(new_n991), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n983), .A2(new_n982), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n978), .A3(new_n973), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n989), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1001), .A2(new_n255), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1007), .B(new_n988), .C1(G900), .C2(new_n255), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1006), .A2(new_n1008), .A3(new_n968), .A4(new_n967), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1003), .A2(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  OAI21_X1  g826(.A(new_n1012), .B1(new_n1001), .B2(new_n959), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n283), .A2(new_n259), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n914), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n893), .A2(new_n894), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1012), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n1015), .A2(new_n684), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1012), .B1(new_n1005), .B2(new_n959), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT126), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1025), .A2(new_n1026), .A3(new_n684), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1018), .B1(new_n984), .B2(new_n866), .ZN(new_n1028));
  OAI21_X1  g842(.A(KEYINPUT126), .B1(new_n1028), .B2(new_n685), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1024), .B1(new_n1027), .B2(new_n1029), .ZN(G57));
endmodule


