

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U554 ( .A1(G8), .A2(n656), .ZN(n692) );
  INV_X1 U555 ( .A(n893), .ZN(n947) );
  NOR2_X2 U556 ( .A1(G164), .A2(G1384), .ZN(n697) );
  NAND2_X1 U557 ( .A1(n693), .A2(n519), .ZN(n694) );
  NOR2_X1 U558 ( .A1(n598), .A2(n597), .ZN(n599) );
  OR2_X1 U559 ( .A1(n692), .A2(n691), .ZN(n519) );
  XNOR2_X1 U560 ( .A(KEYINPUT90), .B(KEYINPUT30), .ZN(n646) );
  XNOR2_X1 U561 ( .A(n647), .B(n646), .ZN(n648) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n638) );
  XNOR2_X1 U563 ( .A(n639), .B(n638), .ZN(n644) );
  INV_X1 U564 ( .A(KEYINPUT69), .ZN(n595) );
  OR2_X1 U565 ( .A1(n695), .A2(n694), .ZN(n699) );
  XOR2_X1 U566 ( .A(KEYINPUT15), .B(n599), .Z(n600) );
  NOR2_X2 U567 ( .A1(G2105), .A2(n524), .ZN(n873) );
  XOR2_X1 U568 ( .A(KEYINPUT17), .B(n521), .Z(n876) );
  XOR2_X1 U569 ( .A(KEYINPUT0), .B(G543), .Z(n570) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n536), .Z(n776) );
  NOR2_X1 U571 ( .A1(n550), .A2(n549), .ZN(G160) );
  INV_X1 U572 ( .A(G2104), .ZN(n524) );
  NAND2_X1 U573 ( .A1(G102), .A2(n873), .ZN(n520) );
  XNOR2_X1 U574 ( .A(n520), .B(KEYINPUT82), .ZN(n523) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n876), .A2(G138), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n523), .A2(n522), .ZN(n529) );
  INV_X1 U578 ( .A(G2105), .ZN(n525) );
  NOR2_X1 U579 ( .A1(n525), .A2(n524), .ZN(n868) );
  NAND2_X1 U580 ( .A1(G114), .A2(n868), .ZN(n527) );
  NOR2_X1 U581 ( .A1(G2104), .A2(n525), .ZN(n869) );
  NAND2_X1 U582 ( .A1(G126), .A2(n869), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U584 ( .A1(n529), .A2(n528), .ZN(G164) );
  NOR2_X1 U585 ( .A1(G543), .A2(G651), .ZN(n530) );
  XOR2_X1 U586 ( .A(KEYINPUT65), .B(n530), .Z(n772) );
  NAND2_X1 U587 ( .A1(n772), .A2(G89), .ZN(n531) );
  XNOR2_X1 U588 ( .A(n531), .B(KEYINPUT4), .ZN(n533) );
  INV_X1 U589 ( .A(G651), .ZN(n535) );
  NOR2_X1 U590 ( .A1(n570), .A2(n535), .ZN(n773) );
  NAND2_X1 U591 ( .A1(G76), .A2(n773), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U593 ( .A(n534), .B(KEYINPUT5), .ZN(n542) );
  NOR2_X1 U594 ( .A1(G543), .A2(n535), .ZN(n536) );
  NAND2_X1 U595 ( .A1(G63), .A2(n776), .ZN(n539) );
  NOR2_X1 U596 ( .A1(n570), .A2(G651), .ZN(n537) );
  XNOR2_X2 U597 ( .A(n537), .B(KEYINPUT66), .ZN(n777) );
  NAND2_X1 U598 ( .A1(G51), .A2(n777), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U600 ( .A(KEYINPUT6), .B(n540), .Z(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U602 ( .A(n543), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U603 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U604 ( .A1(n868), .A2(G113), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G101), .A2(n873), .ZN(n544) );
  XOR2_X1 U606 ( .A(KEYINPUT23), .B(n544), .Z(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G125), .A2(n869), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G137), .A2(n876), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U611 ( .A1(G52), .A2(n777), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n776), .A2(G64), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G90), .A2(n772), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G77), .A2(n773), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U618 ( .A1(n557), .A2(n556), .ZN(G171) );
  INV_X1 U619 ( .A(G171), .ZN(G301) );
  NAND2_X1 U620 ( .A1(n777), .A2(G50), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT76), .B(n558), .Z(n563) );
  NAND2_X1 U622 ( .A1(G88), .A2(n772), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G75), .A2(n773), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U625 ( .A(KEYINPUT77), .B(n561), .Z(n562) );
  NOR2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n776), .A2(G62), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(G303) );
  NAND2_X1 U629 ( .A1(G651), .A2(G74), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G49), .A2(n777), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U632 ( .A1(n776), .A2(n568), .ZN(n569) );
  XNOR2_X1 U633 ( .A(n569), .B(KEYINPUT74), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G87), .A2(n570), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(G288) );
  NAND2_X1 U636 ( .A1(G73), .A2(n773), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(KEYINPUT2), .ZN(n580) );
  NAND2_X1 U638 ( .A1(G61), .A2(n776), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G48), .A2(n777), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G86), .A2(n772), .ZN(n576) );
  XNOR2_X1 U642 ( .A(KEYINPUT75), .B(n576), .ZN(n577) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(G305) );
  NAND2_X1 U645 ( .A1(G85), .A2(n772), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G72), .A2(n773), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G60), .A2(n776), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G47), .A2(n777), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  OR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(G290) );
  INV_X1 U652 ( .A(n697), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G160), .A2(G40), .ZN(n696) );
  NOR2_X2 U654 ( .A1(n587), .A2(n696), .ZN(n601) );
  INV_X1 U655 ( .A(n601), .ZN(n656) );
  BUF_X1 U656 ( .A(n601), .Z(n629) );
  NOR2_X1 U657 ( .A1(n629), .A2(G1348), .ZN(n589) );
  NOR2_X1 U658 ( .A1(G2067), .A2(n656), .ZN(n588) );
  NOR2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n618) );
  NAND2_X1 U660 ( .A1(G54), .A2(n777), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G79), .A2(n773), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U663 ( .A(KEYINPUT70), .B(n592), .ZN(n598) );
  NAND2_X1 U664 ( .A1(G66), .A2(n776), .ZN(n594) );
  NAND2_X1 U665 ( .A1(G92), .A2(n772), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n596) );
  XNOR2_X1 U667 ( .A(n596), .B(n595), .ZN(n597) );
  XOR2_X2 U668 ( .A(KEYINPUT71), .B(n600), .Z(n893) );
  AND2_X1 U669 ( .A1(n601), .A2(G1996), .ZN(n602) );
  XOR2_X1 U670 ( .A(n602), .B(KEYINPUT26), .Z(n615) );
  AND2_X1 U671 ( .A1(n656), .A2(G1341), .ZN(n613) );
  XNOR2_X1 U672 ( .A(KEYINPUT13), .B(KEYINPUT67), .ZN(n607) );
  NAND2_X1 U673 ( .A1(n772), .A2(G81), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n603), .B(KEYINPUT12), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G68), .A2(n773), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n607), .B(n606), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n776), .A2(G56), .ZN(n608) );
  XOR2_X1 U679 ( .A(KEYINPUT14), .B(n608), .Z(n609) );
  NOR2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G43), .A2(n777), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n953) );
  NOR2_X1 U683 ( .A1(n613), .A2(n953), .ZN(n614) );
  AND2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U685 ( .A(n616), .B(KEYINPUT64), .Z(n619) );
  OR2_X1 U686 ( .A1(n947), .A2(n619), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U688 ( .A1(n619), .A2(n947), .ZN(n620) );
  NAND2_X1 U689 ( .A1(n621), .A2(n620), .ZN(n633) );
  NAND2_X1 U690 ( .A1(G65), .A2(n776), .ZN(n623) );
  NAND2_X1 U691 ( .A1(G53), .A2(n777), .ZN(n622) );
  NAND2_X1 U692 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U693 ( .A1(G91), .A2(n772), .ZN(n625) );
  NAND2_X1 U694 ( .A1(G78), .A2(n773), .ZN(n624) );
  NAND2_X1 U695 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n785) );
  NAND2_X1 U697 ( .A1(n629), .A2(G2072), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n628), .B(KEYINPUT27), .ZN(n631) );
  INV_X1 U699 ( .A(G1956), .ZN(n841) );
  NOR2_X1 U700 ( .A1(n841), .A2(n629), .ZN(n630) );
  NOR2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U702 ( .A1(n785), .A2(n634), .ZN(n632) );
  NAND2_X1 U703 ( .A1(n633), .A2(n632), .ZN(n637) );
  NOR2_X1 U704 ( .A1(n785), .A2(n634), .ZN(n635) );
  XOR2_X1 U705 ( .A(n635), .B(KEYINPUT28), .Z(n636) );
  NAND2_X1 U706 ( .A1(n637), .A2(n636), .ZN(n639) );
  XOR2_X1 U707 ( .A(G1961), .B(KEYINPUT88), .Z(n965) );
  NAND2_X1 U708 ( .A1(n965), .A2(n656), .ZN(n640) );
  XNOR2_X1 U709 ( .A(n640), .B(KEYINPUT89), .ZN(n642) );
  XOR2_X1 U710 ( .A(G2078), .B(KEYINPUT25), .Z(n995) );
  NOR2_X1 U711 ( .A1(n656), .A2(n995), .ZN(n641) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n650) );
  OR2_X1 U713 ( .A1(n650), .A2(G301), .ZN(n643) );
  NAND2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n655) );
  NOR2_X1 U715 ( .A1(G1966), .A2(n692), .ZN(n669) );
  NOR2_X1 U716 ( .A1(G2084), .A2(n656), .ZN(n665) );
  NOR2_X1 U717 ( .A1(n669), .A2(n665), .ZN(n645) );
  NAND2_X1 U718 ( .A1(G8), .A2(n645), .ZN(n647) );
  NOR2_X1 U719 ( .A1(n648), .A2(G168), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n649), .B(KEYINPUT91), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n650), .A2(G301), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n653), .B(KEYINPUT31), .ZN(n654) );
  NAND2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n667) );
  NAND2_X1 U725 ( .A1(n667), .A2(G286), .ZN(n662) );
  NOR2_X1 U726 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n657), .B(KEYINPUT92), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n692), .A2(G1971), .ZN(n658) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n660), .A2(G303), .ZN(n661) );
  NAND2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n663), .A2(G8), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n664), .B(KEYINPUT32), .ZN(n673) );
  NAND2_X1 U734 ( .A1(G8), .A2(n665), .ZN(n666) );
  XOR2_X1 U735 ( .A(KEYINPUT87), .B(n666), .Z(n671) );
  INV_X1 U736 ( .A(n667), .ZN(n668) );
  NOR2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n688) );
  NOR2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n946) );
  OR2_X1 U741 ( .A1(G303), .A2(G1971), .ZN(n940) );
  INV_X1 U742 ( .A(n940), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n946), .A2(n674), .ZN(n675) );
  AND2_X1 U744 ( .A1(n688), .A2(n675), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n692), .A2(n676), .ZN(n677) );
  NAND2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n941) );
  NAND2_X1 U747 ( .A1(n677), .A2(n941), .ZN(n678) );
  INV_X1 U748 ( .A(KEYINPUT33), .ZN(n681) );
  NAND2_X1 U749 ( .A1(n678), .A2(n681), .ZN(n684) );
  INV_X1 U750 ( .A(n692), .ZN(n679) );
  NAND2_X1 U751 ( .A1(n679), .A2(n946), .ZN(n680) );
  NOR2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U753 ( .A(n682), .B(KEYINPUT93), .ZN(n683) );
  NAND2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U755 ( .A(G1981), .B(G305), .ZN(n955) );
  NOR2_X1 U756 ( .A1(n685), .A2(n955), .ZN(n695) );
  NOR2_X1 U757 ( .A1(G2090), .A2(G303), .ZN(n686) );
  NAND2_X1 U758 ( .A1(G8), .A2(n686), .ZN(n687) );
  NAND2_X1 U759 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U760 ( .A1(n692), .A2(n689), .ZN(n693) );
  NOR2_X1 U761 ( .A1(G1981), .A2(G305), .ZN(n690) );
  XOR2_X1 U762 ( .A(n690), .B(KEYINPUT24), .Z(n691) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n743) );
  XNOR2_X1 U764 ( .A(G1986), .B(G290), .ZN(n939) );
  NAND2_X1 U765 ( .A1(n743), .A2(n939), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n730) );
  NAND2_X1 U767 ( .A1(G116), .A2(n868), .ZN(n701) );
  NAND2_X1 U768 ( .A1(G128), .A2(n869), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n702), .B(KEYINPUT35), .ZN(n707) );
  NAND2_X1 U771 ( .A1(G140), .A2(n876), .ZN(n704) );
  NAND2_X1 U772 ( .A1(G104), .A2(n873), .ZN(n703) );
  NAND2_X1 U773 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U774 ( .A(KEYINPUT34), .B(n705), .Z(n706) );
  NAND2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U776 ( .A(n708), .B(KEYINPUT36), .Z(n889) );
  XNOR2_X1 U777 ( .A(KEYINPUT37), .B(G2067), .ZN(n731) );
  NOR2_X1 U778 ( .A1(n889), .A2(n731), .ZN(n914) );
  NAND2_X1 U779 ( .A1(n914), .A2(n743), .ZN(n739) );
  NAND2_X1 U780 ( .A1(G107), .A2(n868), .ZN(n710) );
  NAND2_X1 U781 ( .A1(G131), .A2(n876), .ZN(n709) );
  NAND2_X1 U782 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U783 ( .A1(G119), .A2(n869), .ZN(n712) );
  NAND2_X1 U784 ( .A1(G95), .A2(n873), .ZN(n711) );
  NAND2_X1 U785 ( .A1(n712), .A2(n711), .ZN(n713) );
  OR2_X1 U786 ( .A1(n714), .A2(n713), .ZN(n882) );
  AND2_X1 U787 ( .A1(n882), .A2(G1991), .ZN(n726) );
  NAND2_X1 U788 ( .A1(n873), .A2(G105), .ZN(n715) );
  XNOR2_X1 U789 ( .A(KEYINPUT38), .B(n715), .ZN(n721) );
  NAND2_X1 U790 ( .A1(n869), .A2(G129), .ZN(n716) );
  XOR2_X1 U791 ( .A(KEYINPUT83), .B(n716), .Z(n718) );
  NAND2_X1 U792 ( .A1(n868), .A2(G117), .ZN(n717) );
  NAND2_X1 U793 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U794 ( .A(KEYINPUT84), .B(n719), .Z(n720) );
  NAND2_X1 U795 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U796 ( .A(n722), .B(KEYINPUT85), .ZN(n724) );
  NAND2_X1 U797 ( .A1(G141), .A2(n876), .ZN(n723) );
  NAND2_X1 U798 ( .A1(n724), .A2(n723), .ZN(n883) );
  AND2_X1 U799 ( .A1(n883), .A2(G1996), .ZN(n725) );
  NOR2_X1 U800 ( .A1(n726), .A2(n725), .ZN(n912) );
  XOR2_X1 U801 ( .A(n743), .B(KEYINPUT86), .Z(n727) );
  NOR2_X1 U802 ( .A1(n912), .A2(n727), .ZN(n735) );
  INV_X1 U803 ( .A(n735), .ZN(n728) );
  NAND2_X1 U804 ( .A1(n739), .A2(n728), .ZN(n729) );
  NOR2_X1 U805 ( .A1(n730), .A2(n729), .ZN(n747) );
  AND2_X1 U806 ( .A1(n731), .A2(n889), .ZN(n732) );
  XNOR2_X1 U807 ( .A(n732), .B(KEYINPUT95), .ZN(n923) );
  NOR2_X1 U808 ( .A1(G1996), .A2(n883), .ZN(n916) );
  NOR2_X1 U809 ( .A1(G1986), .A2(G290), .ZN(n733) );
  NOR2_X1 U810 ( .A1(G1991), .A2(n882), .ZN(n909) );
  NOR2_X1 U811 ( .A1(n733), .A2(n909), .ZN(n734) );
  NOR2_X1 U812 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U813 ( .A1(n916), .A2(n736), .ZN(n737) );
  XNOR2_X1 U814 ( .A(KEYINPUT94), .B(n737), .ZN(n738) );
  XNOR2_X1 U815 ( .A(n738), .B(KEYINPUT39), .ZN(n740) );
  NAND2_X1 U816 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U817 ( .A1(n923), .A2(n741), .ZN(n742) );
  XNOR2_X1 U818 ( .A(KEYINPUT96), .B(n742), .ZN(n744) );
  NAND2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U820 ( .A(n745), .B(KEYINPUT97), .ZN(n746) );
  OR2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U822 ( .A(n748), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U823 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U824 ( .A1(G111), .A2(n868), .ZN(n750) );
  NAND2_X1 U825 ( .A1(G135), .A2(n876), .ZN(n749) );
  NAND2_X1 U826 ( .A1(n750), .A2(n749), .ZN(n753) );
  NAND2_X1 U827 ( .A1(n869), .A2(G123), .ZN(n751) );
  XOR2_X1 U828 ( .A(KEYINPUT18), .B(n751), .Z(n752) );
  NOR2_X1 U829 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U830 ( .A1(n873), .A2(G99), .ZN(n754) );
  NAND2_X1 U831 ( .A1(n755), .A2(n754), .ZN(n906) );
  XNOR2_X1 U832 ( .A(G2096), .B(n906), .ZN(n756) );
  OR2_X1 U833 ( .A1(G2100), .A2(n756), .ZN(G156) );
  INV_X1 U834 ( .A(G132), .ZN(G219) );
  INV_X1 U835 ( .A(G82), .ZN(G220) );
  INV_X1 U836 ( .A(G57), .ZN(G237) );
  INV_X1 U837 ( .A(n785), .ZN(G299) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n757) );
  XOR2_X1 U839 ( .A(n757), .B(KEYINPUT10), .Z(n905) );
  NAND2_X1 U840 ( .A1(n905), .A2(G567), .ZN(n758) );
  XOR2_X1 U841 ( .A(KEYINPUT11), .B(n758), .Z(G234) );
  INV_X1 U842 ( .A(G860), .ZN(n766) );
  NOR2_X1 U843 ( .A1(n953), .A2(n766), .ZN(n759) );
  XOR2_X1 U844 ( .A(KEYINPUT68), .B(n759), .Z(G153) );
  NOR2_X1 U845 ( .A1(G868), .A2(n947), .ZN(n761) );
  INV_X1 U846 ( .A(G868), .ZN(n763) );
  NOR2_X1 U847 ( .A1(n763), .A2(G301), .ZN(n760) );
  NOR2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U849 ( .A(KEYINPUT72), .B(n762), .ZN(G284) );
  NOR2_X1 U850 ( .A1(G286), .A2(n763), .ZN(n765) );
  NOR2_X1 U851 ( .A1(G868), .A2(G299), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(G297) );
  NAND2_X1 U853 ( .A1(n766), .A2(G559), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n767), .A2(n893), .ZN(n768) );
  XNOR2_X1 U855 ( .A(n768), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U856 ( .A1(G868), .A2(n953), .ZN(n771) );
  NAND2_X1 U857 ( .A1(G868), .A2(n893), .ZN(n769) );
  NOR2_X1 U858 ( .A1(G559), .A2(n769), .ZN(n770) );
  NOR2_X1 U859 ( .A1(n771), .A2(n770), .ZN(G282) );
  NAND2_X1 U860 ( .A1(G93), .A2(n772), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G80), .A2(n773), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n781) );
  NAND2_X1 U863 ( .A1(G67), .A2(n776), .ZN(n779) );
  NAND2_X1 U864 ( .A1(G55), .A2(n777), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n794) );
  NAND2_X1 U867 ( .A1(n893), .A2(G559), .ZN(n792) );
  XNOR2_X1 U868 ( .A(n953), .B(n792), .ZN(n782) );
  NOR2_X1 U869 ( .A1(G860), .A2(n782), .ZN(n783) );
  XOR2_X1 U870 ( .A(KEYINPUT73), .B(n783), .Z(n784) );
  XNOR2_X1 U871 ( .A(n794), .B(n784), .ZN(G145) );
  XOR2_X1 U872 ( .A(KEYINPUT19), .B(n785), .Z(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(G305), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n787), .B(G288), .ZN(n790) );
  XOR2_X1 U875 ( .A(G303), .B(n794), .Z(n788) );
  XNOR2_X1 U876 ( .A(n788), .B(G290), .ZN(n789) );
  XNOR2_X1 U877 ( .A(n790), .B(n789), .ZN(n791) );
  XNOR2_X1 U878 ( .A(n791), .B(n953), .ZN(n895) );
  XOR2_X1 U879 ( .A(n895), .B(n792), .Z(n793) );
  NAND2_X1 U880 ( .A1(G868), .A2(n793), .ZN(n796) );
  OR2_X1 U881 ( .A1(n794), .A2(G868), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n796), .A2(n795), .ZN(G295) );
  NAND2_X1 U883 ( .A1(G2078), .A2(G2084), .ZN(n798) );
  XOR2_X1 U884 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n797) );
  XNOR2_X1 U885 ( .A(n798), .B(n797), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n799), .A2(G2090), .ZN(n800) );
  XOR2_X1 U887 ( .A(KEYINPUT79), .B(n800), .Z(n801) );
  XNOR2_X1 U888 ( .A(KEYINPUT21), .B(n801), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n802), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U890 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U891 ( .A1(G69), .A2(G120), .ZN(n803) );
  NOR2_X1 U892 ( .A1(G237), .A2(n803), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G108), .A2(n804), .ZN(n827) );
  NAND2_X1 U894 ( .A1(G567), .A2(n827), .ZN(n805) );
  XNOR2_X1 U895 ( .A(KEYINPUT81), .B(n805), .ZN(n811) );
  NOR2_X1 U896 ( .A1(G220), .A2(G219), .ZN(n806) );
  XOR2_X1 U897 ( .A(KEYINPUT22), .B(n806), .Z(n807) );
  NOR2_X1 U898 ( .A1(G218), .A2(n807), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G96), .A2(n808), .ZN(n826) );
  NAND2_X1 U900 ( .A1(G2106), .A2(n826), .ZN(n809) );
  XOR2_X1 U901 ( .A(KEYINPUT80), .B(n809), .Z(n810) );
  NOR2_X1 U902 ( .A1(n811), .A2(n810), .ZN(G319) );
  INV_X1 U903 ( .A(G319), .ZN(n813) );
  NAND2_X1 U904 ( .A1(G661), .A2(G483), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n825) );
  NAND2_X1 U906 ( .A1(n825), .A2(G36), .ZN(G176) );
  XNOR2_X1 U907 ( .A(G1341), .B(G2454), .ZN(n814) );
  XNOR2_X1 U908 ( .A(n814), .B(G2430), .ZN(n815) );
  XNOR2_X1 U909 ( .A(n815), .B(G1348), .ZN(n821) );
  XOR2_X1 U910 ( .A(G2443), .B(G2427), .Z(n817) );
  XNOR2_X1 U911 ( .A(G2438), .B(G2446), .ZN(n816) );
  XNOR2_X1 U912 ( .A(n817), .B(n816), .ZN(n819) );
  XOR2_X1 U913 ( .A(G2451), .B(G2435), .Z(n818) );
  XNOR2_X1 U914 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U915 ( .A(n821), .B(n820), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n822), .A2(G14), .ZN(n898) );
  XOR2_X1 U917 ( .A(KEYINPUT98), .B(n898), .Z(G401) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n905), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U920 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G69), .ZN(G235) );
  NOR2_X1 U927 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  XOR2_X1 U929 ( .A(G2100), .B(G2096), .Z(n829) );
  XNOR2_X1 U930 ( .A(KEYINPUT42), .B(G2678), .ZN(n828) );
  XNOR2_X1 U931 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U932 ( .A(KEYINPUT43), .B(G2090), .Z(n831) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n830) );
  XNOR2_X1 U934 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U935 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2084), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(G227) );
  XOR2_X1 U938 ( .A(KEYINPUT41), .B(G1981), .Z(n837) );
  XNOR2_X1 U939 ( .A(G1966), .B(G1961), .ZN(n836) );
  XNOR2_X1 U940 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U941 ( .A(n838), .B(KEYINPUT100), .Z(n840) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n839) );
  XNOR2_X1 U943 ( .A(n840), .B(n839), .ZN(n845) );
  XOR2_X1 U944 ( .A(G1986), .B(G1976), .Z(n843) );
  XOR2_X1 U945 ( .A(n841), .B(G1971), .Z(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U947 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U948 ( .A(KEYINPUT99), .B(G2474), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G124), .A2(n869), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n848), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U952 ( .A1(G112), .A2(n868), .ZN(n849) );
  XOR2_X1 U953 ( .A(KEYINPUT101), .B(n849), .Z(n850) );
  NAND2_X1 U954 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G136), .A2(n876), .ZN(n853) );
  NAND2_X1 U956 ( .A1(G100), .A2(n873), .ZN(n852) );
  NAND2_X1 U957 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U958 ( .A1(n855), .A2(n854), .ZN(G162) );
  XOR2_X1 U959 ( .A(KEYINPUT106), .B(KEYINPUT46), .Z(n867) );
  NAND2_X1 U960 ( .A1(G118), .A2(n868), .ZN(n857) );
  NAND2_X1 U961 ( .A1(G130), .A2(n869), .ZN(n856) );
  NAND2_X1 U962 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U963 ( .A(KEYINPUT102), .B(n858), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G142), .A2(n876), .ZN(n860) );
  NAND2_X1 U965 ( .A1(G106), .A2(n873), .ZN(n859) );
  NAND2_X1 U966 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U967 ( .A(KEYINPUT45), .B(n861), .ZN(n862) );
  XNOR2_X1 U968 ( .A(KEYINPUT103), .B(n862), .ZN(n863) );
  NOR2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n865), .B(KEYINPUT48), .ZN(n866) );
  XNOR2_X1 U971 ( .A(n867), .B(n866), .ZN(n881) );
  NAND2_X1 U972 ( .A1(G115), .A2(n868), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G127), .A2(n869), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n872), .B(KEYINPUT47), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G103), .A2(n873), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n876), .A2(G139), .ZN(n877) );
  XOR2_X1 U979 ( .A(KEYINPUT104), .B(n877), .Z(n878) );
  NOR2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(KEYINPUT105), .B(n880), .Z(n926) );
  XOR2_X1 U982 ( .A(n881), .B(n926), .Z(n885) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n888) );
  XOR2_X1 U985 ( .A(G160), .B(G162), .Z(n886) );
  XNOR2_X1 U986 ( .A(n906), .B(n886), .ZN(n887) );
  XOR2_X1 U987 ( .A(n888), .B(n887), .Z(n891) );
  XOR2_X1 U988 ( .A(n889), .B(G164), .Z(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U990 ( .A1(G37), .A2(n892), .ZN(G395) );
  XOR2_X1 U991 ( .A(G301), .B(n893), .Z(n894) );
  XNOR2_X1 U992 ( .A(n894), .B(G286), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U994 ( .A1(G37), .A2(n897), .ZN(G397) );
  NAND2_X1 U995 ( .A1(G319), .A2(n898), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n899) );
  XOR2_X1 U997 ( .A(KEYINPUT49), .B(n899), .Z(n900) );
  XNOR2_X1 U998 ( .A(n900), .B(KEYINPUT107), .ZN(n901) );
  NOR2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(G108), .ZN(G238) );
  INV_X1 U1004 ( .A(n905), .ZN(G223) );
  XNOR2_X1 U1005 ( .A(G160), .B(G2084), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n910), .B(KEYINPUT108), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n921) );
  XOR2_X1 U1011 ( .A(G2090), .B(G162), .Z(n915) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1013 ( .A(KEYINPUT110), .B(n917), .Z(n919) );
  XOR2_X1 U1014 ( .A(KEYINPUT51), .B(KEYINPUT109), .Z(n918) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n922), .B(KEYINPUT111), .ZN(n924) );
  NAND2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1019 ( .A(KEYINPUT112), .B(n925), .ZN(n931) );
  XOR2_X1 U1020 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1023 ( .A(KEYINPUT50), .B(n929), .Z(n930) );
  NOR2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1025 ( .A(KEYINPUT52), .B(n932), .ZN(n933) );
  INV_X1 U1026 ( .A(KEYINPUT55), .ZN(n1014) );
  NAND2_X1 U1027 ( .A1(n933), .A2(n1014), .ZN(n934) );
  NAND2_X1 U1028 ( .A1(n934), .A2(G29), .ZN(n1022) );
  XOR2_X1 U1029 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n935) );
  XOR2_X1 U1030 ( .A(G16), .B(n935), .Z(n964) );
  XOR2_X1 U1031 ( .A(G299), .B(G1956), .Z(n937) );
  NAND2_X1 U1032 ( .A1(G1971), .A2(G303), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n945) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n943) );
  XOR2_X1 U1036 ( .A(G1961), .B(G171), .Z(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n951) );
  XNOR2_X1 U1039 ( .A(n946), .B(KEYINPUT123), .ZN(n949) );
  XOR2_X1 U1040 ( .A(G1348), .B(n947), .Z(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1043 ( .A(KEYINPUT124), .B(n952), .ZN(n962) );
  XNOR2_X1 U1044 ( .A(n953), .B(G1341), .ZN(n960) );
  XNOR2_X1 U1045 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n958) );
  XOR2_X1 U1046 ( .A(G168), .B(G1966), .Z(n954) );
  NOR2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1048 ( .A(KEYINPUT57), .B(n956), .Z(n957) );
  XNOR2_X1 U1049 ( .A(n958), .B(n957), .ZN(n959) );
  NOR2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1051 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1052 ( .A1(n964), .A2(n963), .ZN(n990) );
  INV_X1 U1053 ( .A(G16), .ZN(n988) );
  XOR2_X1 U1054 ( .A(n965), .B(G5), .Z(n967) );
  XNOR2_X1 U1055 ( .A(G21), .B(G1966), .ZN(n966) );
  NOR2_X1 U1056 ( .A1(n967), .A2(n966), .ZN(n978) );
  XOR2_X1 U1057 ( .A(G1341), .B(G19), .Z(n969) );
  XOR2_X1 U1058 ( .A(G1956), .B(G20), .Z(n968) );
  NAND2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n975) );
  XOR2_X1 U1060 ( .A(G1981), .B(G6), .Z(n973) );
  XOR2_X1 U1061 ( .A(G1348), .B(KEYINPUT125), .Z(n970) );
  XNOR2_X1 U1062 ( .A(G4), .B(n970), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(n971), .B(KEYINPUT59), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(n976), .B(KEYINPUT60), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n985) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G22), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G23), .B(G1976), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n982) );
  XOR2_X1 U1071 ( .A(G1986), .B(G24), .Z(n981) );
  NAND2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(KEYINPUT58), .B(n983), .ZN(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(KEYINPUT61), .B(n986), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n1020) );
  XNOR2_X1 U1078 ( .A(G2090), .B(G35), .ZN(n1006) );
  XNOR2_X1 U1079 ( .A(KEYINPUT113), .B(G2072), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(n991), .B(G33), .ZN(n1000) );
  XNOR2_X1 U1081 ( .A(G2067), .B(G26), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(G1991), .B(G25), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(G28), .A2(n994), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(G27), .B(n995), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(KEYINPUT114), .B(n996), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(KEYINPUT115), .B(G1996), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(G32), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(KEYINPUT53), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(KEYINPUT116), .B(n1007), .Z(n1012) );
  XOR2_X1 U1095 ( .A(G34), .B(KEYINPUT118), .Z(n1009) );
  XNOR2_X1 U1096 ( .A(G2084), .B(KEYINPUT54), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(n1009), .B(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT117), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(n1014), .B(n1013), .Z(n1016) );
  INV_X1 U1101 ( .A(G29), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(G11), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(KEYINPUT119), .B(n1018), .Z(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(n1023), .B(KEYINPUT126), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
  INV_X1 U1110 ( .A(G303), .ZN(G166) );
endmodule

