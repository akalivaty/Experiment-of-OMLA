//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G97), .A2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G58), .C2(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G1), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n223), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT0), .Z(new_n230));
  NOR3_X1   g0030(.A1(new_n222), .A2(new_n225), .A3(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  INV_X1    g0034(.A(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n210), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n209), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n250), .B1(new_n251), .B2(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n218), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT64), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n260), .B(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n254), .A2(new_n257), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n256), .A2(new_n260), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G226), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G179), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT8), .B(G58), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT65), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(new_n272), .B2(G20), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n219), .A2(KEYINPUT65), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n203), .A2(G20), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT66), .B1(G20), .B2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR3_X1   g0080(.A1(KEYINPUT66), .A2(G20), .A3(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n276), .B(new_n277), .C1(new_n278), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n224), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n218), .A2(G20), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n226), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n285), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(G50), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT67), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n283), .A2(new_n285), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n202), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n268), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n266), .A2(G169), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n263), .B2(new_n265), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(G190), .B2(new_n266), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n293), .A2(KEYINPUT69), .A3(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n291), .A2(new_n301), .A3(new_n292), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n299), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n299), .A2(new_n303), .A3(new_n307), .A4(new_n304), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n296), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n310));
  INV_X1    g0110(.A(G107), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n310), .B1(new_n311), .B2(new_n248), .C1(new_n252), .C2(new_n215), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n257), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n262), .A2(new_n259), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n264), .A2(G244), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  XOR2_X1   g0116(.A(new_n316), .B(KEYINPUT68), .Z(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n316), .B(KEYINPUT68), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n267), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n226), .A2(G20), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n218), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G1), .A2(G20), .ZN(new_n324));
  OAI21_X1  g0124(.A(G77), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n287), .ZN(new_n326));
  INV_X1    g0126(.A(new_n282), .ZN(new_n327));
  XOR2_X1   g0127(.A(KEYINPUT15), .B(G87), .Z(new_n328));
  AOI22_X1  g0128(.A1(new_n327), .A2(new_n270), .B1(new_n328), .B2(new_n275), .ZN(new_n329));
  INV_X1    g0129(.A(new_n285), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n325), .B1(G77), .B2(new_n326), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n319), .A2(new_n321), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n317), .A2(G200), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n320), .B2(G190), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n309), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n275), .A2(G77), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n339), .B1(new_n219), .B2(G68), .C1(new_n202), .C2(new_n282), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n285), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT11), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n287), .A2(new_n214), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT12), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n330), .A2(G68), .A3(new_n286), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n343), .A2(new_n345), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(KEYINPUT3), .A2(G33), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  OAI211_X1 g0151(.A(G226), .B(new_n249), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(G232), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n257), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n264), .A2(G238), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n314), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT71), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n355), .A2(new_n257), .B1(G238), .B2(new_n264), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n363), .A2(KEYINPUT71), .A3(KEYINPUT13), .A4(new_n314), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G190), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(KEYINPUT13), .A3(new_n314), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n360), .A2(G200), .A3(new_n367), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n349), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n365), .A2(G179), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT72), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n360), .A2(G169), .A3(new_n367), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n372), .A2(KEYINPUT14), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT72), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n365), .A2(new_n374), .A3(G179), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(KEYINPUT14), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n371), .A2(new_n373), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n369), .B1(new_n377), .B2(new_n348), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n309), .A2(KEYINPUT70), .A3(new_n332), .A4(new_n335), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n350), .A2(new_n351), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT7), .B1(new_n380), .B2(new_n219), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  NOR4_X1   g0182(.A1(new_n350), .A2(new_n351), .A3(new_n382), .A4(G20), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n327), .A2(G159), .ZN(new_n385));
  INV_X1    g0185(.A(G58), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n214), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n387), .B2(new_n201), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT16), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n385), .A4(new_n388), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n285), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n270), .A2(new_n286), .A3(new_n330), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n287), .A2(new_n269), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n248), .A2(G223), .A3(new_n249), .ZN(new_n397));
  INV_X1    g0197(.A(G87), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n397), .B1(new_n272), .B2(new_n398), .C1(new_n252), .C2(new_n235), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n257), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n264), .A2(G232), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n314), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n318), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n402), .A2(G179), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n396), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n396), .A2(KEYINPUT18), .A3(new_n404), .A4(new_n403), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT17), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n402), .A2(G200), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n400), .A2(G190), .A3(new_n314), .A4(new_n401), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n410), .A2(new_n411), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n393), .A2(new_n413), .A3(new_n394), .A4(new_n395), .ZN(new_n415));
  INV_X1    g0215(.A(new_n412), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT17), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n409), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n338), .A2(new_n378), .A3(new_n379), .A4(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n219), .B(G68), .C1(new_n350), .C2(new_n351), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT80), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT19), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n219), .B1(new_n354), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G87), .B2(new_n206), .ZN(new_n427));
  INV_X1    g0227(.A(G97), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n273), .B2(new_n274), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n429), .B2(KEYINPUT19), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n285), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n328), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n287), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n288), .B1(G1), .B2(new_n272), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G87), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n431), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n218), .A2(G45), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n256), .A2(G250), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT78), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n438), .B2(new_n258), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n256), .A2(new_n440), .A3(G250), .A4(new_n438), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT79), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT79), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n442), .A2(new_n446), .A3(new_n443), .ZN(new_n447));
  OAI211_X1 g0247(.A(G244), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n448));
  OAI211_X1 g0248(.A(G238), .B(new_n249), .C1(new_n350), .C2(new_n351), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G116), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n257), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n445), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G200), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n442), .A2(new_n446), .A3(new_n443), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n446), .B1(new_n442), .B2(new_n443), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(G190), .A3(new_n452), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n437), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n431), .B(new_n433), .C1(new_n434), .C2(new_n432), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n453), .A2(new_n318), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n267), .A3(new_n452), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(G257), .A3(new_n256), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT5), .B(G41), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n471), .A2(G274), .A3(new_n256), .A4(new_n466), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT76), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n470), .A2(KEYINPUT76), .A3(new_n472), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(G250), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT75), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT75), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n248), .A2(new_n480), .A3(G250), .A4(G1698), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G244), .B(new_n249), .C1(new_n350), .C2(new_n351), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT74), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n486), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n248), .A2(G244), .A3(new_n249), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n257), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n477), .A2(new_n491), .A3(KEYINPUT77), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT77), .B1(new_n477), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g0293(.A(G190), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT73), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n326), .A2(G97), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n434), .A2(new_n428), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(G107), .B1(new_n381), .B2(new_n383), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n311), .A2(KEYINPUT6), .A3(G97), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n428), .A2(new_n311), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(new_n205), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n501), .B2(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G20), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n498), .B(new_n503), .C1(new_n251), .C2(new_n282), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n497), .B1(new_n504), .B2(new_n285), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n496), .A2(new_n495), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n477), .A2(new_n491), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G200), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n494), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT77), .ZN(new_n511));
  INV_X1    g0311(.A(new_n483), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n487), .A2(new_n489), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n256), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n470), .A2(KEYINPUT76), .A3(new_n472), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT76), .B1(new_n470), .B2(new_n472), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n511), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n477), .A2(new_n491), .A3(KEYINPUT77), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n318), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n505), .A2(new_n506), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n477), .A2(new_n491), .A3(new_n267), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n464), .A2(new_n510), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT25), .B1(new_n326), .B2(G107), .ZN(new_n525));
  AND2_X1   g0325(.A1(KEYINPUT87), .A2(G87), .ZN(new_n526));
  OAI211_X1 g0326(.A(KEYINPUT22), .B(new_n526), .C1(new_n350), .C2(new_n351), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n450), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n219), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n219), .B(new_n526), .C1(new_n350), .C2(new_n351), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT22), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(G20), .A3(new_n311), .ZN(new_n534));
  NOR2_X1   g0334(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n529), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(KEYINPUT89), .A3(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n528), .A2(new_n219), .B1(new_n531), .B2(new_n530), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n538), .A2(KEYINPUT89), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(KEYINPUT89), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n540), .A2(new_n536), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n285), .A3(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G257), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n545));
  OAI211_X1 g0345(.A(G250), .B(new_n249), .C1(new_n350), .C2(new_n351), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G294), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n224), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n471), .A2(new_n466), .B1(new_n549), .B2(new_n255), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n548), .A2(new_n257), .B1(new_n550), .B2(G264), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n551), .A2(new_n472), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G190), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n326), .A2(KEYINPUT25), .A3(G107), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n435), .B2(G107), .ZN(new_n555));
  AND4_X1   g0355(.A1(new_n525), .A2(new_n544), .A3(new_n553), .A4(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n552), .A2(new_n297), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT90), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n551), .A2(G179), .A3(new_n472), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n318), .B1(new_n551), .B2(new_n472), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(KEYINPUT90), .B(new_n561), .C1(new_n552), .C2(new_n318), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n544), .A2(new_n525), .A3(new_n555), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n559), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n524), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT85), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n326), .A2(G116), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n435), .A2(G116), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n482), .B(new_n219), .C1(G33), .C2(new_n428), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT84), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n272), .A2(G97), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n578), .A2(KEYINPUT84), .A3(new_n219), .A4(new_n482), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT83), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n209), .A2(G20), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n285), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n285), .A2(new_n582), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT83), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n580), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT20), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n285), .A2(new_n581), .A3(new_n582), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n581), .B1(new_n285), .B2(new_n582), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT20), .B1(new_n591), .B2(new_n580), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n573), .B(new_n574), .C1(new_n588), .C2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(G257), .B(new_n249), .C1(new_n350), .C2(new_n351), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n248), .A2(KEYINPUT82), .A3(G257), .A4(new_n249), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n380), .A2(G303), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n248), .A2(G264), .A3(G1698), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n597), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n257), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n469), .A2(new_n256), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n472), .B1(new_n603), .B2(new_n210), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT81), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT81), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n606), .B(new_n472), .C1(new_n603), .C2(new_n210), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n602), .A2(new_n605), .A3(G179), .A4(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n571), .B1(new_n594), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n608), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(KEYINPUT85), .A3(new_n593), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n602), .A2(new_n605), .A3(new_n607), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G200), .ZN(new_n614));
  INV_X1    g0414(.A(G190), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n594), .B(new_n614), .C1(new_n615), .C2(new_n613), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n593), .A2(G169), .A3(new_n613), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n617), .A2(KEYINPUT86), .A3(KEYINPUT21), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT21), .B1(new_n617), .B2(KEYINPUT86), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n612), .B(new_n616), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n570), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n421), .A2(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n421), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n452), .A2(KEYINPUT91), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT91), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n451), .A2(new_n626), .A3(new_n257), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(G169), .B1(new_n628), .B2(new_n457), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n453), .A2(G179), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT92), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n451), .A2(new_n626), .A3(new_n257), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n626), .B1(new_n451), .B2(new_n257), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n445), .A2(new_n447), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n318), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT92), .B1(new_n637), .B2(new_n462), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n460), .B1(new_n632), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n628), .A2(new_n457), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G200), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n641), .A2(new_n458), .A3(new_n437), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n639), .A2(new_n559), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n510), .A2(new_n523), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT93), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n510), .A2(new_n523), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT93), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n637), .A2(KEYINPUT92), .A3(new_n462), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n642), .B1(new_n651), .B2(new_n460), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n647), .A2(new_n648), .A3(new_n652), .A4(new_n559), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n567), .B1(new_n563), .B2(new_n562), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n612), .B(new_n654), .C1(new_n618), .C2(new_n619), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n646), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n652), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n464), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT26), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n659), .A2(new_n661), .A3(new_n639), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n624), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n377), .A2(new_n348), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n332), .B2(new_n369), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n418), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT94), .B1(new_n407), .B2(new_n408), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n407), .A2(KEYINPUT94), .A3(new_n408), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n306), .A2(new_n308), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n296), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n664), .A2(new_n672), .ZN(G369));
  OAI21_X1  g0473(.A(new_n612), .B1(new_n618), .B2(new_n619), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n324), .A2(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n594), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n674), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n620), .B2(new_n682), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n684), .A2(KEYINPUT95), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(KEYINPUT95), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n556), .A2(new_n558), .B1(new_n566), .B2(new_n567), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n567), .A2(new_n680), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n566), .A2(new_n567), .A3(new_n680), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(G330), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n674), .A2(new_n688), .A3(new_n681), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n654), .B2(new_n680), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(KEYINPUT97), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n205), .A2(new_n398), .A3(new_n209), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT96), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n227), .A2(G41), .ZN(new_n701));
  OR3_X1    g0501(.A1(new_n700), .A2(new_n218), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n701), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(new_n223), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n698), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n698), .B2(new_n702), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT28), .Z(new_n707));
  AOI21_X1  g0507(.A(new_n680), .B1(new_n656), .B2(new_n662), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n460), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n649), .B2(new_n650), .ZN(new_n712));
  INV_X1    g0512(.A(new_n553), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n567), .A2(new_n557), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n712), .A2(new_n714), .A3(new_n642), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n612), .B(new_n568), .C1(new_n618), .C2(new_n619), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n510), .A2(KEYINPUT100), .A3(new_n523), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT100), .B1(new_n510), .B2(new_n523), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n639), .A2(new_n658), .A3(new_n643), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT26), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n658), .A2(new_n657), .A3(new_n464), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT99), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n639), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n712), .A2(KEYINPUT99), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n723), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n681), .B1(new_n720), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT29), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n710), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G330), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n457), .A2(new_n551), .A3(new_n452), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n734), .B(new_n610), .C1(new_n492), .C2(new_n493), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT30), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n518), .A2(new_n519), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n737), .A2(new_n738), .A3(new_n610), .A4(new_n734), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n640), .A2(new_n508), .A3(new_n267), .A4(new_n613), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n552), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n733), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT98), .B1(new_n744), .B2(new_n680), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n742), .B1(new_n736), .B2(new_n739), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT98), .ZN(new_n747));
  NOR4_X1   g0547(.A1(new_n746), .A2(new_n747), .A3(new_n733), .A4(new_n681), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n688), .A2(new_n523), .A3(new_n510), .A4(new_n464), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT31), .B1(new_n750), .B2(new_n620), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n740), .A2(new_n743), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n680), .B1(new_n752), .B2(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n732), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n731), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n707), .B1(new_n756), .B2(G1), .ZN(G364));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n224), .B1(G20), .B2(new_n318), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n227), .A2(new_n248), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n223), .A2(G45), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n764), .B(new_n765), .C1(new_n243), .C2(G45), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n228), .A2(G355), .A3(new_n248), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G116), .B2(new_n228), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT101), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n762), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n218), .B1(new_n322), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n701), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n219), .A2(new_n267), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G190), .A3(new_n297), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n380), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n615), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G326), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n219), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(G303), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n781), .A2(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G190), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n778), .B(new_n786), .C1(G329), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n779), .A2(G190), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(KEYINPUT33), .B(G317), .Z(new_n793));
  NAND3_X1  g0593(.A1(new_n783), .A2(new_n615), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n792), .A2(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n267), .A2(new_n297), .A3(G190), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(G294), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n775), .A2(new_n787), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n790), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n794), .A2(new_n311), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n789), .A2(G159), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT32), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n803), .B(new_n805), .C1(G68), .C2(new_n791), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n776), .A2(new_n386), .B1(new_n801), .B2(new_n251), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT102), .Z(new_n808));
  INV_X1    g0608(.A(new_n798), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n248), .B1(new_n809), .B2(new_n428), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G50), .B2(new_n780), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n806), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n784), .A2(new_n398), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n802), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n774), .B1(new_n814), .B2(new_n761), .ZN(new_n815));
  INV_X1    g0615(.A(new_n760), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n770), .B(new_n815), .C1(new_n687), .C2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(G330), .B1(new_n685), .B2(new_n686), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n774), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n687), .A2(G330), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(G396));
  NAND4_X1  g0621(.A1(new_n319), .A2(new_n321), .A3(new_n331), .A4(new_n681), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n319), .A2(new_n321), .A3(new_n331), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n333), .A2(new_n334), .B1(new_n331), .B2(new_n680), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n708), .A2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n680), .B(new_n825), .C1(new_n656), .C2(new_n662), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(new_n755), .Z(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n774), .ZN(new_n831));
  INV_X1    g0631(.A(new_n801), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n780), .A2(G137), .B1(new_n832), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n834), .B2(new_n776), .C1(new_n278), .C2(new_n792), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT34), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n809), .A2(new_n386), .B1(new_n794), .B2(new_n214), .ZN(new_n837));
  INV_X1    g0637(.A(new_n784), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n380), .B(new_n837), .C1(G50), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n836), .B(new_n839), .C1(new_n840), .C2(new_n788), .ZN(new_n841));
  INV_X1    g0641(.A(G294), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n776), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(KEYINPUT103), .B(G283), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n792), .A2(new_n845), .B1(new_n781), .B2(new_n785), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G107), .B2(new_n838), .ZN(new_n847));
  INV_X1    g0647(.A(new_n794), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G87), .B1(new_n798), .B2(G97), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n380), .B1(new_n801), .B2(new_n209), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G311), .B2(new_n789), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n847), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n841), .B1(new_n843), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n774), .B1(new_n853), .B2(new_n761), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n761), .A2(new_n758), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n854), .B1(G77), .B2(new_n856), .C1(new_n826), .C2(new_n759), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n831), .A2(new_n857), .ZN(G384));
  OAI211_X1 g0658(.A(G20), .B(new_n549), .C1(new_n502), .C2(KEYINPUT35), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n209), .B(new_n859), .C1(KEYINPUT35), .C2(new_n502), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT36), .Z(new_n861));
  OAI21_X1  g0661(.A(G77), .B1(new_n386), .B2(new_n214), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n862), .A2(new_n223), .B1(G50), .B2(new_n214), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(G1), .A3(new_n226), .ZN(new_n864));
  INV_X1    g0664(.A(new_n678), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n396), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n405), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n415), .A2(new_n416), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT37), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n868), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(new_n405), .A4(new_n866), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n866), .B1(new_n409), .B2(new_n418), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n869), .A2(new_n872), .ZN(new_n877));
  INV_X1    g0677(.A(new_n418), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT94), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n409), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n407), .A2(KEYINPUT94), .A3(new_n408), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n877), .B1(new_n882), .B2(new_n866), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n876), .B1(new_n883), .B2(new_n874), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n349), .A2(new_n681), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n378), .A2(new_n886), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n885), .B(new_n369), .C1(new_n377), .C2(new_n348), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n681), .B1(new_n746), .B2(new_n733), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n622), .B2(KEYINPUT31), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n746), .A2(new_n733), .A3(new_n681), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n889), .B(new_n826), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT40), .B1(new_n884), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n751), .B2(new_n753), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n887), .A2(new_n888), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n895), .A2(new_n825), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n874), .B1(new_n873), .B2(new_n875), .ZN(new_n899));
  INV_X1    g0699(.A(new_n875), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(KEYINPUT38), .A3(new_n877), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n894), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n421), .A2(new_n895), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n904), .B(new_n905), .Z(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(G330), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n880), .A2(new_n881), .A3(new_n678), .ZN(new_n908));
  INV_X1    g0708(.A(new_n822), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n889), .B(new_n902), .C1(new_n828), .C2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n899), .B2(new_n901), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n884), .B2(new_n911), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n665), .A2(new_n680), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n908), .B(new_n910), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n907), .B(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT104), .B1(new_n731), .B2(new_n624), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT104), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n920), .B(new_n421), .C1(new_n710), .C2(new_n730), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n672), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n918), .B(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n861), .B(new_n864), .C1(new_n925), .C2(new_n323), .ZN(G367));
  AOI22_X1  g0726(.A1(new_n791), .A2(G159), .B1(new_n838), .B2(G58), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n834), .B2(new_n781), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n809), .A2(new_n214), .B1(new_n794), .B2(new_n251), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n248), .B1(new_n801), .B2(new_n202), .C1(new_n278), .C2(new_n776), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(G137), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n931), .B1(new_n932), .B2(new_n788), .ZN(new_n933));
  INV_X1    g0733(.A(G317), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n788), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n784), .A2(new_n209), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n380), .B1(new_n785), .B2(new_n776), .C1(new_n936), .C2(KEYINPUT46), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n935), .B(new_n937), .C1(KEYINPUT46), .C2(new_n936), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n794), .A2(new_n428), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n792), .A2(new_n842), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n832), .A2(new_n844), .B1(G107), .B2(new_n798), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n939), .B(new_n940), .C1(KEYINPUT109), .C2(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n938), .B(new_n943), .C1(KEYINPUT109), .C2(new_n942), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n781), .A2(new_n800), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n933), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT47), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n774), .B1(new_n947), .B2(new_n761), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n762), .B1(new_n228), .B2(new_n432), .C1(new_n239), .C2(new_n764), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n639), .A2(new_n437), .A3(new_n681), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n652), .B1(new_n437), .B2(new_n681), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n948), .B(new_n949), .C1(new_n816), .C2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n658), .A2(new_n680), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT105), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n717), .A2(new_n718), .B1(new_n507), .B2(new_n681), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n694), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT42), .Z(new_n962));
  INV_X1    g0762(.A(new_n959), .ZN(new_n963));
  OAI211_X1 g0763(.A(KEYINPUT106), .B(new_n523), .C1(new_n963), .C2(new_n568), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT106), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n568), .B1(new_n957), .B2(new_n958), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(new_n966), .B2(new_n658), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n964), .A2(new_n681), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n692), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n818), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n959), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n969), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n972), .B1(new_n969), .B2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n955), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n969), .A2(new_n973), .ZN(new_n978));
  INV_X1    g0778(.A(new_n972), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n954), .A3(new_n974), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT44), .B1(new_n963), .B2(new_n695), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT44), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n959), .A2(new_n696), .A3(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n987));
  NAND3_X1  g0787(.A1(new_n959), .A2(new_n696), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n987), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n963), .B2(new_n695), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n986), .A2(new_n693), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n983), .A2(new_n985), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n988), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n971), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n674), .A2(new_n681), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n694), .B1(new_n997), .B2(new_n692), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n818), .B(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n756), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n701), .B(KEYINPUT41), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n771), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT108), .B1(new_n982), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n977), .A2(new_n981), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n772), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT108), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n953), .B1(new_n1004), .B2(new_n1008), .ZN(G387));
  INV_X1    g0809(.A(new_n756), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(new_n999), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n999), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n701), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n798), .A2(new_n844), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n776), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1016), .A2(G317), .B1(new_n832), .B2(G303), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1017), .A2(KEYINPUT110), .B1(G311), .B2(new_n791), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(KEYINPUT110), .B2(new_n1017), .C1(new_n777), .C2(new_n781), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT48), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1015), .B1(new_n842), .B2(new_n784), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT111), .Z(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n1025));
  XNOR2_X1  g0825(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n248), .B1(new_n848), .B2(G116), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n782), .C2(new_n788), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n776), .A2(new_n202), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n248), .B1(new_n788), .B2(new_n278), .C1(new_n214), .C2(new_n801), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n939), .B(new_n1030), .C1(G77), .C2(new_n838), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n780), .A2(G159), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n791), .A2(new_n270), .B1(new_n328), .B2(new_n798), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1028), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n761), .ZN(new_n1036));
  OR3_X1    g0836(.A1(new_n269), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT50), .B1(new_n269), .B2(G50), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n465), .A3(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n700), .B(new_n1039), .C1(G68), .C2(G77), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n763), .B1(new_n236), .B2(new_n465), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n700), .A2(new_n228), .A3(new_n248), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n228), .A2(G107), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n762), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n774), .B1(new_n970), .B2(new_n760), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1036), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1014), .B(new_n1047), .C1(new_n771), .C2(new_n999), .ZN(G393));
  INV_X1    g0848(.A(new_n995), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n772), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n959), .A2(new_n816), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT113), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n762), .B1(new_n428), .B2(new_n228), .C1(new_n246), .C2(new_n764), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(KEYINPUT113), .ZN(new_n1054));
  INV_X1    g0854(.A(G159), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n781), .A2(new_n278), .B1(new_n1055), .B2(new_n776), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT51), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n809), .A2(new_n251), .B1(new_n794), .B2(new_n398), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n248), .B1(new_n788), .B2(new_n834), .C1(new_n269), .C2(new_n801), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(G50), .C2(new_n791), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1057), .B(new_n1060), .C1(new_n214), .C2(new_n784), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n781), .A2(new_n934), .B1(new_n800), .B2(new_n776), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT52), .Z(new_n1063));
  OAI221_X1 g0863(.A(new_n380), .B1(new_n788), .B2(new_n777), .C1(new_n842), .C2(new_n801), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n803), .B1(G116), .B2(new_n798), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n784), .B2(new_n845), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n792), .A2(new_n785), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1061), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n774), .B1(new_n1069), .B2(new_n761), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1012), .A2(new_n995), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT114), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n701), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1049), .A2(new_n1011), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n1072), .B2(KEYINPUT114), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1050), .B(new_n1071), .C1(new_n1074), .C2(new_n1076), .ZN(G390));
  AOI21_X1  g0877(.A(new_n909), .B1(new_n708), .B2(new_n826), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n915), .B1(new_n1078), .B2(new_n896), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n913), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n747), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n892), .A2(KEYINPUT98), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n733), .B1(new_n570), .B2(new_n621), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1082), .B(new_n1083), .C1(new_n1084), .C2(new_n890), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1085), .A2(G330), .A3(new_n826), .A4(new_n889), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT116), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n755), .A2(KEYINPUT116), .A3(new_n826), .A4(new_n889), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n884), .A2(new_n914), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n824), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n332), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n681), .B(new_n1093), .C1(new_n720), .C2(new_n728), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n822), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n889), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT115), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n418), .B1(new_n669), .B2(new_n668), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n866), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT38), .B1(new_n1100), .B2(new_n877), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n915), .B1(new_n1101), .B2(new_n876), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n896), .B1(new_n1094), .B2(new_n822), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT115), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1080), .B(new_n1090), .C1(new_n1097), .C2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1091), .A2(KEYINPUT115), .A3(new_n1096), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1104), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1107), .A2(new_n1108), .B1(new_n913), .B2(new_n1079), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n897), .A2(G330), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1106), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n772), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n913), .A2(new_n758), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n781), .A2(new_n795), .B1(new_n251), .B2(new_n809), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G107), .B2(new_n791), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n832), .A2(G97), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n813), .B1(G68), .B2(new_n848), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n380), .B1(new_n788), .B2(new_n842), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G116), .B2(new_n1016), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n784), .A2(new_n278), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT53), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n776), .A2(new_n840), .B1(new_n801), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G125), .B2(new_n789), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n791), .A2(G137), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n780), .A2(G128), .B1(G159), .B2(new_n798), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1123), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n248), .B1(new_n794), .B2(new_n202), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT117), .Z(new_n1131));
  OAI21_X1  g0931(.A(new_n1121), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n774), .B1(new_n1132), .B2(new_n761), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1114), .B(new_n1133), .C1(new_n270), .C2(new_n856), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1113), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n905), .A2(G330), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n672), .B(new_n1136), .C1(new_n919), .C2(new_n921), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1085), .A2(G330), .A3(new_n826), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n896), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1078), .B1(new_n1139), .B2(new_n1110), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n895), .A2(new_n825), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n889), .B1(new_n1141), .B2(G330), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1095), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1140), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1137), .A2(new_n1145), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1112), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n703), .B1(new_n1112), .B2(new_n1146), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1135), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(G378));
  AOI21_X1  g0950(.A(new_n873), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n901), .B1(new_n1151), .B2(KEYINPUT38), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n898), .B1(new_n1152), .B2(new_n897), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT38), .B1(new_n900), .B2(new_n877), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n898), .B1(new_n876), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n893), .ZN(new_n1156));
  OAI21_X1  g0956(.A(G330), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT56), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT55), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n293), .A2(new_n865), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n309), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n296), .B(new_n1162), .C1(new_n306), .C2(new_n308), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1159), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n309), .A2(new_n1160), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1166), .A2(new_n1163), .A3(KEYINPUT55), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1158), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1161), .A2(new_n1164), .A3(new_n1159), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT55), .B1(new_n1166), .B2(new_n1163), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n1170), .A3(KEYINPUT56), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1157), .A2(new_n1172), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1174), .B(G330), .C1(new_n1153), .C2(new_n1156), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n916), .A3(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1176), .A2(KEYINPUT121), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(KEYINPUT121), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT120), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n1180), .B2(new_n917), .ZN(new_n1181));
  AOI211_X1 g0981(.A(KEYINPUT120), .B(new_n916), .C1(new_n1173), .C2(new_n1175), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1177), .A2(new_n1178), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1112), .A2(new_n1146), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1137), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n703), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1180), .A2(new_n917), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT119), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n1176), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1173), .A2(KEYINPUT119), .A3(new_n916), .A4(new_n1175), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1137), .B1(new_n1112), .B2(new_n1146), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1184), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1188), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1191), .A2(new_n772), .A3(new_n1192), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n380), .B1(new_n788), .B2(new_n795), .C1(new_n386), .C2(new_n794), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G41), .B(new_n1198), .C1(G77), .C2(new_n838), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT118), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1016), .A2(G107), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n791), .A2(G97), .B1(new_n780), .B2(G116), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n832), .A2(new_n328), .B1(G68), .B2(new_n798), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT58), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n202), .B1(new_n350), .B2(G41), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n780), .A2(G125), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n784), .B2(new_n1124), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n791), .A2(G132), .B1(new_n832), .B2(G137), .ZN(new_n1209));
  INV_X1    g1009(.A(G128), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1209), .B1(new_n1210), .B2(new_n776), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1208), .B(new_n1211), .C1(G150), .C2(new_n798), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT59), .ZN(new_n1213));
  AOI21_X1  g1013(.A(G41), .B1(new_n848), .B2(G159), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G33), .B1(new_n789), .B2(G124), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1205), .A2(new_n1206), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n774), .B1(new_n1217), .B2(new_n761), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(G50), .B2(new_n856), .C1(new_n1172), .C2(new_n759), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1197), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1196), .A2(new_n1221), .ZN(G375));
  INV_X1    g1022(.A(KEYINPUT122), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n889), .B2(new_n759), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n855), .A2(new_n214), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n896), .A2(KEYINPUT122), .A3(new_n758), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n776), .A2(new_n795), .B1(new_n801), .B2(new_n311), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n791), .A2(G116), .B1(new_n328), .B2(new_n798), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n428), .B2(new_n784), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(G303), .C2(new_n789), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n380), .B1(new_n794), .B2(new_n251), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT123), .Z(new_n1232));
  OAI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(new_n842), .C2(new_n781), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n248), .B1(new_n801), .B2(new_n278), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n781), .A2(new_n840), .B1(new_n794), .B2(new_n386), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(G137), .C2(new_n1016), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n792), .A2(new_n1124), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n809), .A2(new_n202), .B1(new_n784), .B2(new_n1055), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1236), .B(new_n1239), .C1(new_n1210), .C2(new_n788), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1233), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n774), .B1(new_n1241), .B2(new_n761), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1145), .B2(new_n771), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT124), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT124), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1246), .B(new_n1243), .C1(new_n1145), .C2(new_n771), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1146), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1137), .A2(new_n1145), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1001), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(G381));
  AOI21_X1  g1052(.A(new_n1220), .B1(new_n1188), .B2(new_n1195), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1149), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NOR4_X1   g1055(.A1(G387), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(G381), .A2(G384), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(G407));
  NAND2_X1  g1058(.A1(new_n1255), .A2(new_n679), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(G407), .A2(G213), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT125), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(G407), .A2(new_n1259), .A3(new_n1262), .A4(G213), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(G409));
  INV_X1    g1064(.A(G213), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(G343), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1183), .A2(new_n772), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1269), .A2(new_n1001), .A3(new_n1192), .A4(new_n1191), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1149), .A2(new_n1268), .A3(new_n1270), .A4(new_n1219), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1267), .B(new_n1271), .C1(new_n1253), .C2(new_n1149), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1249), .B1(new_n1273), .B2(KEYINPUT60), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1137), .B2(new_n1145), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n701), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1248), .B(G384), .C1(new_n1274), .C2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1146), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1273), .A2(KEYINPUT60), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n701), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1283), .B2(new_n1248), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT63), .B1(new_n1272), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G375), .A2(G378), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1291));
  AND4_X1   g1091(.A1(new_n1113), .A2(new_n1291), .A3(new_n1134), .A4(new_n1219), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1266), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1288), .A2(new_n1289), .A3(new_n1293), .A4(new_n1285), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1287), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1288), .A2(KEYINPUT127), .A3(new_n1293), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1149), .B1(new_n1196), .B2(new_n1221), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1271), .A2(new_n1267), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1266), .A2(G2897), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1248), .B1(new_n1274), .B2(new_n1278), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(new_n831), .A3(new_n857), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1301), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n1279), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1296), .A2(new_n1300), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT61), .ZN(new_n1309));
  INV_X1    g1109(.A(G390), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G387), .A2(new_n1310), .ZN(new_n1311));
  XOR2_X1   g1111(.A(G393), .B(G396), .Z(new_n1312));
  OAI211_X1 g1112(.A(G390), .B(new_n953), .C1(new_n1004), .C2(new_n1008), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1312), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1295), .A2(new_n1308), .A3(new_n1309), .A4(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(KEYINPUT62), .B1(new_n1272), .B2(new_n1286), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT61), .B1(new_n1272), .B2(new_n1307), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1288), .A2(new_n1320), .A3(new_n1293), .A4(new_n1285), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1318), .A2(new_n1319), .A3(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1316), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1317), .A2(new_n1324), .ZN(G405));
  OAI21_X1  g1125(.A(new_n1285), .B1(new_n1255), .B2(new_n1298), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1288), .A2(new_n1254), .A3(new_n1286), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1316), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1316), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(G402));
endmodule


