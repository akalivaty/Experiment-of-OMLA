//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n214), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n214), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n212), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n206), .A2(new_n207), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n222), .B(new_n225), .C1(new_n227), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G226), .B(G232), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  AOI22_X1  g0046(.A1(new_n246), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT67), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n248), .B1(new_n249), .B2(G20), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n212), .A2(KEYINPUT67), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n226), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT11), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT12), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(new_n260), .B2(G68), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n256), .B1(new_n211), .B2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n262), .B(new_n264), .C1(new_n266), .C2(new_n202), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT74), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n268), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n259), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G232), .A3(G1698), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G97), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G226), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n273), .B(new_n274), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT66), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n279), .A2(KEYINPUT66), .A3(G1), .A4(G13), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT13), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n280), .A2(new_n287), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n290), .B1(new_n292), .B2(G238), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n285), .A2(new_n286), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n286), .B1(new_n285), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g0095(.A(G200), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n285), .A2(new_n293), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n286), .A2(KEYINPUT73), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n285), .B(new_n293), .C1(KEYINPUT73), .C2(new_n286), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G190), .A3(new_n300), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n271), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(G169), .B1(new_n294), .B2(new_n295), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT14), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n305), .B(G169), .C1(new_n294), .C2(new_n295), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n299), .A2(G179), .A3(new_n300), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n271), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n302), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n289), .B1(new_n291), .B2(new_n277), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n272), .A2(G223), .A3(G1698), .ZN(new_n312));
  INV_X1    g0112(.A(G222), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n312), .B1(new_n253), .B2(new_n272), .C1(new_n276), .C2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n314), .B2(new_n284), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(G179), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n261), .A2(new_n207), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n266), .B2(new_n207), .ZN(new_n319));
  INV_X1    g0119(.A(new_n252), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n320), .A2(new_n322), .B1(G150), .B2(new_n246), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n208), .A2(G20), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n319), .B1(new_n325), .B2(new_n256), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n315), .A2(G169), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n317), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n326), .A2(KEYINPUT9), .B1(new_n315), .B2(G190), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  OAI22_X1  g0131(.A1(new_n326), .A2(KEYINPUT9), .B1(new_n315), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT10), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n326), .A2(KEYINPUT9), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT10), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n316), .A2(G200), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n334), .A2(new_n329), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n328), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G244), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n289), .B1(new_n291), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n272), .A2(G232), .A3(new_n275), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n272), .A2(G238), .A3(G1698), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT68), .B(G107), .Z(new_n343));
  OAI211_X1 g0143(.A(new_n341), .B(new_n342), .C1(new_n272), .C2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n340), .B1(new_n344), .B2(new_n284), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n331), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n252), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n246), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n321), .A2(new_n349), .B1(new_n212), .B2(new_n253), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n256), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n211), .A2(G20), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n352), .A2(new_n255), .A3(G77), .A4(new_n226), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT69), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n261), .A2(new_n253), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n351), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT70), .B1(new_n346), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n356), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT70), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n358), .B(new_n359), .C1(new_n331), .C2(new_n345), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n345), .A2(G190), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n356), .B1(new_n345), .B2(G169), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT71), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n356), .B(KEYINPUT71), .C1(new_n345), .C2(G169), .ZN(new_n366));
  INV_X1    g0166(.A(G179), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n345), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n362), .A2(new_n369), .A3(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n362), .A2(new_n369), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT72), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n310), .A2(new_n338), .A3(new_n370), .A4(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n322), .A2(new_n261), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n266), .B2(new_n322), .ZN(new_n376));
  INV_X1    g0176(.A(new_n256), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n201), .A2(new_n202), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n206), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n246), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G33), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT7), .B1(new_n385), .B2(new_n212), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT75), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n202), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n272), .B2(G20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT75), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n381), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n377), .B1(new_n393), .B2(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n202), .B1(new_n390), .B2(new_n391), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(new_n381), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n376), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT78), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n280), .A2(G232), .A3(new_n287), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n289), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n399), .B1(new_n289), .B2(new_n400), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n401), .A2(new_n402), .A3(G190), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n382), .A2(new_n384), .A3(G223), .A4(new_n275), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT76), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n272), .A2(KEYINPUT76), .A3(G223), .A4(new_n275), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n272), .A2(G226), .A3(G1698), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n406), .A2(new_n407), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT77), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n410), .A2(new_n411), .A3(new_n284), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n410), .B2(new_n284), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n403), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n284), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n401), .A2(new_n402), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n331), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT79), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n398), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n398), .A2(new_n419), .A3(new_n420), .A4(KEYINPUT17), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(G169), .B1(new_n415), .B2(new_n416), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n415), .A2(KEYINPUT77), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n410), .A2(new_n411), .A3(new_n284), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n416), .A2(new_n367), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n426), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n379), .A2(new_n380), .ZN(new_n433));
  INV_X1    g0233(.A(new_n392), .ZN(new_n434));
  OAI21_X1  g0234(.A(G68), .B1(new_n390), .B2(KEYINPUT75), .ZN(new_n435));
  OAI211_X1 g0235(.A(KEYINPUT16), .B(new_n433), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(new_n397), .A3(new_n256), .ZN(new_n437));
  INV_X1    g0237(.A(new_n376), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n432), .A2(new_n439), .A3(KEYINPUT18), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT18), .B1(new_n432), .B2(new_n439), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n425), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT80), .B1(new_n374), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n338), .A2(new_n370), .A3(new_n373), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT80), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n423), .A2(new_n424), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n440), .A2(new_n441), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n445), .A2(new_n446), .A3(new_n449), .A4(new_n310), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT21), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n272), .A2(G264), .A3(G1698), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n385), .A2(G303), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n382), .A2(new_n384), .A3(G257), .A4(new_n275), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n284), .ZN(new_n457));
  XOR2_X1   g0257(.A(KEYINPUT5), .B(G41), .Z(new_n458));
  NAND3_X1  g0258(.A1(new_n211), .A2(G45), .A3(G274), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OR2_X1    g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n280), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n211), .A2(G45), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n280), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n460), .B1(new_n466), .B2(G270), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n457), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G169), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n260), .A2(G116), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n211), .A2(G33), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n377), .A2(new_n260), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n212), .C1(G33), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT84), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n249), .A2(G97), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(KEYINPUT84), .A3(new_n212), .A4(new_n476), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n255), .A2(new_n226), .B1(G20), .B2(new_n474), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT20), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n480), .A2(KEYINPUT20), .A3(new_n482), .A4(new_n483), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n475), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n452), .B1(new_n469), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n487), .ZN(new_n490));
  INV_X1    g0290(.A(new_n475), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(KEYINPUT21), .A3(G169), .A4(new_n468), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n457), .A2(new_n467), .A3(G179), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n492), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n489), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT85), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n331), .B1(new_n457), .B2(new_n467), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n457), .A2(new_n467), .ZN(new_n500));
  OAI211_X1 g0300(.A(KEYINPUT85), .B(new_n488), .C1(new_n500), .C2(new_n331), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(G190), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT86), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT86), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n499), .A2(new_n501), .A3(new_n505), .A4(new_n502), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n496), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n272), .A2(new_n212), .A3(G87), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT22), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT22), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n272), .A2(new_n510), .A3(new_n212), .A4(G87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  INV_X1    g0313(.A(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(G20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G116), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(G20), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n343), .A2(G20), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(KEYINPUT23), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g0320(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n521), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n512), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n256), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n261), .A2(new_n514), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n526), .A2(KEYINPUT25), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(KEYINPUT25), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n528), .C1(new_n514), .C2(new_n473), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n460), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n382), .A2(new_n384), .A3(G257), .A4(G1698), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT88), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n272), .A2(KEYINPUT88), .A3(G257), .A4(G1698), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G294), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n272), .A2(G250), .A3(new_n275), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n535), .A2(new_n536), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n284), .ZN(new_n540));
  INV_X1    g0340(.A(G264), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n463), .B2(new_n465), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT90), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT90), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n545), .B(new_n542), .C1(new_n539), .C2(new_n284), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n532), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n331), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n542), .B1(new_n539), .B2(new_n284), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n532), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT89), .ZN(new_n551));
  INV_X1    g0351(.A(G190), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT89), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n549), .A2(new_n553), .A3(new_n532), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n531), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n524), .A2(new_n256), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n529), .B1(new_n557), .B2(new_n522), .ZN(new_n558));
  AND4_X1   g0358(.A1(new_n553), .A2(new_n540), .A3(new_n532), .A4(new_n543), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n553), .B1(new_n549), .B2(new_n532), .ZN(new_n560));
  OAI21_X1  g0360(.A(G169), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G179), .B(new_n532), .C1(new_n544), .C2(new_n546), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n382), .A2(new_n384), .A3(G250), .A4(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n382), .A2(new_n384), .A3(G244), .A4(new_n275), .ZN(new_n566));
  NOR2_X1   g0366(.A1(KEYINPUT81), .A2(KEYINPUT4), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n476), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n284), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n460), .B1(new_n466), .B2(G257), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G169), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(new_n367), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n246), .A2(G77), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT6), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n577), .A2(new_n477), .A3(G107), .ZN(new_n578));
  XNOR2_X1  g0378(.A(G97), .B(G107), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n576), .B1(new_n580), .B2(new_n212), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n343), .B1(new_n390), .B2(new_n391), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n256), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n260), .A2(G97), .ZN(new_n584));
  INV_X1    g0384(.A(new_n473), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(G97), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n574), .A2(new_n575), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n570), .A2(G190), .A3(new_n571), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(new_n583), .A3(new_n586), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n331), .B1(new_n570), .B2(new_n571), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT82), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n583), .A2(new_n586), .ZN(new_n593));
  INV_X1    g0393(.A(new_n591), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT82), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .A4(new_n589), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n588), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT83), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n382), .A2(new_n384), .A3(G244), .A4(G1698), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n382), .A2(new_n384), .A3(G238), .A4(new_n275), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(new_n516), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n284), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n280), .A2(G250), .A3(new_n464), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n459), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n598), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n602), .A2(new_n598), .A3(new_n605), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n573), .A3(new_n608), .ZN(new_n609));
  AOI211_X1 g0409(.A(KEYINPUT83), .B(new_n604), .C1(new_n601), .C2(new_n284), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n367), .B1(new_n610), .B2(new_n606), .ZN(new_n611));
  INV_X1    g0411(.A(new_n347), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n260), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT19), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n252), .B2(new_n477), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n272), .A2(new_n212), .A3(G68), .ZN(new_n616));
  XNOR2_X1  g0416(.A(KEYINPUT68), .B(G107), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n617), .A2(G87), .A3(G97), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n274), .A2(new_n614), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(G20), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n615), .B(new_n616), .C1(new_n618), .C2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n613), .B1(new_n621), .B2(new_n256), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n585), .A2(new_n612), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n609), .A2(new_n611), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n607), .A2(G200), .A3(new_n608), .ZN(new_n626));
  OAI21_X1  g0426(.A(G190), .B1(new_n610), .B2(new_n606), .ZN(new_n627));
  INV_X1    g0427(.A(G87), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n473), .A2(new_n628), .ZN(new_n629));
  AOI211_X1 g0429(.A(new_n613), .B(new_n629), .C1(new_n621), .C2(new_n256), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n626), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n597), .A2(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n451), .A2(new_n507), .A3(new_n564), .A4(new_n633), .ZN(G372));
  NAND2_X1  g0434(.A1(new_n561), .A2(new_n562), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n531), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT92), .ZN(new_n637));
  INV_X1    g0437(.A(new_n496), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT92), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n563), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n602), .A2(new_n605), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n573), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n611), .A2(new_n624), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(G200), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n627), .A2(new_n630), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT91), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n644), .A2(new_n646), .A3(KEYINPUT91), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n548), .A2(new_n555), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n649), .A2(new_n650), .B1(new_n651), .B2(new_n558), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n641), .A2(new_n597), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n644), .A2(new_n646), .A3(KEYINPUT91), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT91), .B1(new_n644), .B2(new_n646), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n654), .B(new_n588), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n644), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n625), .A2(new_n631), .A3(new_n588), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(KEYINPUT26), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n451), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n308), .A2(new_n309), .ZN(new_n664));
  INV_X1    g0464(.A(new_n302), .ZN(new_n665));
  INV_X1    g0465(.A(new_n369), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n442), .B1(new_n667), .B2(new_n447), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n333), .A2(new_n337), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n328), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n670), .ZN(G369));
  AND2_X1   g0471(.A1(new_n212), .A2(G13), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n211), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n531), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n564), .A2(new_n679), .B1(new_n563), .B2(new_n678), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT93), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT93), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n678), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n638), .A2(new_n488), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n492), .A2(new_n678), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n685), .B1(new_n507), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n638), .A2(new_n678), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n637), .A2(new_n640), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(new_n678), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n223), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n618), .A2(new_n474), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(G1), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n228), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n701), .B1(new_n702), .B2(new_n698), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT28), .Z(new_n704));
  AOI211_X1 g0504(.A(KEYINPUT29), .B(new_n678), .C1(new_n653), .C2(new_n661), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT29), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n636), .A2(new_n638), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n652), .A2(KEYINPUT95), .A3(new_n597), .A4(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT95), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n559), .A2(new_n560), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n710), .A2(new_n552), .B1(new_n547), .B2(new_n331), .ZN(new_n711));
  OAI22_X1  g0511(.A1(new_n655), .A2(new_n656), .B1(new_n711), .B2(new_n531), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n597), .B1(new_n563), .B2(new_n496), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n644), .B1(new_n659), .B2(KEYINPUT26), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n588), .B1(new_n655), .B2(new_n656), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(KEYINPUT26), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n708), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n706), .B1(new_n718), .B2(new_n684), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n705), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT94), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  INV_X1    g0522(.A(new_n572), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n723), .B(new_n494), .C1(new_n606), .C2(new_n610), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n544), .A2(new_n546), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n721), .B(new_n722), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n468), .A2(new_n367), .A3(new_n642), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n547), .A2(new_n572), .A3(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n724), .A2(new_n725), .A3(new_n722), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n730), .B1(new_n731), .B2(KEYINPUT94), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n684), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n633), .A2(new_n564), .A3(new_n507), .A4(new_n684), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(KEYINPUT31), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n730), .A2(new_n728), .ZN(new_n737));
  INV_X1    g0537(.A(new_n731), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n736), .B(new_n684), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n720), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n704), .B1(new_n742), .B2(new_n211), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT96), .ZN(G364));
  AOI21_X1  g0544(.A(new_n211), .B1(new_n672), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n697), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n689), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n687), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(G330), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n223), .A2(new_n272), .ZN(new_n751));
  INV_X1    g0551(.A(G355), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n751), .A2(new_n752), .B1(G116), .B2(new_n223), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n696), .A2(new_n272), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G45), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(new_n228), .B2(new_n756), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n241), .A2(new_n756), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n753), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n226), .B1(G20), .B2(new_n573), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n747), .B1(new_n759), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT97), .Z(new_n768));
  NAND2_X1  g0568(.A1(new_n552), .A2(G20), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n367), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n212), .A2(new_n552), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n771), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n773), .A2(G311), .B1(new_n776), .B2(G322), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n367), .A2(new_n331), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n770), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n331), .A2(G179), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n774), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n780), .A2(new_n781), .B1(new_n784), .B2(G303), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n777), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n778), .A2(new_n774), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n272), .B(new_n786), .C1(G326), .C2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(KEYINPUT98), .B1(G179), .B2(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(KEYINPUT98), .A2(G179), .A3(G200), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n770), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT99), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(new_n792), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n552), .B1(new_n800), .B2(new_n790), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n212), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G294), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n770), .A2(new_n782), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT100), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G283), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n789), .A2(new_n799), .A3(new_n804), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n798), .A2(G159), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT32), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n806), .A2(new_n514), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n783), .A2(new_n628), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n772), .A2(new_n253), .B1(new_n775), .B2(new_n201), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(G50), .C2(new_n788), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n803), .A2(G97), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n385), .B1(new_n780), .B2(G68), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n813), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n809), .B1(new_n811), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n768), .B1(new_n820), .B2(new_n764), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n749), .B2(new_n763), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n750), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  INV_X1    g0624(.A(KEYINPUT102), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n678), .A2(new_n356), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n369), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n362), .A2(new_n369), .A3(new_n826), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n662), .A2(new_n684), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n678), .B1(new_n653), .B2(new_n661), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n829), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n741), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n741), .A2(new_n832), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n825), .B(new_n830), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n834), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n830), .A2(new_n825), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n741), .A2(new_n832), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n747), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n835), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n798), .A2(G311), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n272), .B1(new_n784), .B2(G107), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(KEYINPUT101), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n807), .B2(G87), .ZN(new_n845));
  INV_X1    g0645(.A(G283), .ZN(new_n846));
  INV_X1    g0646(.A(G294), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n779), .A2(new_n846), .B1(new_n775), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G303), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n772), .A2(new_n474), .B1(new_n787), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n848), .B(new_n850), .C1(KEYINPUT101), .C2(new_n843), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n842), .A2(new_n845), .A3(new_n817), .A4(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n780), .A2(G150), .B1(new_n776), .B2(G143), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  INV_X1    g0654(.A(G159), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n853), .B1(new_n854), .B2(new_n787), .C1(new_n855), .C2(new_n772), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT34), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n806), .A2(new_n202), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n385), .B(new_n858), .C1(G50), .C2(new_n784), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n859), .C1(new_n201), .C2(new_n802), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n797), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n852), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n764), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n764), .A2(new_n760), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n840), .B1(new_n253), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n864), .B(new_n866), .C1(new_n761), .C2(new_n829), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n841), .A2(new_n867), .ZN(G384));
  AND2_X1   g0668(.A1(new_n733), .A2(KEYINPUT31), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n735), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n436), .A2(new_n256), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n393), .A2(KEYINPUT16), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n438), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT103), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n676), .ZN(new_n877));
  OAI211_X1 g0677(.A(KEYINPUT103), .B(new_n438), .C1(new_n872), .C2(new_n873), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n425), .B2(new_n442), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n430), .B1(new_n427), .B2(new_n428), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n676), .B1(new_n882), .B2(new_n426), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n876), .A2(new_n883), .A3(new_n878), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n398), .A2(new_n419), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n432), .A2(new_n439), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n439), .A2(new_n877), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n885), .A2(new_n887), .A3(new_n888), .A4(new_n881), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n871), .B1(new_n880), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n884), .A2(new_n885), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n889), .B1(new_n893), .B2(new_n881), .ZN(new_n894));
  INV_X1    g0694(.A(new_n879), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n447), .B2(new_n448), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n896), .A3(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n308), .A2(new_n309), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n899), .B(new_n665), .C1(new_n271), .C2(new_n684), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n664), .A2(new_n678), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n900), .A2(new_n901), .B1(new_n828), .B2(new_n827), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n870), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n439), .B(new_n877), .C1(new_n447), .C2(new_n448), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n889), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n871), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n897), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n870), .A2(new_n912), .A3(KEYINPUT40), .A4(new_n902), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n905), .A2(new_n451), .A3(new_n870), .A4(new_n913), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n905), .A2(G330), .A3(new_n913), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n451), .B(G330), .C1(new_n735), .C2(new_n869), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n451), .B1(new_n705), .B2(new_n719), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n670), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n899), .A2(new_n678), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n911), .A2(new_n923), .A3(new_n897), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n923), .B1(new_n892), .B2(new_n897), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT104), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI211_X1 g0727(.A(KEYINPUT104), .B(new_n923), .C1(new_n892), .C2(new_n897), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n442), .A2(new_n877), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n900), .A2(new_n901), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n369), .A2(new_n678), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n931), .B1(new_n830), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n930), .B1(new_n934), .B2(new_n898), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n921), .A2(new_n936), .B1(new_n211), .B2(new_n672), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n921), .ZN(new_n938));
  INV_X1    g0738(.A(new_n580), .ZN(new_n939));
  OAI211_X1 g0739(.A(G116), .B(new_n227), .C1(new_n939), .C2(KEYINPUT35), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(KEYINPUT35), .B2(new_n939), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT36), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n228), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n207), .A2(G68), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n211), .B(G13), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n938), .A2(new_n942), .A3(new_n945), .ZN(G367));
  OR2_X1    g0746(.A1(new_n692), .A2(new_n713), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT42), .ZN(new_n948));
  INV_X1    g0748(.A(new_n588), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n597), .B1(new_n593), .B2(new_n684), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n636), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n947), .A2(KEYINPUT42), .B1(new_n684), .B2(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n655), .A2(new_n656), .B1(new_n630), .B2(new_n684), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n644), .A2(new_n630), .A3(new_n684), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n948), .A2(new_n952), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n588), .A2(new_n678), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n950), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n690), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT43), .ZN(new_n962));
  INV_X1    g0762(.A(new_n955), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n948), .A2(new_n952), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n957), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n961), .B1(new_n957), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n692), .A2(new_n694), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n960), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n969), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n968), .A2(new_n960), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n690), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n689), .A2(new_n691), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n683), .B(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n742), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n697), .B(KEYINPUT41), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n745), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n967), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(G317), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n797), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n385), .B1(new_n772), .B2(new_n846), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n805), .A2(new_n477), .B1(new_n775), .B2(new_n849), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(G311), .C2(new_n788), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT107), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n784), .A2(KEYINPUT46), .A3(G116), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n783), .B2(new_n474), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(new_n847), .C2(new_n779), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n988), .B1(new_n989), .B2(new_n993), .C1(new_n343), .C2(new_n802), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n985), .B(new_n994), .C1(new_n989), .C2(new_n993), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n779), .A2(new_n855), .B1(new_n772), .B2(new_n207), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n272), .B1(new_n805), .B2(new_n253), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n996), .A2(KEYINPUT108), .B1(new_n997), .B2(KEYINPUT109), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(KEYINPUT108), .B2(new_n996), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n803), .A2(G68), .ZN(new_n1000));
  INV_X1    g0800(.A(G150), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n201), .A2(new_n783), .B1(new_n775), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G143), .B2(new_n788), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1000), .B(new_n1003), .C1(KEYINPUT109), .C2(new_n997), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n999), .B(new_n1004), .C1(G137), .C2(new_n798), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n995), .A2(new_n1005), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT47), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(KEYINPUT47), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n764), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n755), .A2(new_n237), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n763), .B(new_n765), .C1(new_n223), .C2(new_n347), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1009), .B(new_n747), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT110), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n955), .B2(new_n763), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n983), .A2(new_n1014), .ZN(G387));
  OAI21_X1  g0815(.A(new_n754), .B1(new_n234), .B2(new_n756), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n700), .B2(new_n751), .ZN(new_n1017));
  AOI21_X1  g0817(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1018));
  OR3_X1    g0818(.A1(new_n321), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1019));
  OAI21_X1  g0819(.A(KEYINPUT50), .B1(new_n321), .B2(G50), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n700), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1017), .A2(new_n1021), .B1(new_n514), .B2(new_n696), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n747), .B1(new_n1022), .B2(new_n766), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G303), .A2(new_n773), .B1(new_n788), .B2(G322), .ZN(new_n1024));
  INV_X1    g0824(.A(G311), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n779), .C1(new_n984), .C2(new_n775), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT112), .Z(new_n1027));
  AND2_X1   g0827(.A1(new_n1027), .A2(KEYINPUT48), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(KEYINPUT48), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n802), .A2(new_n846), .B1(new_n847), .B2(new_n783), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n385), .B1(new_n805), .B2(new_n474), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n798), .B2(G326), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n797), .A2(new_n1001), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G159), .A2(new_n788), .B1(new_n776), .B2(G50), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n784), .A2(G77), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n272), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G97), .B2(new_n807), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n803), .A2(new_n612), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n321), .A2(new_n779), .B1(new_n772), .B2(new_n202), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT111), .Z(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1036), .B1(new_n1037), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1023), .B1(new_n1046), .B2(new_n764), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n681), .A2(new_n682), .A3(new_n762), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n746), .A2(new_n978), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n742), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n978), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n697), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1050), .A2(new_n978), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(G393));
  INV_X1    g0854(.A(new_n690), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n969), .B(new_n970), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n973), .B(KEYINPUT44), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n976), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n1051), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n976), .A2(new_n1050), .A3(new_n978), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n697), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1058), .A2(new_n746), .A3(new_n976), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n272), .B1(new_n772), .B2(new_n321), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n779), .A2(new_n207), .B1(new_n783), .B2(new_n202), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n807), .C2(G87), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n798), .A2(G143), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n803), .A2(G77), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n787), .A2(new_n1001), .B1(new_n775), .B2(new_n855), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n272), .B(new_n812), .C1(G283), .C2(new_n784), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n773), .A2(G294), .B1(new_n780), .B2(G303), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n802), .B2(new_n474), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT113), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n798), .A2(G322), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n787), .A2(new_n984), .B1(new_n775), .B2(new_n1025), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT52), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1071), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n764), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n754), .A2(new_n244), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n766), .B1(G97), .B2(new_n696), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n840), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1083), .B(new_n1086), .C1(new_n959), .C2(new_n763), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1063), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1062), .A2(new_n1088), .ZN(G390));
  NAND3_X1  g0889(.A1(new_n919), .A2(new_n670), .A3(new_n916), .ZN(new_n1090));
  OAI211_X1 g0890(.A(G330), .B(new_n829), .C1(new_n735), .C2(new_n739), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n931), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n902), .B(G330), .C1(new_n735), .C2(new_n869), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n830), .A2(new_n933), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n931), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n740), .A2(G330), .A3(new_n829), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n718), .A2(new_n684), .A3(new_n829), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n933), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(G330), .B(new_n829), .C1(new_n735), .C2(new_n869), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n931), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1098), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1090), .B1(new_n1096), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT38), .B1(new_n906), .B2(new_n909), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n880), .A2(new_n891), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(KEYINPUT38), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(new_n922), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n1101), .B2(new_n931), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n880), .A2(new_n891), .A3(new_n871), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT38), .B1(new_n894), .B2(new_n896), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT39), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(KEYINPUT104), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n925), .A2(new_n926), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n1115), .A3(new_n924), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n922), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1110), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1093), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1098), .B(new_n1110), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1105), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n922), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n912), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n927), .A2(new_n928), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n932), .B1(new_n831), .B2(new_n829), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1123), .B1(new_n1127), .B2(new_n931), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1125), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1105), .B(new_n1121), .C1(new_n1129), .C2(new_n1093), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n697), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT114), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1122), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(KEYINPUT114), .A3(new_n697), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1121), .B(new_n746), .C1(new_n1129), .C2(new_n1093), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n840), .B1(new_n321), .B2(new_n865), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n272), .B1(new_n805), .B2(new_n207), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT115), .Z(new_n1139));
  NAND2_X1  g0939(.A1(new_n784), .A2(G150), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT53), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  INV_X1    g0942(.A(G128), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n772), .A2(new_n1142), .B1(new_n787), .B2(new_n1143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n779), .A2(new_n854), .B1(new_n775), .B2(new_n861), .ZN(new_n1145));
  NOR4_X1   g0945(.A1(new_n1139), .A2(new_n1141), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(G125), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n797), .C1(new_n855), .C2(new_n802), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n798), .A2(G294), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n858), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n779), .A2(new_n343), .B1(new_n787), .B2(new_n846), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n772), .A2(new_n477), .B1(new_n775), .B2(new_n474), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n272), .A4(new_n814), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1149), .A2(new_n1150), .A3(new_n1068), .A4(new_n1153), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1148), .A2(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1137), .B1(new_n765), .B2(new_n1155), .C1(new_n1116), .C2(new_n761), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1136), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT116), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT116), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1136), .A2(new_n1159), .A3(new_n1156), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1135), .A2(new_n1161), .ZN(G378));
  INV_X1    g0962(.A(new_n915), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n338), .A2(KEYINPUT119), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n338), .A2(KEYINPUT119), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n326), .A2(new_n676), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1166), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1169), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n929), .A2(new_n935), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n929), .B2(new_n935), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1163), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1113), .A2(KEYINPUT104), .B1(new_n1108), .B2(new_n923), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1123), .B1(new_n1178), .B2(new_n1115), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n934), .A2(new_n898), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n930), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1173), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n929), .A2(new_n935), .A3(new_n1174), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n915), .A3(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1177), .A2(new_n1185), .A3(new_n746), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n840), .B1(new_n207), .B2(new_n865), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n805), .A2(new_n201), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n272), .A2(G41), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1039), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT117), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1188), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n1191), .B2(new_n1190), .C1(new_n797), .C2(new_n846), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT118), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n780), .A2(G97), .B1(new_n788), .B2(G116), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n773), .A2(new_n612), .B1(new_n776), .B2(G107), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1194), .A2(new_n1000), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(G33), .A2(G41), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1189), .A2(G50), .A3(new_n1200), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n779), .A2(new_n861), .B1(new_n783), .B2(new_n1142), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n773), .A2(G137), .B1(new_n776), .B2(G128), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1147), .B2(new_n787), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(G150), .C2(new_n803), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  INV_X1    g1007(.A(G124), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1200), .B1(new_n855), .B2(new_n805), .C1(new_n797), .C2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1206), .B2(KEYINPUT59), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1201), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1199), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1198), .B2(new_n1197), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1187), .B1(new_n765), .B2(new_n1213), .C1(new_n1173), .C2(new_n761), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1186), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1090), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1130), .A2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1218), .A2(KEYINPUT57), .A3(new_n1185), .A4(new_n1177), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n697), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1177), .A2(new_n1185), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1221), .B2(new_n1218), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1216), .B1(new_n1220), .B2(new_n1222), .ZN(G375));
  INV_X1    g1023(.A(new_n1105), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1096), .A2(new_n1090), .A3(new_n1104), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n980), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1096), .A2(new_n1104), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n746), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G294), .A2(new_n788), .B1(new_n784), .B2(G97), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n474), .B2(new_n779), .C1(new_n846), .C2(new_n775), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n272), .B(new_n1230), .C1(new_n617), .C2(new_n773), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n807), .A2(G77), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1042), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G303), .B2(new_n798), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1188), .A2(new_n385), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT120), .Z(new_n1236));
  OAI22_X1  g1036(.A1(new_n772), .A2(new_n1001), .B1(new_n783), .B2(new_n855), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n779), .A2(new_n1142), .B1(new_n787), .B2(new_n861), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(G137), .C2(new_n776), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1236), .B(new_n1239), .C1(new_n207), .C2(new_n802), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G128), .B2(new_n798), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n764), .B1(new_n1234), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n840), .B1(new_n202), .B2(new_n865), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(new_n1097), .C2(new_n761), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1226), .A2(new_n1228), .A3(new_n1244), .ZN(G381));
  OR2_X1    g1045(.A1(G393), .A2(G396), .ZN(new_n1246));
  OR4_X1    g1046(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT57), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1130), .A2(new_n1217), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1177), .A2(new_n1185), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(new_n697), .A3(new_n1219), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1133), .A2(new_n1134), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1216), .ZN(new_n1254));
  OR3_X1    g1054(.A1(new_n1247), .A2(G387), .A3(new_n1254), .ZN(G407));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G343), .C2(new_n1254), .ZN(G409));
  XNOR2_X1  g1056(.A(G393), .B(new_n823), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1062), .A2(new_n1088), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1258), .B1(new_n1062), .B2(new_n1088), .ZN(new_n1261));
  OAI21_X1  g1061(.A(G387), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G390), .A2(new_n1257), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1014), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n967), .B2(new_n982), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1265), .A3(new_n1259), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n677), .A2(G213), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G375), .A2(G378), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1186), .A2(KEYINPUT121), .A3(new_n1214), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1221), .A2(new_n980), .A3(new_n1218), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT121), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1215), .A2(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1253), .A2(new_n1271), .A3(new_n1272), .A4(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1270), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT122), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1269), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1270), .A2(KEYINPUT122), .A3(new_n1275), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT123), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G384), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n841), .A2(KEYINPUT123), .A3(new_n867), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1282), .A2(new_n1228), .A3(new_n1244), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT60), .ZN(new_n1284));
  OR2_X1    g1084(.A1(new_n1225), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1225), .A2(new_n1284), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n697), .A3(new_n1224), .A4(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1281), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1283), .A2(new_n1287), .A3(new_n1281), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1278), .B(new_n1279), .C1(new_n1288), .C2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1269), .A2(G2897), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT124), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1269), .A2(KEYINPUT124), .A3(G2897), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1296), .B(new_n1297), .C1(new_n1290), .C2(new_n1288), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1288), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1299), .A2(new_n1295), .A3(new_n1289), .A4(new_n1294), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1276), .B2(new_n1269), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1290), .A2(new_n1288), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1276), .A2(new_n1303), .A3(new_n1269), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1293), .B(new_n1302), .C1(new_n1304), .C2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1267), .B1(new_n1292), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1301), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1291), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1262), .A2(new_n1266), .A3(new_n1293), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1304), .B2(KEYINPUT63), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT125), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1274), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1315), .A2(G378), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1253), .B1(new_n1252), .B2(new_n1216), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1277), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(new_n1279), .A3(new_n1268), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1310), .B1(new_n1319), .B2(new_n1301), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1303), .ZN(new_n1321));
  OAI211_X1 g1121(.A(KEYINPUT125), .B(new_n1313), .C1(new_n1320), .C2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1307), .B1(new_n1314), .B2(new_n1323), .ZN(G405));
  NAND2_X1  g1124(.A1(new_n1270), .A2(new_n1254), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1325), .A2(new_n1303), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT126), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1326), .B(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1325), .A2(new_n1303), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1329), .B(KEYINPUT127), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(new_n1267), .ZN(G402));
endmodule


