//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n547, new_n549, new_n550, new_n551, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT65), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n462), .A2(new_n470), .A3(G137), .A4(new_n464), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n462), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT66), .Z(new_n477));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  MUX2_X1   g055(.A(G100), .B(G112), .S(G2105), .Z(new_n481));
  AOI22_X1  g056(.A1(G136), .A2(new_n480), .B1(new_n481), .B2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(KEYINPUT67), .A2(KEYINPUT4), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT67), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n480), .B2(G138), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(new_n486), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n485), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(G114), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G102), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n474), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT68), .B1(new_n491), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n485), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n489), .A2(new_n486), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n462), .A2(G138), .A3(new_n464), .A4(new_n487), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n503), .A2(new_n504), .A3(new_n497), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n499), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n507), .A2(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n515), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT69), .B(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n511), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n512), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n510), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n524), .A2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n517), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n533), .A2(new_n511), .B1(new_n513), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(KEYINPUT70), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(KEYINPUT70), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n540), .A2(new_n511), .B1(new_n513), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n517), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT71), .Z(G188));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n554), .B(new_n555), .C1(new_n511), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n508), .A2(new_n509), .ZN(new_n558));
  INV_X1    g133(.A(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n560), .A2(new_n553), .A3(KEYINPUT9), .A4(G53), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n525), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n525), .A2(new_n558), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n566), .A2(G651), .B1(new_n567), .B2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(G299));
  NAND2_X1  g144(.A1(new_n560), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n513), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(KEYINPUT73), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(KEYINPUT73), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G288));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n578), .A2(new_n511), .B1(new_n513), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n517), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G60), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n525), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n517), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(new_n588), .B2(new_n587), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n567), .A2(G85), .B1(new_n560), .B2(G47), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n525), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n560), .B2(G54), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(KEYINPUT75), .B(KEYINPUT10), .Z(new_n599));
  OR3_X1    g174(.A1(new_n513), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n513), .B2(new_n598), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g179(.A(new_n603), .B1(G171), .B2(G868), .ZN(G321));
  MUX2_X1   g180(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g181(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g182(.A(new_n602), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT76), .B(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(G860), .B2(new_n609), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT77), .Z(G148));
  INV_X1    g186(.A(new_n545), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n609), .ZN(new_n613));
  MUX2_X1   g188(.A(new_n612), .B(new_n613), .S(G868), .Z(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n480), .A2(G2104), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  MUX2_X1   g196(.A(G99), .B(G111), .S(G2105), .Z(new_n622));
  AOI22_X1  g197(.A1(new_n475), .A2(G123), .B1(G2104), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G135), .ZN(new_n624));
  INV_X1    g199(.A(new_n480), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND3_X1  g202(.A1(new_n620), .A2(new_n621), .A3(new_n627), .ZN(G156));
  INV_X1    g203(.A(G14), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2427), .ZN(new_n632));
  INV_X1    g207(.A(G2430), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n636), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT78), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT79), .Z(new_n645));
  AOI211_X1 g220(.A(new_n629), .B(new_n645), .C1(new_n643), .C2(new_n641), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT18), .ZN(new_n653));
  INV_X1    g228(.A(new_n649), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n650), .B1(new_n656), .B2(new_n647), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n648), .B2(new_n655), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n648), .A2(new_n651), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n654), .B1(new_n659), .B2(KEYINPUT17), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n653), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2096), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT80), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n666), .A2(new_n669), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT20), .Z(new_n673));
  AOI211_X1 g248(.A(new_n671), .B(new_n673), .C1(new_n666), .C2(new_n670), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT81), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(G229));
  NOR2_X1   g256(.A1(G16), .A2(G24), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n592), .B2(G16), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT83), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1986), .ZN(new_n685));
  MUX2_X1   g260(.A(G95), .B(G107), .S(G2105), .Z(new_n686));
  AOI22_X1  g261(.A1(new_n475), .A2(G119), .B1(G2104), .B2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G131), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n625), .ZN(new_n689));
  MUX2_X1   g264(.A(G25), .B(new_n689), .S(G29), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT82), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT35), .B(G1991), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT84), .Z(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G303), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT85), .B(G1971), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G23), .B(new_n573), .S(G16), .Z(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT33), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(G6), .A2(G16), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n583), .B2(G16), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n700), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n685), .B(new_n694), .C1(KEYINPUT34), .C2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT86), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(KEYINPUT34), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT36), .Z(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G32), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT26), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n475), .A2(G129), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n480), .A2(G141), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n717), .B(new_n720), .C1(G105), .C2(new_n460), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n715), .B1(new_n721), .B2(new_n714), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT27), .B(G1996), .Z(new_n723));
  INV_X1    g298(.A(G2084), .ZN(new_n724));
  AND2_X1   g299(.A1(KEYINPUT24), .A2(G34), .ZN(new_n725));
  NOR2_X1   g300(.A1(KEYINPUT24), .A2(G34), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n714), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G160), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n714), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n722), .A2(new_n723), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G2072), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n714), .A2(G33), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n462), .A2(G127), .ZN(new_n733));
  AND2_X1   g308(.A1(G115), .A2(G2104), .ZN(new_n734));
  OAI21_X1  g309(.A(G2105), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT25), .ZN(new_n739));
  INV_X1    g314(.A(new_n460), .ZN(new_n740));
  INV_X1    g315(.A(G103), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n460), .A2(KEYINPUT25), .A3(G103), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n742), .A2(new_n743), .B1(G139), .B2(new_n480), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n737), .A2(new_n738), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n732), .B1(new_n745), .B2(G29), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n730), .B1(new_n731), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n731), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT89), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT90), .Z(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G35), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G162), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT29), .Z(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT92), .Z(new_n757));
  NOR2_X1   g332(.A1(new_n754), .A2(new_n755), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n714), .A2(G26), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT28), .Z(new_n760));
  MUX2_X1   g335(.A(G104), .B(G116), .S(G2105), .Z(new_n761));
  AOI22_X1  g336(.A1(new_n475), .A2(G128), .B1(G2104), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G140), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n625), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n760), .B1(new_n764), .B2(G29), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT87), .B(G2067), .Z(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT31), .B(G11), .Z(new_n768));
  INV_X1    g343(.A(G28), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(KEYINPUT30), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT91), .Z(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n769), .B2(KEYINPUT30), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n768), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n773), .B1(new_n714), .B2(new_n626), .C1(new_n765), .C2(new_n766), .ZN(new_n774));
  INV_X1    g349(.A(G1341), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n545), .A2(G16), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G16), .B2(G19), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n767), .B(new_n774), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n775), .ZN(new_n779));
  NOR2_X1   g354(.A1(G168), .A2(new_n695), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n695), .B2(G21), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n779), .B1(new_n782), .B2(G1966), .ZN(new_n783));
  INV_X1    g358(.A(G1966), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n781), .A2(new_n784), .B1(new_n722), .B2(new_n723), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n778), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n729), .A2(new_n724), .ZN(new_n787));
  NOR2_X1   g362(.A1(G4), .A2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n608), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1348), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n758), .A2(new_n786), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n695), .A2(G20), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT93), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT23), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G299), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1956), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n695), .A2(G5), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G171), .B2(new_n695), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n796), .B1(G1961), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G1961), .B2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n714), .A2(G27), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G164), .B2(new_n714), .ZN(new_n802));
  INV_X1    g377(.A(G2078), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n757), .A2(new_n791), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n713), .A2(new_n751), .A3(new_n805), .ZN(G311));
  INV_X1    g381(.A(G311), .ZN(G150));
  INV_X1    g382(.A(G55), .ZN(new_n808));
  INV_X1    g383(.A(G93), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n808), .A2(new_n511), .B1(new_n513), .B2(new_n809), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n517), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT96), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n612), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n545), .A2(new_n813), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n608), .A2(G559), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n822), .B(new_n823), .Z(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT94), .ZN(new_n826));
  AOI21_X1  g401(.A(G860), .B1(new_n824), .B2(KEYINPUT39), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n818), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT97), .Z(G145));
  XNOR2_X1  g404(.A(new_n689), .B(new_n617), .ZN(new_n830));
  MUX2_X1   g405(.A(G106), .B(G118), .S(G2105), .Z(new_n831));
  AOI22_X1  g406(.A1(new_n475), .A2(G130), .B1(G2104), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G142), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n625), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n830), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n491), .A2(new_n498), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n764), .B(new_n836), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n835), .B(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n721), .B(new_n745), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n483), .B(new_n626), .ZN(new_n841));
  XNOR2_X1  g416(.A(G160), .B(KEYINPUT98), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(G37), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n840), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT99), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(G395));
  NOR2_X1   g423(.A1(new_n814), .A2(G868), .ZN(new_n849));
  XNOR2_X1  g424(.A(G299), .B(new_n608), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT41), .Z(new_n851));
  XOR2_X1   g426(.A(new_n821), .B(new_n613), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n850), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT42), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n592), .B(new_n573), .ZN(new_n857));
  XNOR2_X1  g432(.A(G305), .B(G303), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n856), .B(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n849), .B1(new_n861), .B2(G868), .ZN(G331));
  XOR2_X1   g437(.A(G331), .B(KEYINPUT101), .Z(G295));
  XNOR2_X1  g438(.A(G301), .B(G168), .ZN(new_n864));
  INV_X1    g439(.A(new_n821), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(new_n854), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n866), .A2(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n867), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n869), .B1(new_n873), .B2(new_n851), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n860), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n874), .A2(new_n860), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n876), .A2(KEYINPUT103), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT103), .B1(new_n876), .B2(new_n877), .ZN(new_n879));
  OAI211_X1 g454(.A(KEYINPUT43), .B(new_n875), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n873), .A2(new_n854), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n851), .B2(new_n868), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n877), .B(new_n875), .C1(new_n883), .C2(new_n860), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n885), .B(new_n875), .C1(new_n878), .C2(new_n879), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n881), .B1(new_n884), .B2(KEYINPUT43), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n888), .A2(KEYINPUT104), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT104), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(G397));
  XNOR2_X1  g467(.A(KEYINPUT105), .B(G1384), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n836), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT45), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(G113), .A2(G2104), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n466), .A2(new_n467), .ZN(new_n898));
  INV_X1    g473(.A(G125), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n900), .A2(G2105), .B1(G101), .B2(new_n460), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n901), .A2(G40), .A3(new_n469), .A4(new_n471), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n764), .B(G2067), .Z(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n721), .B2(new_n905), .ZN(new_n906));
  OR3_X1    g481(.A1(new_n904), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT46), .B1(new_n904), .B2(G1996), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT47), .Z(new_n910));
  XNOR2_X1  g485(.A(new_n721), .B(G1996), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n911), .A2(new_n905), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n689), .A2(new_n693), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT125), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n764), .A2(G2067), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n904), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n689), .A2(new_n693), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(new_n918), .A3(new_n913), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n904), .A2(G1986), .A3(G290), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n919), .A2(new_n903), .B1(KEYINPUT48), .B2(new_n920), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n920), .A2(KEYINPUT48), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n910), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT126), .ZN(new_n925));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n503), .B2(new_n497), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n902), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G8), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT49), .ZN(new_n931));
  OAI21_X1  g506(.A(G1981), .B1(new_n580), .B2(new_n582), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n580), .A2(G1981), .A3(new_n582), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n934), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n932), .A3(KEYINPUT49), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n930), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1976), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n938), .A2(new_n939), .A3(new_n576), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n930), .B1(new_n940), .B2(new_n934), .ZN(new_n941));
  INV_X1    g516(.A(G40), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n465), .A2(new_n472), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n836), .A3(new_n926), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n944), .B(G8), .C1(new_n939), .C2(new_n573), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n576), .B2(G1976), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n938), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n945), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT107), .B1(new_n949), .B2(new_n946), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n951), .A3(KEYINPUT52), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n948), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n955), .B(new_n926), .C1(new_n503), .C2(new_n497), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n956), .A2(new_n943), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n491), .A2(KEYINPUT68), .A3(new_n498), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n504), .B1(new_n503), .B2(new_n497), .ZN(new_n959));
  AOI21_X1  g534(.A(G1384), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n957), .B(new_n755), .C1(new_n960), .C2(new_n955), .ZN(new_n961));
  OAI211_X1 g536(.A(KEYINPUT45), .B(new_n893), .C1(new_n503), .C2(new_n497), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n943), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n926), .B1(new_n499), .B2(new_n505), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n895), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n961), .B1(new_n965), .B2(G1971), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(G303), .A2(G8), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT55), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n962), .A2(new_n943), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n960), .B2(KEYINPUT45), .ZN(new_n973));
  INV_X1    g548(.A(G1971), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(KEYINPUT106), .A3(new_n961), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n968), .A2(G8), .A3(new_n971), .A4(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n941), .B1(new_n954), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(G286), .A2(G8), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT116), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n957), .B(new_n724), .C1(new_n960), .C2(new_n955), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT45), .B(new_n926), .C1(new_n499), .C2(new_n505), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n902), .B1(new_n895), .B2(new_n927), .ZN(new_n984));
  AOI21_X1  g559(.A(G1966), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n980), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(G8), .B1(new_n982), .B2(new_n985), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT117), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n989), .B(G8), .C1(new_n982), .C2(new_n985), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n980), .A2(KEYINPUT51), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n988), .A2(KEYINPUT118), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n983), .A2(new_n984), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n784), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n929), .B1(new_n994), .B2(new_n981), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT51), .B1(new_n995), .B2(new_n980), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n980), .A2(KEYINPUT51), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n995), .B2(new_n989), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT118), .B1(new_n999), .B2(new_n988), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n986), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n972), .B(new_n803), .C1(new_n960), .C2(KEYINPUT45), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n983), .A2(KEYINPUT53), .A3(new_n803), .A4(new_n984), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n957), .B1(new_n960), .B2(new_n955), .ZN(new_n1006));
  INV_X1    g581(.A(G1961), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G171), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT120), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n896), .A2(new_n972), .A3(KEYINPUT53), .A4(new_n803), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1004), .A2(new_n1008), .A3(G301), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1009), .A2(new_n1016), .A3(G171), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1011), .A2(new_n1015), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT54), .B1(new_n1009), .B2(G171), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1004), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT122), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT122), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1004), .A2(new_n1008), .A3(new_n1025), .A4(new_n1012), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1022), .B1(new_n1027), .B2(G171), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n960), .A2(new_n955), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n902), .B1(KEYINPUT50), .B2(new_n927), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n755), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n929), .B1(new_n975), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT108), .B1(new_n1032), .B2(new_n971), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT108), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n927), .A2(KEYINPUT50), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n943), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n955), .B2(new_n960), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1037), .A2(new_n755), .B1(new_n973), .B2(new_n974), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1034), .B(new_n970), .C1(new_n1038), .C2(new_n929), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n977), .A2(new_n1033), .A3(new_n953), .A4(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1028), .A2(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1001), .A2(new_n1021), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT111), .B1(new_n1037), .B2(G1956), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n1045));
  INV_X1    g620(.A(G1956), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT56), .B(G2072), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT114), .B1(new_n965), .B2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n972), .B(new_n1048), .C1(new_n960), .C2(KEYINPUT45), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1043), .B(new_n1047), .C1(new_n1049), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1045), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1056));
  AOI211_X1 g631(.A(KEYINPUT111), .B(G1956), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1050), .B(new_n1051), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(KEYINPUT115), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n562), .A2(KEYINPUT112), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n568), .B1(new_n562), .B2(KEYINPUT112), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n563), .A2(KEYINPUT57), .A3(new_n568), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1058), .A2(new_n1069), .A3(new_n1059), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n944), .A2(G2067), .ZN(new_n1072));
  INV_X1    g647(.A(G1348), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1006), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(new_n602), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1061), .A2(new_n1070), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT61), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1053), .A2(new_n1070), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1069), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT58), .B(G1341), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n973), .A2(G1996), .B1(new_n928), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n545), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT59), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1085), .A3(new_n545), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n608), .B(new_n1072), .C1(new_n1006), .C2(new_n1073), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT60), .B1(new_n1075), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT60), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1074), .A2(new_n1090), .A3(new_n608), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1080), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1071), .A2(KEYINPUT61), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1061), .B2(new_n1070), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1076), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n978), .B1(new_n1042), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n990), .A2(new_n991), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n995), .A2(new_n989), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(new_n992), .A3(new_n996), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1098), .B1(new_n1103), .B2(new_n986), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1098), .A3(new_n986), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1040), .B1(new_n1017), .B2(new_n1011), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1105), .A2(KEYINPUT123), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n1104), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n995), .A2(G168), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT109), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT63), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n954), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n968), .A2(G8), .A3(new_n976), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n970), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1113), .A2(new_n1115), .A3(new_n977), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1040), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(KEYINPUT110), .A3(new_n1113), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1114), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT110), .B1(new_n1119), .B2(new_n1113), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1097), .A2(new_n1108), .A3(new_n1111), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n1125));
  XOR2_X1   g700(.A(new_n592), .B(G1986), .Z(new_n1126));
  OAI21_X1  g701(.A(new_n903), .B1(new_n919), .B2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1125), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n925), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT127), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT127), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1132), .B(new_n925), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g709(.A(G319), .ZN(new_n1136));
  NOR4_X1   g710(.A1(G401), .A2(G229), .A3(new_n1136), .A4(G227), .ZN(new_n1137));
  NAND4_X1  g711(.A1(new_n1137), .A2(new_n880), .A3(new_n846), .A4(new_n886), .ZN(G225));
  INV_X1    g712(.A(G225), .ZN(G308));
endmodule


