//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1337, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n207), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT66), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n207), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n226), .B(new_n233), .C1(KEYINPUT1), .C2(new_n220), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n222), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G58), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(new_n209), .ZN(new_n253));
  OAI21_X1  g0053(.A(G20), .B1(new_n253), .B2(new_n201), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G159), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT7), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n260), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(KEYINPUT76), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n263), .B2(new_n231), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT76), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT76), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(new_n265), .A3(G33), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n268), .A2(new_n259), .A3(new_n231), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G68), .ZN(new_n272));
  OAI211_X1 g0072(.A(KEYINPUT16), .B(new_n258), .C1(new_n264), .C2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT16), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n259), .B1(new_n262), .B2(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n266), .A2(new_n267), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n209), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n274), .B1(new_n278), .B2(new_n257), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n230), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n273), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  XOR2_X1   g0082(.A(KEYINPUT8), .B(G58), .Z(new_n283));
  INV_X1    g0083(.A(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G20), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G13), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(new_n231), .A3(G1), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n281), .ZN(new_n289));
  INV_X1    g0089(.A(new_n283), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n286), .A2(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n282), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  AND2_X1   g0093(.A1(G1), .A2(G13), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G41), .ZN(new_n297));
  INV_X1    g0097(.A(G45), .ZN(new_n298));
  AOI21_X1  g0098(.A(G1), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(new_n295), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n284), .B1(G41), .B2(G45), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(G232), .A3(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n260), .A2(new_n211), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n268), .A2(new_n270), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G223), .A2(G1698), .ZN(new_n307));
  INV_X1    g0107(.A(G226), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(G1698), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n305), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n304), .B1(new_n310), .B2(new_n301), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G169), .ZN(new_n312));
  OAI211_X1 g0112(.A(G179), .B(new_n304), .C1(new_n310), .C2(new_n301), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n292), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT18), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT18), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n292), .A2(new_n317), .A3(new_n314), .ZN(new_n318));
  INV_X1    g0118(.A(G190), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n319), .B(new_n304), .C1(new_n310), .C2(new_n301), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n300), .A2(new_n303), .ZN(new_n321));
  INV_X1    g0121(.A(new_n305), .ZN(new_n322));
  INV_X1    g0122(.A(new_n309), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n263), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n301), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n320), .B1(new_n326), .B2(G200), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n282), .A2(new_n327), .A3(new_n291), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT17), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n282), .A2(new_n327), .A3(KEYINPUT17), .A4(new_n291), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n316), .A2(new_n318), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  INV_X1    g0133(.A(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n308), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n334), .A2(G232), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n262), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n325), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n301), .A2(G238), .A3(new_n302), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n300), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n301), .B1(new_n337), .B2(new_n338), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT13), .B1(new_n346), .B2(new_n342), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n333), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n347), .ZN(new_n350));
  INV_X1    g0150(.A(G179), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n348), .A2(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(G169), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT75), .B1(new_n353), .B2(KEYINPUT14), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT75), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n348), .A2(new_n355), .A3(new_n349), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n352), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n260), .A2(G20), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(G77), .B1(G20), .B2(new_n209), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n231), .A2(new_n260), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n202), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n281), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT11), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT74), .B1(new_n288), .B2(new_n209), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT12), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n289), .A2(G68), .A3(new_n285), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n362), .B2(new_n363), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n357), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n350), .A2(G200), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n370), .C1(new_n319), .C2(new_n350), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n289), .A2(G50), .A3(new_n285), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n287), .A2(G1), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G20), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n375), .B1(G50), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n281), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n283), .A2(new_n358), .B1(G150), .B2(new_n255), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n203), .A2(G20), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g0183(.A(new_n383), .B(KEYINPUT9), .Z(new_n384));
  NAND2_X1  g0184(.A1(new_n301), .A2(new_n302), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n300), .B1(new_n385), .B2(new_n308), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G222), .A2(G1698), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n334), .A2(G223), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n262), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n301), .B1(new_n276), .B2(new_n215), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n319), .ZN(new_n392));
  XOR2_X1   g0192(.A(KEYINPUT71), .B(G200), .Z(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n392), .B1(new_n394), .B2(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n384), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT10), .B1(new_n395), .B2(KEYINPUT73), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n397), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n391), .A2(G169), .ZN(new_n400));
  AOI211_X1 g0200(.A(new_n383), .B(new_n400), .C1(new_n351), .C2(new_n391), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n301), .A2(G244), .A3(new_n302), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n300), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n262), .A2(G238), .A3(G1698), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n262), .A2(G232), .A3(new_n334), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT68), .B(G107), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n406), .B(new_n407), .C1(new_n262), .C2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n405), .B1(new_n410), .B2(new_n325), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n411), .A2(G169), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT15), .B(G87), .Z(new_n413));
  INV_X1    g0213(.A(KEYINPUT70), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT15), .B(G87), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT70), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n415), .A2(new_n358), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n360), .A2(KEYINPUT69), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT69), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n255), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n283), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G20), .A2(G77), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n281), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n288), .A2(new_n215), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n289), .A2(G77), .A3(new_n285), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n412), .A2(new_n428), .A3(KEYINPUT72), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n422), .A2(new_n423), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n415), .A2(new_n358), .A3(new_n417), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n379), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n426), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n432), .A2(new_n433), .B1(new_n411), .B2(G169), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT72), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n411), .A2(new_n351), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n429), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n432), .A2(new_n433), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n411), .A2(G190), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(new_n393), .C2(new_n411), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  OR4_X1    g0242(.A1(new_n332), .A2(new_n374), .A3(new_n403), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n210), .A2(new_n334), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n216), .A2(G1698), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n306), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G116), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n301), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n284), .A2(new_n293), .A3(G45), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n212), .B1(new_n298), .B2(G1), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n301), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT83), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n301), .A2(new_n455), .A3(new_n451), .A4(new_n452), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n394), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n306), .A2(new_n231), .A3(G68), .ZN(new_n459));
  OR2_X1    g0259(.A1(KEYINPUT68), .A2(G107), .ZN(new_n460));
  INV_X1    g0260(.A(G97), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT68), .A2(G107), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n460), .A2(new_n211), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT19), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n231), .B1(new_n338), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n358), .A2(G97), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n463), .A2(new_n465), .B1(new_n466), .B2(new_n464), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n415), .A2(new_n417), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n468), .A2(new_n281), .B1(new_n288), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n457), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n446), .B1(new_n268), .B2(new_n270), .ZN(new_n472));
  INV_X1    g0272(.A(new_n449), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n325), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(G190), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n284), .A2(G33), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n379), .A2(new_n377), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G87), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n458), .A2(new_n470), .A3(new_n475), .A4(new_n478), .ZN(new_n479));
  AOI211_X1 g0279(.A(G20), .B(new_n209), .C1(new_n268), .C2(new_n270), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n211), .A2(new_n461), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n465), .B1(new_n408), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n466), .A2(new_n464), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n281), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n415), .A2(new_n417), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n477), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n469), .A2(new_n288), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n333), .B1(new_n450), .B2(new_n457), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n471), .A2(new_n351), .A3(new_n474), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n479), .A2(new_n492), .A3(KEYINPUT84), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT84), .B1(new_n479), .B2(new_n492), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(KEYINPUT4), .A2(G244), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n266), .A2(new_n267), .A3(new_n496), .A4(new_n334), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n216), .A2(G1698), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n306), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n266), .A2(new_n267), .A3(G250), .A4(G1698), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT78), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT78), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n262), .A2(new_n506), .A3(G250), .A4(G1698), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT79), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n500), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n502), .B1(new_n263), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n497), .A2(new_n498), .ZN(new_n512));
  AND4_X1   g0312(.A1(KEYINPUT79), .A2(new_n511), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n325), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n284), .B(G45), .C1(new_n297), .C2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT80), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G41), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(KEYINPUT80), .A3(new_n284), .A4(G45), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n518), .A2(G41), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n517), .A2(new_n520), .A3(new_n296), .A4(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT81), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n515), .B2(new_n516), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n526), .A2(KEYINPUT81), .A3(new_n296), .A4(new_n520), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n325), .B1(new_n526), .B2(new_n520), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G257), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n514), .A2(new_n351), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT79), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n510), .B1(new_n268), .B2(new_n270), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n512), .B1(new_n535), .B2(KEYINPUT4), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n505), .A2(new_n507), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n511), .A2(KEYINPUT79), .A3(new_n508), .A4(new_n512), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n301), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n333), .B1(new_n540), .B2(new_n531), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n289), .A2(new_n476), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n377), .A2(new_n461), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT77), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(KEYINPUT77), .A3(new_n544), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n461), .A2(new_n217), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n552), .B2(KEYINPUT6), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n275), .A2(new_n277), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(new_n409), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n547), .A2(new_n548), .B1(new_n556), .B2(new_n281), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n533), .A2(new_n541), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(G200), .B1(new_n540), .B2(new_n531), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n538), .A2(new_n539), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n531), .B1(new_n561), .B2(new_n325), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n560), .A2(KEYINPUT82), .B1(new_n562), .B2(G190), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n514), .A2(KEYINPUT82), .A3(G190), .A4(new_n532), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n557), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n495), .B(new_n559), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  XNOR2_X1  g0366(.A(KEYINPUT87), .B(KEYINPUT22), .ZN(new_n567));
  AND4_X1   g0367(.A1(new_n231), .A2(new_n262), .A3(new_n567), .A4(G87), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n306), .A2(new_n231), .A3(G87), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(KEYINPUT22), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n231), .A2(G107), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G116), .ZN(new_n574));
  INV_X1    g0374(.A(new_n358), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n408), .A2(new_n231), .ZN(new_n576));
  OAI221_X1 g0376(.A(new_n573), .B1(new_n574), .B2(new_n575), .C1(new_n576), .C2(new_n572), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n570), .A2(KEYINPUT24), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT24), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n262), .A2(new_n567), .A3(new_n231), .A4(G87), .ZN(new_n580));
  AOI211_X1 g0380(.A(G20), .B(new_n211), .C1(new_n268), .C2(new_n270), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT22), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n576), .A2(new_n572), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n573), .B1(new_n575), .B2(new_n574), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n579), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n281), .B1(new_n578), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G200), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n525), .A2(new_n527), .ZN(new_n590));
  INV_X1    g0390(.A(G257), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G1698), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(G250), .B2(G1698), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n270), .B2(new_n268), .ZN(new_n594));
  INV_X1    g0394(.A(G294), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n260), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n325), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n526), .A2(new_n520), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(G264), .A3(new_n301), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n589), .B1(new_n590), .B2(new_n600), .ZN(new_n601));
  OAI22_X1  g0401(.A1(new_n263), .A2(new_n593), .B1(new_n260), .B2(new_n595), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(new_n325), .B1(new_n529), .B2(G264), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n319), .A3(new_n528), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n376), .B(new_n571), .C1(KEYINPUT88), .C2(KEYINPUT25), .ZN(new_n606));
  NAND2_X1  g0406(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n608), .A2(new_n609), .B1(new_n477), .B2(G107), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n588), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(G169), .B1(new_n590), .B2(new_n600), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n603), .A2(G179), .A3(new_n528), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT24), .B1(new_n570), .B2(new_n577), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n583), .A2(new_n579), .A3(new_n586), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n379), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n610), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n525), .A2(new_n527), .B1(new_n529), .B2(G270), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n591), .A2(new_n334), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n218), .A2(G1698), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n268), .B2(new_n270), .ZN(new_n626));
  INV_X1    g0426(.A(G303), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n262), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n622), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n276), .A2(G303), .ZN(new_n630));
  OAI211_X1 g0430(.A(KEYINPUT85), .B(new_n630), .C1(new_n263), .C2(new_n625), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n631), .A3(new_n325), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n621), .A2(new_n632), .A3(G190), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n589), .B1(new_n621), .B2(new_n632), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT86), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n377), .B2(G116), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n288), .A2(KEYINPUT86), .A3(new_n574), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n477), .A2(G116), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n498), .B(new_n231), .C1(G33), .C2(new_n461), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n574), .A2(G20), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n281), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT20), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n633), .A2(new_n634), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n621), .A2(new_n632), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n333), .B1(new_n638), .B2(new_n643), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(KEYINPUT21), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n644), .A2(new_n621), .A3(new_n632), .A4(G179), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT21), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n645), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n620), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n443), .A2(new_n566), .A3(new_n653), .ZN(G372));
  INV_X1    g0454(.A(new_n443), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n479), .A2(new_n492), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT84), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n479), .A2(new_n492), .A3(KEYINPUT84), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n660), .A2(new_n559), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT91), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n559), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n557), .B1(new_n562), .B2(new_n351), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(KEYINPUT91), .A3(new_n541), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n470), .A2(new_n475), .A3(new_n478), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT89), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n449), .B1(new_n263), .B2(new_n446), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n325), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n668), .B(new_n325), .C1(new_n472), .C2(new_n473), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n471), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n394), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n333), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n489), .A2(new_n491), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n667), .A2(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n664), .A2(new_n666), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n662), .B1(new_n678), .B2(new_n661), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT90), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n680), .B(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n559), .B1(new_n563), .B2(new_n565), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n588), .A2(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n646), .A2(new_n647), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT21), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n649), .A3(new_n648), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n611), .B(new_n677), .C1(new_n684), .C2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n682), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n679), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n655), .A2(new_n691), .ZN(new_n692));
  AOI221_X4 g0492(.A(KEYINPUT18), .B1(new_n312), .B2(new_n313), .C1(new_n282), .C2(new_n291), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n317), .B1(new_n292), .B2(new_n314), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n437), .B1(new_n434), .B2(new_n435), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT72), .B1(new_n412), .B2(new_n428), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n429), .A2(new_n436), .A3(KEYINPUT92), .A4(new_n437), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n373), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n371), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n330), .A2(new_n331), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n696), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n398), .A2(new_n399), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n402), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n692), .A2(new_n708), .ZN(G369));
  NAND2_X1  g0509(.A1(new_n376), .A2(new_n231), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G213), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G343), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n644), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n652), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n688), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n716), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n684), .A2(new_n715), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT93), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n620), .ZN(new_n725));
  INV_X1    g0525(.A(new_n715), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n588), .B2(new_n610), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT94), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n684), .A2(new_n726), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n718), .A2(new_n715), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n732), .B1(new_n728), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(G399));
  INV_X1    g0535(.A(new_n223), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G41), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n463), .A2(G116), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(G1), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n228), .B2(new_n738), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT28), .ZN(new_n742));
  INV_X1    g0542(.A(new_n689), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n560), .A2(KEYINPUT82), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n562), .A2(G190), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n540), .A2(new_n319), .A3(new_n531), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n558), .B1(new_n747), .B2(KEYINPUT82), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n746), .A2(new_n748), .B1(new_n541), .B2(new_n665), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n743), .A2(new_n749), .A3(KEYINPUT97), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT97), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n683), .B2(new_n689), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT96), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n674), .A2(new_n667), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n680), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n559), .B2(new_n663), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n661), .B1(new_n757), .B2(new_n666), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n665), .A2(new_n658), .A3(new_n659), .A4(new_n541), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n682), .B1(new_n759), .B2(KEYINPUT26), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n754), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n678), .A2(KEYINPUT26), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n680), .B(KEYINPUT90), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n660), .A2(new_n559), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(new_n661), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n762), .A2(new_n765), .A3(KEYINPUT96), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n753), .B1(new_n761), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT29), .B1(new_n767), .B2(new_n715), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT29), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n691), .A2(new_n769), .A3(new_n726), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(G179), .B1(new_n603), .B2(new_n528), .ZN(new_n772));
  AND3_X1   g0572(.A1(new_n772), .A2(new_n673), .A3(new_n646), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n514), .A2(new_n532), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n600), .A2(new_n457), .A3(new_n450), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n621), .A2(new_n632), .A3(G179), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(KEYINPUT95), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT95), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n621), .A2(new_n632), .A3(new_n779), .A4(G179), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n562), .A2(new_n776), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n775), .A2(new_n781), .A3(KEYINPUT30), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n778), .A2(new_n780), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT30), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n783), .A2(new_n784), .A3(new_n562), .A4(new_n776), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n782), .A2(new_n785), .A3(KEYINPUT31), .A4(new_n715), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n620), .A2(new_n652), .A3(new_n726), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n566), .B2(new_n787), .ZN(new_n788));
  AND4_X1   g0588(.A1(new_n562), .A2(new_n776), .A3(new_n778), .A4(new_n780), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n772), .A2(new_n673), .A3(new_n646), .ZN(new_n790));
  OAI21_X1  g0590(.A(KEYINPUT30), .B1(new_n562), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n726), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(KEYINPUT31), .B1(new_n792), .B2(new_n782), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G330), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n771), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n742), .B1(new_n799), .B2(G1), .ZN(G364));
  NOR2_X1   g0600(.A1(new_n719), .A2(G330), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n287), .A2(G20), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n284), .B1(new_n802), .B2(G45), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n737), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n721), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G13), .A2(G33), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n719), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n262), .A2(new_n223), .ZN(new_n812));
  INV_X1    g0612(.A(G355), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n812), .A2(new_n813), .B1(G116), .B2(new_n223), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n247), .A2(new_n298), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n263), .A2(new_n223), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n298), .B2(new_n229), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n230), .B1(G20), .B2(new_n333), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n809), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n805), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n231), .A2(G179), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n394), .A2(G190), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n211), .ZN(new_n825));
  NAND2_X1  g0625(.A1(G20), .A2(G179), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT98), .Z(new_n827));
  NOR2_X1   g0627(.A1(new_n319), .A2(G200), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(G190), .A2(G200), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n252), .A2(new_n829), .B1(new_n831), .B2(new_n215), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n394), .A2(new_n319), .A3(new_n823), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n825), .B(new_n832), .C1(G107), .C2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n231), .B1(new_n828), .B2(new_n351), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(KEYINPUT100), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(KEYINPUT100), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(G97), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n823), .A2(new_n830), .ZN(new_n843));
  INV_X1    g0643(.A(G159), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(new_n276), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n827), .A2(G200), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n319), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(G190), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G50), .A2(new_n850), .B1(new_n851), .B2(G68), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n835), .A2(new_n842), .A3(new_n848), .A4(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(G283), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n833), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n843), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n262), .B(new_n855), .C1(G329), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(G322), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n627), .A2(new_n824), .B1(new_n829), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n831), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(G311), .B2(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(KEYINPUT101), .B(G326), .Z(new_n862));
  NAND2_X1  g0662(.A1(new_n850), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(KEYINPUT33), .B(G317), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n841), .A2(G294), .B1(new_n851), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n857), .A2(new_n861), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n853), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n822), .B1(new_n867), .B2(new_n819), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n806), .B1(new_n811), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(G396));
  NAND2_X1  g0670(.A1(new_n691), .A2(new_n726), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n439), .A2(new_n726), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n441), .B(new_n873), .C1(new_n698), .C2(new_n699), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT103), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n700), .A2(new_n701), .A3(new_n872), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT103), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n438), .A2(new_n877), .A3(new_n441), .A4(new_n873), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n726), .B(new_n881), .C1(new_n679), .C2(new_n690), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n805), .B1(new_n883), .B2(new_n797), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n797), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n819), .A2(new_n807), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT102), .Z(new_n887));
  OAI21_X1  g0687(.A(new_n805), .B1(new_n887), .B2(G77), .ZN(new_n888));
  INV_X1    g0688(.A(G311), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n276), .B1(new_n889), .B2(new_n843), .C1(new_n829), .C2(new_n595), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(G97), .B2(new_n841), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n834), .A2(G87), .ZN(new_n892));
  INV_X1    g0692(.A(new_n824), .ZN(new_n893));
  AOI22_X1  g0693(.A1(G107), .A2(new_n893), .B1(new_n860), .B2(G116), .ZN(new_n894));
  AOI22_X1  g0694(.A1(G283), .A2(new_n851), .B1(new_n850), .B2(G303), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n891), .A2(new_n892), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n829), .ZN(new_n897));
  AOI22_X1  g0697(.A1(G143), .A2(new_n897), .B1(new_n860), .B2(G159), .ZN(new_n898));
  INV_X1    g0698(.A(new_n850), .ZN(new_n899));
  INV_X1    g0699(.A(G137), .ZN(new_n900));
  INV_X1    g0700(.A(G150), .ZN(new_n901));
  INV_X1    g0701(.A(new_n851), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n898), .B1(new_n899), .B2(new_n900), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT34), .Z(new_n904));
  INV_X1    g0704(.A(G132), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n306), .B1(new_n905), .B2(new_n843), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n833), .A2(new_n209), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n906), .B(new_n907), .C1(G50), .C2(new_n893), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n252), .B2(new_n840), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n896), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n888), .B1(new_n910), .B2(new_n819), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n808), .B2(new_n881), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n885), .A2(new_n912), .ZN(G384));
  OR2_X1    g0713(.A1(new_n553), .A2(KEYINPUT35), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n553), .A2(KEYINPUT35), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n914), .A2(G116), .A3(new_n232), .A4(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT36), .Z(new_n917));
  OR3_X1    g0717(.A1(new_n228), .A2(new_n215), .A3(new_n253), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n202), .A2(G68), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n284), .B(G13), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n443), .B1(new_n768), .B2(new_n770), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(new_n707), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n713), .B1(new_n282), .B2(new_n291), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n312), .A2(new_n313), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n926), .A2(new_n713), .B1(new_n282), .B2(new_n291), .ZN(new_n927));
  INV_X1    g0727(.A(new_n328), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT37), .ZN(new_n930));
  INV_X1    g0730(.A(new_n713), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n292), .B1(new_n314), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n930), .B1(new_n932), .B2(KEYINPUT105), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n332), .A2(new_n925), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT105), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT37), .B1(new_n927), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n328), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n273), .A2(new_n281), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT7), .B1(new_n306), .B2(G20), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G68), .A3(new_n271), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT16), .B1(new_n942), .B2(new_n258), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n291), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n931), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n695), .B2(new_n704), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT38), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n930), .B1(new_n927), .B2(new_n928), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n944), .B1(new_n314), .B2(new_n931), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(KEYINPUT37), .A3(new_n328), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n946), .A2(new_n947), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n924), .B1(new_n939), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n371), .A2(new_n715), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n947), .B1(new_n946), .B2(new_n951), .ZN(new_n955));
  INV_X1    g0755(.A(new_n945), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n332), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n928), .A2(new_n930), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n937), .A2(new_n930), .B1(new_n958), .B2(new_n949), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT38), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n955), .A2(KEYINPUT39), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n953), .A2(new_n954), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n696), .A2(new_n713), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n370), .A2(new_n726), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n373), .B(new_n966), .C1(new_n357), .C2(new_n370), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n345), .A2(new_n347), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n353), .A2(KEYINPUT14), .B1(new_n968), .B2(G179), .ZN(new_n969));
  INV_X1    g0769(.A(new_n356), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n355), .B1(new_n348), .B2(new_n349), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n373), .B(new_n969), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT104), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n965), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n967), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n973), .B1(new_n972), .B2(new_n965), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT38), .B1(new_n957), .B2(new_n959), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n952), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n438), .A2(new_n715), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n977), .B(new_n979), .C1(new_n882), .C2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n964), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n923), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n955), .A2(new_n960), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n967), .A2(new_n974), .ZN(new_n986));
  INV_X1    g0786(.A(new_n976), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n879), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT107), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n784), .B1(new_n773), .B2(new_n774), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n715), .B1(new_n990), .B2(new_n781), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n789), .A2(new_n791), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT31), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n792), .A2(KEYINPUT107), .A3(new_n782), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n985), .B(new_n988), .C1(new_n996), .C2(new_n788), .ZN(new_n997));
  XNOR2_X1  g0797(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n881), .B1(new_n975), .B2(new_n976), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n788), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT40), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n332), .A2(new_n925), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n933), .A2(new_n929), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n938), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n947), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1005), .B1(new_n1009), .B2(new_n960), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1000), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n655), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n795), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n984), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n284), .B2(new_n802), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n984), .A2(new_n1017), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n921), .B1(new_n1019), .B2(new_n1020), .ZN(G367));
  NOR2_X1   g0821(.A1(new_n239), .A2(new_n816), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n820), .B1(new_n469), .B2(new_n223), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n805), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n841), .A2(G68), .B1(G159), .B2(new_n851), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n202), .A2(new_n831), .B1(new_n829), .B2(new_n901), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n833), .A2(new_n215), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n850), .A2(G143), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n262), .B1(new_n843), .B2(new_n900), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n893), .B2(G58), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1025), .A2(new_n1028), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n840), .A2(new_n409), .B1(new_n854), .B2(new_n831), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT113), .Z(new_n1034));
  NOR2_X1   g0834(.A1(new_n824), .A2(new_n574), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1035), .A2(KEYINPUT46), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G294), .B2(new_n851), .ZN(new_n1037));
  INV_X1    g0837(.A(G317), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n263), .B1(new_n1038), .B2(new_n843), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n833), .A2(new_n461), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G303), .C2(new_n897), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(KEYINPUT46), .A2(new_n1035), .B1(new_n850), .B2(G311), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1037), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1032), .B1(new_n1034), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT47), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1024), .B1(new_n1045), .B2(new_n819), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n726), .B1(new_n470), .B2(new_n478), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT108), .Z(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(new_n756), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n763), .A2(new_n1048), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1046), .B1(new_n1051), .B2(new_n810), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n557), .A2(new_n726), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n683), .A2(new_n1053), .B1(new_n559), .B2(new_n726), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1054), .A2(KEYINPUT110), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(KEYINPUT110), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n728), .A2(new_n733), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n732), .ZN(new_n1059));
  XOR2_X1   g0859(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n1060));
  XOR2_X1   g0860(.A(new_n1059), .B(new_n1060), .Z(new_n1061));
  OR2_X1    g0861(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n734), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT45), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n730), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1064), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n730), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1059), .B(new_n1060), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n728), .B(new_n733), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(new_n721), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n799), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n799), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n737), .B(KEYINPUT41), .Z(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n804), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1051), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT43), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT109), .Z(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1062), .A2(new_n1058), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(KEYINPUT42), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n559), .B1(new_n1057), .B2(new_n619), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n726), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT42), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1062), .A2(new_n1089), .A3(new_n1058), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1090), .A2(KEYINPUT111), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(KEYINPUT111), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1086), .B(new_n1088), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1084), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1093), .A2(new_n1084), .A3(new_n1095), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1097), .A2(new_n1067), .A3(new_n1062), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1098), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1100), .A2(new_n1096), .B1(new_n730), .B2(new_n1057), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1052), .B1(new_n1079), .B2(new_n1102), .ZN(G387));
  OR2_X1    g0903(.A1(new_n728), .A2(new_n810), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n243), .A2(new_n298), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1105), .A2(new_n816), .B1(new_n739), .B2(new_n812), .ZN(new_n1106));
  OR3_X1    g0906(.A1(new_n290), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1107));
  AOI21_X1  g0907(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT50), .B1(new_n290), .B2(G50), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1107), .A2(new_n739), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1106), .A2(new_n1110), .B1(new_n217), .B2(new_n736), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n805), .B1(new_n1111), .B2(new_n821), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n263), .B(new_n1040), .C1(G150), .C2(new_n856), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n202), .A2(new_n829), .B1(new_n831), .B2(new_n209), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G77), .B2(new_n893), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n841), .A2(new_n486), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G159), .A2(new_n850), .B1(new_n851), .B2(new_n283), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n306), .B1(new_n862), .B2(new_n856), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n840), .A2(new_n854), .B1(new_n595), .B2(new_n824), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G303), .A2(new_n860), .B1(new_n897), .B2(G317), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n899), .B2(new_n858), .C1(new_n889), .C2(new_n902), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT48), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1123), .B2(new_n1122), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT49), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1119), .B1(new_n574), .B2(new_n833), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1118), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1112), .B1(new_n1129), .B2(new_n819), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1072), .A2(new_n804), .B1(new_n1104), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1073), .A2(new_n737), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n799), .A2(new_n1072), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(G393));
  NAND3_X1  g0934(.A1(new_n1065), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1075), .A2(new_n737), .A3(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n820), .B1(new_n461), .B2(new_n223), .C1(new_n250), .C2(new_n816), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n899), .A2(new_n1038), .B1(new_n829), .B2(new_n889), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT52), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n902), .A2(new_n627), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n840), .A2(new_n574), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n276), .B1(new_n858), .B2(new_n843), .C1(new_n833), .C2(new_n217), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n854), .A2(new_n824), .B1(new_n831), .B2(new_n595), .ZN(new_n1143));
  NOR4_X1   g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n899), .A2(new_n901), .B1(new_n829), .B2(new_n844), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT51), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n841), .A2(G77), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n202), .B2(new_n902), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n263), .B1(G143), .B2(new_n856), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n892), .A2(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n209), .A2(new_n824), .B1(new_n831), .B2(new_n290), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1148), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1139), .A2(new_n1144), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n819), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n805), .B(new_n1137), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n1057), .B2(new_n809), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n1070), .B2(new_n804), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1136), .A2(new_n1157), .ZN(G390));
  NAND2_X1  g0958(.A1(new_n882), .A2(new_n981), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n977), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n954), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n953), .A2(new_n961), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g0965(.A(G330), .B(new_n881), .C1(new_n788), .C2(new_n793), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1166), .A2(new_n977), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n761), .A2(new_n766), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n753), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n726), .A3(new_n881), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n977), .B1(new_n1171), .B2(new_n981), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1009), .A2(new_n960), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1162), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1165), .B(new_n1167), .C1(new_n1172), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1164), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n767), .A2(new_n715), .A3(new_n879), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1160), .B1(new_n1178), .B2(new_n980), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1174), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n795), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n988), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1175), .B(new_n804), .C1(new_n1181), .C2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n805), .B1(new_n887), .B2(new_n283), .ZN(new_n1185));
  INV_X1    g0985(.A(G125), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n262), .B1(new_n843), .B2(new_n1186), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n202), .A2(new_n833), .B1(new_n829), .B2(new_n905), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT54), .B(G143), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1187), .B(new_n1188), .C1(new_n860), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n850), .A2(G128), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n841), .A2(G159), .B1(G137), .B2(new_n851), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n824), .A2(new_n901), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT53), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n907), .B1(G97), .B2(new_n860), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n574), .B2(new_n829), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n262), .B(new_n825), .C1(G294), .C2(new_n856), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G283), .A2(new_n850), .B1(new_n851), .B2(new_n408), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1147), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1196), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1185), .B1(new_n1202), .B2(new_n819), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1176), .B2(new_n808), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1184), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1175), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n655), .A2(new_n1182), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n922), .A2(new_n707), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n715), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n980), .B1(new_n1210), .B2(new_n881), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT115), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n795), .B(new_n879), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1212), .B1(new_n1213), .B2(new_n1160), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1182), .A2(new_n881), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(KEYINPUT115), .A3(new_n977), .ZN(new_n1216));
  AND4_X1   g1016(.A1(new_n1211), .A2(new_n1214), .A3(new_n1167), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1183), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1166), .A2(new_n977), .ZN(new_n1219));
  OAI211_X1 g1019(.A(KEYINPUT114), .B(new_n1159), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT114), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1182), .A2(new_n988), .B1(new_n1166), .B2(new_n977), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1159), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1209), .B1(new_n1217), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n738), .B1(new_n1206), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1165), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1218), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1211), .A2(new_n1214), .A3(new_n1167), .A4(new_n1216), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n1224), .A3(new_n1220), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1229), .A2(new_n1175), .A3(new_n1209), .A4(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1205), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(G378));
  OAI21_X1  g1034(.A(new_n1209), .B1(new_n1206), .B2(new_n1226), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n963), .B(new_n962), .C1(new_n1161), .C2(new_n979), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n795), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1237));
  XOR2_X1   g1037(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1238));
  OR2_X1    g1038(.A1(new_n403), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n403), .A2(new_n1238), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n383), .A2(new_n713), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT118), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1239), .A2(new_n1243), .A3(new_n1240), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1000), .A2(new_n1237), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1247), .B1(new_n1000), .B2(new_n1237), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1236), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1011), .A2(G330), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n998), .B1(new_n1004), .B2(new_n985), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1000), .A2(new_n1237), .A3(new_n1247), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n983), .A3(new_n1255), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1250), .A2(new_n1256), .A3(KEYINPUT57), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1235), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1250), .A2(new_n1256), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1232), .B2(new_n1209), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1258), .B(new_n737), .C1(new_n1260), .C2(KEYINPUT57), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n306), .A2(G41), .ZN(new_n1262));
  AOI211_X1 g1062(.A(G50), .B(new_n1262), .C1(new_n260), .C2(new_n297), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n824), .A2(new_n215), .B1(new_n854), .B2(new_n843), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n461), .A2(new_n902), .B1(new_n899), .B2(new_n574), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(G68), .C2(new_n841), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n833), .A2(new_n252), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n486), .A2(new_n860), .B1(new_n897), .B2(G107), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1266), .A2(new_n1262), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT58), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1263), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n897), .A2(G128), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n1273), .B1(new_n900), .B2(new_n831), .C1(new_n824), .C2(new_n1189), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G132), .B2(new_n851), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n841), .A2(G150), .B1(G125), .B2(new_n850), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT116), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1277), .A2(KEYINPUT116), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1275), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT59), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT117), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1283), .A2(G124), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(G124), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI211_X1 g1086(.A(G33), .B(G41), .C1(new_n1286), .C2(new_n856), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1282), .B(new_n1287), .C1(new_n844), .C2(new_n833), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1281), .A2(KEYINPUT59), .ZN(new_n1289));
  OAI221_X1 g1089(.A(new_n1272), .B1(new_n1271), .B2(new_n1270), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n819), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n804), .B(new_n737), .C1(new_n202), .C2(new_n886), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1291), .B(new_n1292), .C1(new_n1251), .C2(new_n808), .ZN(new_n1293));
  XOR2_X1   g1093(.A(new_n1293), .B(KEYINPUT119), .Z(new_n1294));
  INV_X1    g1094(.A(new_n1259), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n804), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1261), .A2(new_n1296), .ZN(G375));
  NAND2_X1  g1097(.A1(new_n1231), .A2(new_n804), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n805), .B1(new_n887), .B2(G68), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n262), .B(new_n1027), .C1(G303), .C2(new_n856), .ZN(new_n1300));
  OAI22_X1  g1100(.A1(new_n461), .A2(new_n824), .B1(new_n829), .B2(new_n854), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n408), .B2(new_n860), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(G116), .A2(new_n851), .B1(new_n850), .B2(G294), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1300), .A2(new_n1302), .A3(new_n1303), .A4(new_n1116), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n263), .B(new_n1267), .C1(G128), .C2(new_n856), .ZN(new_n1305));
  OAI22_X1  g1105(.A1(new_n844), .A2(new_n824), .B1(new_n829), .B2(new_n900), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(G150), .B2(new_n860), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n851), .A2(new_n1190), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n841), .A2(G50), .B1(G132), .B2(new_n850), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1305), .A2(new_n1307), .A3(new_n1308), .A4(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1304), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1299), .B1(new_n1311), .B2(new_n819), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1160), .B2(new_n808), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1298), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT120), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1231), .B2(new_n1209), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n708), .B(new_n1207), .C1(new_n771), .C2(new_n443), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1318), .A2(new_n1319), .A3(KEYINPUT120), .A4(new_n1230), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1226), .A2(new_n1078), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1315), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1323), .B(KEYINPUT121), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(G381));
  INV_X1    g1125(.A(G375), .ZN(new_n1326));
  NOR4_X1   g1126(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1052), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1102), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n798), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n803), .B1(new_n1330), .B2(new_n1077), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1328), .B1(new_n1329), .B2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1327), .A2(new_n1332), .A3(new_n1324), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1233), .B(new_n1326), .C1(new_n1333), .C2(KEYINPUT122), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1333), .A2(KEYINPUT122), .ZN(new_n1335));
  OR2_X1    g1135(.A1(new_n1334), .A2(new_n1335), .ZN(G407));
  NAND2_X1  g1136(.A1(new_n1326), .A2(new_n1233), .ZN(new_n1337));
  OAI211_X1 g1137(.A(G407), .B(G213), .C1(G343), .C2(new_n1337), .ZN(G409));
  NOR2_X1   g1138(.A1(new_n1231), .A2(new_n1209), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n738), .B1(new_n1339), .B2(KEYINPUT60), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT60), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1341), .B1(new_n1231), .B2(new_n1209), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1340), .B1(new_n1321), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1315), .ZN(new_n1344));
  INV_X1    g1144(.A(G384), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1343), .A2(G384), .A3(new_n1315), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1346), .A2(KEYINPUT125), .A3(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT125), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1226), .A2(KEYINPUT60), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1350), .A2(new_n1317), .A3(new_n1320), .ZN(new_n1351));
  AOI211_X1 g1151(.A(new_n1345), .B(new_n1314), .C1(new_n1351), .C2(new_n1340), .ZN(new_n1352));
  AOI21_X1  g1152(.A(G384), .B1(new_n1343), .B2(new_n1315), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1349), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1348), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(G213), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1356), .A2(G343), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(G2897), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1355), .A2(new_n1358), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1250), .A2(new_n1256), .A3(KEYINPUT123), .ZN(new_n1360));
  AOI21_X1  g1160(.A(KEYINPUT123), .B1(new_n1250), .B2(new_n1256), .ZN(new_n1361));
  NOR3_X1   g1161(.A1(new_n1360), .A2(new_n1361), .A3(new_n803), .ZN(new_n1362));
  OAI21_X1  g1162(.A(KEYINPUT124), .B1(new_n1362), .B2(new_n1294), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1235), .A2(new_n1078), .A3(new_n1295), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT123), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1259), .A2(new_n1365), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1250), .A2(new_n1256), .A3(KEYINPUT123), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1366), .A2(new_n804), .A3(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT124), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1294), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1368), .A2(new_n1369), .A3(new_n1370), .ZN(new_n1371));
  NAND4_X1  g1171(.A1(new_n1363), .A2(new_n1233), .A3(new_n1364), .A4(new_n1371), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1357), .ZN(new_n1373));
  AND2_X1   g1173(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(G375), .A2(G378), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1358), .ZN(new_n1377));
  AOI22_X1  g1177(.A1(new_n1374), .A2(new_n1375), .B1(new_n1376), .B2(new_n1377), .ZN(new_n1378));
  AOI21_X1  g1178(.A(KEYINPUT61), .B1(new_n1359), .B2(new_n1378), .ZN(new_n1379));
  OAI21_X1  g1179(.A(G390), .B1(new_n1332), .B2(KEYINPUT127), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT127), .ZN(new_n1381));
  AND2_X1   g1181(.A1(new_n1136), .A2(new_n1157), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(G387), .A2(new_n1381), .A3(new_n1382), .ZN(new_n1383));
  XNOR2_X1  g1183(.A(G393), .B(G396), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1380), .A2(new_n1383), .A3(new_n1384), .ZN(new_n1385));
  INV_X1    g1185(.A(KEYINPUT126), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(G390), .A2(new_n1386), .ZN(new_n1387));
  INV_X1    g1187(.A(new_n1387), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1384), .B1(new_n1388), .B2(G387), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1382), .A2(KEYINPUT126), .ZN(new_n1390));
  NAND3_X1  g1190(.A1(new_n1332), .A2(new_n1390), .A3(new_n1387), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1389), .A2(new_n1391), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1385), .A2(new_n1392), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1394));
  AOI21_X1  g1194(.A(new_n1233), .B1(new_n1261), .B2(new_n1296), .ZN(new_n1395));
  NOR2_X1   g1195(.A1(new_n1394), .A2(new_n1395), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1355), .A2(new_n1396), .ZN(new_n1397));
  INV_X1    g1197(.A(KEYINPUT63), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1397), .A2(new_n1398), .ZN(new_n1399));
  NAND3_X1  g1199(.A1(new_n1355), .A2(new_n1396), .A3(KEYINPUT63), .ZN(new_n1400));
  NAND4_X1  g1200(.A1(new_n1379), .A2(new_n1393), .A3(new_n1399), .A4(new_n1400), .ZN(new_n1401));
  INV_X1    g1201(.A(KEYINPUT61), .ZN(new_n1402));
  AOI21_X1  g1202(.A(new_n1377), .B1(new_n1348), .B2(new_n1354), .ZN(new_n1403));
  OAI21_X1  g1203(.A(new_n1377), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1404));
  OAI21_X1  g1204(.A(new_n1404), .B1(new_n1394), .B2(new_n1395), .ZN(new_n1405));
  OAI21_X1  g1205(.A(new_n1402), .B1(new_n1403), .B2(new_n1405), .ZN(new_n1406));
  INV_X1    g1206(.A(KEYINPUT62), .ZN(new_n1407));
  AND3_X1   g1207(.A1(new_n1355), .A2(new_n1396), .A3(new_n1407), .ZN(new_n1408));
  AOI21_X1  g1208(.A(new_n1407), .B1(new_n1355), .B2(new_n1396), .ZN(new_n1409));
  NOR3_X1   g1209(.A1(new_n1406), .A2(new_n1408), .A3(new_n1409), .ZN(new_n1410));
  OAI21_X1  g1210(.A(new_n1401), .B1(new_n1410), .B2(new_n1393), .ZN(G405));
  NAND2_X1  g1211(.A1(new_n1337), .A2(new_n1375), .ZN(new_n1412));
  NAND2_X1  g1212(.A1(new_n1412), .A2(new_n1376), .ZN(new_n1413));
  INV_X1    g1213(.A(new_n1355), .ZN(new_n1414));
  OAI21_X1  g1214(.A(new_n1413), .B1(new_n1414), .B2(new_n1412), .ZN(new_n1415));
  NAND3_X1  g1215(.A1(new_n1415), .A2(new_n1392), .A3(new_n1385), .ZN(new_n1416));
  OAI211_X1 g1216(.A(new_n1393), .B(new_n1413), .C1(new_n1414), .C2(new_n1412), .ZN(new_n1417));
  NAND2_X1  g1217(.A1(new_n1416), .A2(new_n1417), .ZN(G402));
endmodule


