//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT64), .Z(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G68), .A2(G238), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n205), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n208), .B(new_n219), .C1(new_n222), .C2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(new_n216), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G264), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G50), .B(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G58), .ZN(new_n236));
  INV_X1    g0036(.A(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  INV_X1    g0039(.A(G107), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n238), .B(new_n243), .Z(G351));
  AND2_X1   g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(new_n220), .ZN(new_n246));
  AND2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT66), .B(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G257), .ZN(new_n251));
  NOR3_X1   g0051(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  OAI211_X1 g0052(.A(G264), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n253));
  OR2_X1    g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G303), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n246), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n259), .B(G45), .C1(new_n260), .C2(KEYINPUT5), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT5), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G41), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT65), .B1(new_n245), .B2(new_n220), .ZN(new_n266));
  AND2_X1   g0066(.A1(G1), .A2(G13), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT65), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n262), .A2(new_n265), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G270), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n270), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n264), .B1(new_n261), .B2(KEYINPUT76), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n263), .A2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT76), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(new_n259), .A4(G45), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n273), .A2(new_n274), .A3(G274), .A4(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n258), .A2(new_n272), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n280), .A2(new_n220), .B1(G20), .B2(new_n242), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G283), .ZN(new_n282));
  INV_X1    g0082(.A(G97), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n282), .B(new_n221), .C1(G33), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT20), .ZN(new_n286));
  OR2_X1    g0086(.A1(new_n286), .A2(KEYINPUT79), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(KEYINPUT79), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n242), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n281), .A2(KEYINPUT79), .A3(new_n284), .A4(new_n286), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n221), .A2(G1), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n294), .A2(G13), .B1(new_n259), .B2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n280), .A2(new_n220), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(G116), .A3(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n289), .A2(new_n292), .A3(new_n293), .A4(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n279), .A2(G169), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT21), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n299), .A2(G169), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT21), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(new_n279), .ZN(new_n304));
  INV_X1    g0104(.A(new_n299), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n279), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n301), .A2(new_n304), .B1(G179), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n279), .A2(G200), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n308), .B(new_n305), .C1(new_n309), .C2(new_n279), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G45), .ZN(new_n312));
  AOI21_X1  g0112(.A(G1), .B1(new_n260), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n273), .A2(G274), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n266), .B2(new_n270), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G238), .ZN(new_n316));
  INV_X1    g0116(.A(G1698), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n250), .A2(new_n216), .B1(new_n227), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT3), .B(G33), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n318), .A2(new_n319), .B1(G33), .B2(G97), .ZN(new_n320));
  INV_X1    g0120(.A(new_n246), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n314), .B(new_n316), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT13), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(KEYINPUT66), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT66), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G1698), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n328));
  INV_X1    g0128(.A(G33), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n328), .A2(new_n249), .B1(new_n329), .B2(new_n283), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n246), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n331), .A2(new_n332), .A3(new_n314), .A4(new_n316), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n323), .A2(new_n333), .A3(KEYINPUT70), .ZN(new_n334));
  OR3_X1    g0134(.A1(new_n322), .A2(KEYINPUT70), .A3(KEYINPUT13), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(G169), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT14), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n323), .A2(new_n333), .A3(G179), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n334), .A2(new_n335), .A3(new_n339), .A4(G169), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n280), .A2(KEYINPUT67), .A3(new_n220), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT67), .B1(new_n280), .B2(new_n220), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n221), .A2(G68), .ZN(new_n345));
  NOR2_X1   g0145(.A1(G20), .A2(G33), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n221), .A2(G33), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n347), .A2(new_n215), .B1(new_n348), .B2(new_n237), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n344), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT11), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n294), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n297), .A2(G68), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n350), .B2(new_n351), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n290), .A2(G68), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT12), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n352), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n341), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n334), .A2(new_n335), .A3(G200), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n323), .A2(new_n333), .A3(G190), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT7), .B1(new_n249), .B2(new_n221), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NOR4_X1   g0166(.A1(new_n247), .A2(new_n248), .A3(new_n366), .A4(G20), .ZN(new_n367));
  OAI21_X1  g0167(.A(G68), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n346), .A2(G159), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G58), .A2(G68), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n371), .B2(new_n201), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n368), .A2(KEYINPUT16), .A3(new_n369), .A4(new_n372), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(new_n296), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT8), .B(G58), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n290), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n344), .A2(new_n294), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n379), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n327), .A2(new_n319), .A3(G223), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G87), .ZN(new_n385));
  OAI211_X1 g0185(.A(G226), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n246), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n315), .A2(G232), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n314), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G169), .ZN(new_n391));
  INV_X1    g0191(.A(G179), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n390), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n383), .A2(KEYINPUT18), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT18), .B1(new_n383), .B2(new_n393), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT73), .ZN(new_n397));
  INV_X1    g0197(.A(G200), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n390), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n388), .A2(new_n309), .A3(new_n389), .A4(new_n314), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(KEYINPUT71), .A3(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n388), .A2(new_n314), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT71), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n309), .A4(new_n389), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n401), .A2(new_n377), .A3(new_n382), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(KEYINPUT72), .A2(KEYINPUT17), .ZN(new_n406));
  OR2_X1    g0206(.A1(KEYINPUT72), .A2(KEYINPUT17), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n405), .B2(new_n407), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n397), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n401), .A2(new_n377), .A3(new_n382), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n411), .A2(KEYINPUT72), .A3(KEYINPUT17), .A4(new_n404), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT73), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n396), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n317), .B1(new_n254), .B2(new_n255), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G223), .ZN(new_n417));
  INV_X1    g0217(.A(G222), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n327), .A2(new_n319), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n417), .B1(new_n237), .B2(new_n319), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n246), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n315), .A2(G226), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n314), .A3(new_n422), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n423), .A2(new_n309), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n381), .A2(G50), .ZN(new_n425));
  INV_X1    g0225(.A(G150), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n378), .A2(new_n348), .B1(new_n426), .B2(new_n347), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n221), .B1(new_n201), .B2(new_n215), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n344), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n425), .B(new_n429), .C1(G50), .C2(new_n290), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT9), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n423), .A2(G200), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n430), .A2(new_n431), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n424), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT10), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n416), .A2(G238), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n436), .B1(new_n240), .B2(new_n319), .C1(new_n227), .C2(new_n419), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n246), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n315), .A2(G244), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n314), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G169), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n379), .A2(new_n346), .B1(G20), .B2(G77), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT15), .B(G87), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(new_n348), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(new_n296), .B1(new_n237), .B2(new_n291), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n297), .A2(G77), .A3(new_n353), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n442), .B(new_n448), .C1(G179), .C2(new_n440), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n423), .A2(new_n441), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n430), .B1(new_n423), .B2(G179), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n440), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT68), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n455), .A3(G190), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT68), .B1(new_n440), .B2(new_n309), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n448), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n440), .A2(G200), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n435), .A2(new_n449), .A3(new_n453), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT69), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n415), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n364), .B(new_n463), .C1(new_n462), .C2(new_n461), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT75), .ZN(new_n465));
  OAI21_X1  g0265(.A(G107), .B1(new_n365), .B2(new_n367), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT6), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n283), .A2(new_n240), .ZN(new_n468));
  NOR2_X1   g0268(.A1(G97), .A2(G107), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n240), .A2(KEYINPUT6), .A3(G97), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G20), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n346), .A2(G77), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n466), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n296), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n295), .B(G97), .C1(new_n342), .C2(new_n343), .ZN(new_n477));
  OR3_X1    g0277(.A1(new_n290), .A2(KEYINPUT74), .A3(G97), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT74), .B1(new_n290), .B2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n465), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  AOI211_X1 g0283(.A(KEYINPUT75), .B(new_n481), .C1(new_n475), .C2(new_n296), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n327), .A2(new_n319), .A3(G244), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n416), .A2(G250), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n327), .A2(new_n319), .A3(KEYINPUT4), .A4(G244), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n487), .A2(new_n282), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n246), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n273), .B(G257), .C1(new_n261), .C2(new_n264), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n492), .A2(new_n278), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n491), .A2(new_n309), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(G200), .B1(new_n491), .B2(new_n493), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n483), .A2(new_n484), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n327), .A2(new_n319), .A3(G250), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n319), .A2(G257), .A3(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n246), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n271), .A2(G264), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n278), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n398), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n501), .A2(new_n309), .A3(new_n502), .A4(new_n278), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n295), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n344), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G107), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT23), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n221), .B2(G107), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n240), .A2(KEYINPUT23), .A3(G20), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n329), .A2(new_n242), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n221), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n221), .B(G87), .C1(new_n247), .C2(new_n248), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n515), .A2(KEYINPUT22), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(KEYINPUT22), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT80), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n515), .B(KEYINPUT22), .ZN(new_n522));
  NAND2_X1  g0322(.A1(KEYINPUT80), .A2(KEYINPUT24), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(new_n520), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n522), .A2(new_n514), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n525), .A3(new_n296), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n290), .A2(G107), .ZN(new_n527));
  XNOR2_X1  g0327(.A(new_n527), .B(KEYINPUT25), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n506), .A2(new_n509), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n491), .A2(G179), .A3(new_n493), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n441), .B1(new_n491), .B2(new_n493), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n366), .B1(new_n319), .B2(G20), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n249), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(G107), .B1(new_n472), .B2(G20), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n297), .B1(new_n535), .B2(new_n474), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n530), .A2(new_n531), .B1(new_n536), .B2(new_n481), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n496), .A2(new_n529), .A3(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n266), .A2(new_n270), .B1(new_n259), .B2(G45), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n259), .A2(G45), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n268), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n539), .A2(G250), .B1(G274), .B2(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n327), .A2(new_n319), .A3(G238), .ZN(new_n543));
  OAI211_X1 g0343(.A(G244), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n544));
  INV_X1    g0344(.A(new_n513), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n246), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G200), .ZN(new_n549));
  NAND3_X1  g0349(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n221), .ZN(new_n551));
  NOR4_X1   g0351(.A1(KEYINPUT77), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT77), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G87), .A2(G97), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n240), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n551), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n319), .A2(new_n221), .A3(G68), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n348), .B2(new_n283), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT78), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT78), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(new_n558), .C1(new_n348), .C2(new_n283), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n556), .A2(new_n557), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(new_n296), .B1(new_n291), .B2(new_n444), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n542), .A2(new_n547), .A3(G190), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n508), .A2(G87), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n549), .A2(new_n564), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n444), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n508), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n513), .B1(new_n416), .B2(G244), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n327), .A2(new_n319), .A3(G238), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n321), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n245), .A2(KEYINPUT65), .A3(new_n220), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n575));
  OAI211_X1 g0375(.A(G250), .B(new_n540), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n541), .A2(G274), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n573), .A2(new_n578), .A3(new_n392), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n441), .B1(new_n542), .B2(new_n547), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n567), .B1(new_n570), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n277), .B(G274), .C1(new_n574), .C2(new_n575), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n584), .A2(new_n274), .B1(new_n500), .B2(new_n246), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n441), .B1(new_n585), .B2(new_n502), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n503), .A2(new_n392), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT81), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n503), .A2(G169), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT81), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n392), .C2(new_n503), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n526), .A2(new_n509), .A3(new_n528), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n582), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n311), .A2(new_n464), .A3(new_n538), .A4(new_n594), .ZN(G372));
  INV_X1    g0395(.A(KEYINPUT83), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n589), .B1(new_n392), .B2(new_n503), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n306), .A2(G179), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n303), .B1(new_n302), .B2(new_n279), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n303), .A2(new_n279), .A3(G169), .A4(new_n299), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n596), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT82), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n579), .B2(new_n580), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n542), .A2(new_n547), .A3(G179), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n573), .A2(new_n578), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(KEYINPUT82), .C1(new_n607), .C2(new_n441), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n570), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n567), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n593), .A2(new_n597), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n307), .A2(new_n612), .A3(KEYINPUT83), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n603), .A2(new_n538), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n582), .ZN(new_n615));
  INV_X1    g0415(.A(new_n537), .ZN(new_n616));
  XNOR2_X1  g0416(.A(KEYINPUT84), .B(KEYINPUT26), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT75), .B1(new_n536), .B2(new_n481), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n476), .A2(new_n465), .A3(new_n482), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n619), .B(new_n620), .C1(new_n531), .C2(new_n530), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n621), .A2(new_n609), .A3(new_n610), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n618), .B1(new_n622), .B2(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(new_n609), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n614), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n464), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n360), .A2(new_n449), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n408), .A2(new_n409), .A3(new_n397), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT73), .B1(new_n412), .B2(new_n413), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n627), .B(new_n363), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n394), .B2(new_n395), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n383), .A2(new_n393), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT18), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n383), .A2(KEYINPUT18), .A3(new_n393), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(KEYINPUT85), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n630), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n452), .B1(new_n638), .B2(new_n435), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n626), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT86), .ZN(G369));
  INV_X1    g0441(.A(new_n593), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n588), .B2(new_n591), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n642), .B2(new_n506), .ZN(new_n644));
  INV_X1    g0444(.A(G13), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(G20), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n259), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n307), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n652), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n644), .B1(new_n642), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n643), .A2(new_n652), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n654), .B1(new_n658), .B2(new_n653), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n652), .A2(new_n299), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n311), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n307), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n644), .A2(new_n653), .B1(new_n598), .B2(new_n655), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(G399));
  OR3_X1    g0467(.A1(new_n552), .A2(new_n555), .A3(G116), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT87), .Z(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n206), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(G1), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n223), .B2(new_n673), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n625), .A2(new_n655), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT88), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n611), .A2(new_n537), .A3(new_n496), .A4(new_n529), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n602), .B1(new_n592), .B2(new_n593), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n624), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n615), .A2(new_n616), .ZN(new_n684));
  INV_X1    g0484(.A(new_n617), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n622), .A2(KEYINPUT26), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n655), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n253), .B(new_n256), .C1(new_n419), .C2(new_n251), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n690), .A2(new_n246), .B1(new_n271), .B2(G270), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n491), .A2(new_n493), .B1(new_n691), .B2(new_n278), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n392), .A3(new_n503), .A4(new_n548), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n491), .A2(new_n607), .A3(new_n493), .A4(G179), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n585), .A2(new_n691), .A3(new_n502), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n258), .A2(new_n272), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n503), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n492), .A2(new_n278), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n246), .B2(new_n490), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n699), .A2(new_n701), .A3(KEYINPUT30), .A4(new_n579), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n693), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n652), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n538), .A2(new_n594), .A3(new_n311), .A4(new_n655), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(KEYINPUT31), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(G330), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n689), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n676), .B1(new_n712), .B2(G1), .ZN(G364));
  NOR2_X1   g0513(.A1(new_n671), .A2(new_n319), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n224), .A2(new_n312), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n714), .B(new_n715), .C1(new_n238), .C2(new_n312), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n319), .A2(G355), .A3(new_n206), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n716), .B(new_n717), .C1(G116), .C2(new_n206), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G13), .A2(G33), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G20), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n220), .B1(G20), .B2(new_n441), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n259), .B1(new_n646), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n672), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT89), .Z(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n221), .A2(G179), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n398), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G107), .ZN(new_n734));
  INV_X1    g0534(.A(G87), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n309), .A2(new_n398), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n730), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n734), .B(new_n319), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT90), .Z(new_n739));
  NOR2_X1   g0539(.A1(G190), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n730), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G159), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT32), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n309), .A2(G179), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n221), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n221), .A2(new_n392), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n736), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n746), .A2(new_n283), .B1(new_n748), .B2(new_n215), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(G190), .A3(new_n398), .ZN(new_n750));
  INV_X1    g0550(.A(G58), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n747), .A2(new_n731), .ZN(new_n752));
  INV_X1    g0552(.A(G68), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n744), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n747), .A2(new_n740), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n739), .B(new_n755), .C1(new_n237), .C2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G294), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n746), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G303), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n737), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  INV_X1    g0562(.A(G329), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n750), .A2(new_n762), .B1(new_n741), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n756), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n761), .B(new_n764), .C1(G311), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n732), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n748), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n319), .B(new_n768), .C1(G326), .C2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n752), .ZN(new_n771));
  INV_X1    g0571(.A(G317), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT33), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n772), .A2(KEYINPUT33), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n766), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n757), .B1(new_n759), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n729), .B1(new_n777), .B2(new_n722), .ZN(new_n778));
  INV_X1    g0578(.A(new_n721), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n724), .B(new_n778), .C1(new_n662), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n663), .A2(new_n729), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n662), .A2(G330), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(G396));
  NOR2_X1   g0583(.A1(new_n449), .A2(new_n652), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n448), .A2(new_n652), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n460), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(new_n786), .B2(new_n449), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n625), .A2(new_n655), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n678), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n787), .B(KEYINPUT93), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n711), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n729), .B1(new_n793), .B2(KEYINPUT94), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(KEYINPUT94), .B2(new_n793), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n792), .A2(new_n711), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G137), .A2(new_n769), .B1(new_n765), .B2(G159), .ZN(new_n798));
  INV_X1    g0598(.A(G143), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n798), .B1(new_n799), .B2(new_n750), .C1(new_n426), .C2(new_n752), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT92), .Z(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n733), .A2(G68), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n803), .B(new_n319), .C1(new_n804), .C2(new_n741), .ZN(new_n805));
  INV_X1    g0605(.A(new_n746), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(G58), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n802), .B(new_n807), .C1(new_n215), .C2(new_n737), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n249), .B1(new_n737), .B2(new_n240), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G303), .A2(new_n769), .B1(new_n771), .B2(G283), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n242), .B2(new_n756), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT91), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n732), .A2(new_n735), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n750), .A2(new_n758), .B1(new_n741), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n814), .B(new_n816), .C1(G97), .C2(new_n806), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n813), .B(new_n817), .C1(new_n812), .C2(new_n811), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n808), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n729), .B1(new_n819), .B2(new_n722), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n722), .A2(new_n719), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(G77), .B2(new_n822), .C1(new_n720), .C2(new_n787), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n797), .A2(new_n823), .ZN(G384));
  INV_X1    g0624(.A(KEYINPUT39), .ZN(new_n825));
  INV_X1    g0625(.A(new_n650), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n383), .A2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n405), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT37), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT97), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n633), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n383), .A2(KEYINPUT97), .A3(new_n393), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n828), .A2(new_n829), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n393), .A2(new_n826), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n375), .A2(new_n344), .A3(new_n376), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n835), .A2(new_n382), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n405), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n836), .A2(new_n650), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n839), .B1(new_n415), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(KEYINPUT38), .B(new_n839), .C1(new_n415), .C2(new_n841), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n825), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n827), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n632), .A2(new_n637), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n412), .A2(new_n413), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n405), .A2(new_n633), .A3(new_n827), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT98), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT98), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n851), .A2(new_n854), .A3(KEYINPUT37), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(new_n833), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n843), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n858), .A2(new_n825), .A3(new_n845), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n846), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n360), .A2(new_n652), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n848), .A2(new_n650), .ZN(new_n864));
  INV_X1    g0664(.A(new_n396), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n628), .B2(new_n629), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n840), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n867), .B2(new_n839), .ZN(new_n868));
  INV_X1    g0668(.A(new_n845), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n784), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n788), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n359), .A2(new_n652), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n360), .A2(new_n363), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n363), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n359), .B(new_n652), .C1(new_n341), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n863), .A2(new_n864), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n689), .A2(new_n464), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n639), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n880), .B(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  INV_X1    g0684(.A(new_n787), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n874), .B2(new_n876), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT100), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n706), .A2(KEYINPUT31), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n704), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n708), .B(KEYINPUT99), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT99), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n708), .B(new_n892), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n707), .A2(new_n893), .A3(KEYINPUT100), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n886), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n884), .B1(new_n870), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n858), .A2(new_n845), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n889), .A2(new_n887), .A3(new_n890), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT100), .B1(new_n707), .B2(new_n893), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n897), .A2(new_n900), .A3(KEYINPUT40), .A4(new_n886), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n464), .A2(new_n900), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n883), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n883), .A2(new_n905), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(KEYINPUT101), .B2(new_n907), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n908), .B1(KEYINPUT101), .B2(new_n907), .C1(new_n259), .C2(new_n646), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n472), .B(KEYINPUT95), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n242), .B1(new_n910), .B2(KEYINPUT35), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(new_n222), .C1(KEYINPUT35), .C2(new_n910), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  OR3_X1    g0713(.A1(new_n753), .A2(KEYINPUT96), .A3(G50), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT96), .B1(new_n753), .B2(G50), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n370), .A2(G77), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n914), .B(new_n915), .C1(new_n223), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n645), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n909), .A2(new_n913), .A3(new_n918), .ZN(G367));
  NAND3_X1  g0719(.A1(new_n619), .A2(new_n620), .A3(new_n652), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n496), .A2(new_n537), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n621), .B2(new_n655), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT102), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n664), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n564), .A2(new_n566), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n652), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n611), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n609), .A2(new_n925), .A3(new_n652), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n923), .A2(new_n643), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n652), .B1(new_n931), .B2(new_n537), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n644), .A2(new_n922), .A3(new_n653), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT42), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n930), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n924), .B(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n672), .B(KEYINPUT41), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n659), .B(new_n663), .Z(new_n940));
  NAND2_X1  g0740(.A1(new_n664), .A2(KEYINPUT103), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n666), .A2(new_n922), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT45), .Z(new_n944));
  NOR2_X1   g0744(.A1(new_n666), .A2(new_n922), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n712), .B(new_n940), .C1(new_n942), .C2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n942), .B2(new_n947), .ZN(new_n949));
  INV_X1    g0749(.A(new_n712), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n939), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n938), .B1(new_n951), .B2(new_n725), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n732), .A2(new_n283), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G283), .B2(new_n765), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n772), .B2(new_n741), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n319), .B(new_n955), .C1(G294), .C2(new_n771), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT46), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n737), .A2(new_n957), .A3(new_n242), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n957), .B1(new_n737), .B2(new_n242), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n240), .B2(new_n746), .ZN(new_n960));
  XNOR2_X1  g0760(.A(KEYINPUT104), .B(G311), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n958), .B(new_n960), .C1(new_n769), .C2(new_n961), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n956), .B(new_n962), .C1(new_n760), .C2(new_n750), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n756), .A2(new_n215), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n319), .B1(new_n732), .B2(new_n237), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT105), .Z(new_n966));
  INV_X1    g0766(.A(G137), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n737), .A2(new_n751), .B1(new_n741), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT106), .ZN(new_n969));
  AOI22_X1  g0769(.A1(G143), .A2(new_n769), .B1(new_n771), .B2(G159), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n746), .A2(new_n753), .ZN(new_n971));
  INV_X1    g0771(.A(new_n750), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n971), .B1(G150), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n966), .A2(new_n969), .A3(new_n970), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n963), .B1(new_n964), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n729), .B1(new_n976), .B2(new_n722), .ZN(new_n977));
  INV_X1    g0777(.A(new_n714), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n723), .B1(new_n206), .B2(new_n444), .C1(new_n233), .C2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n927), .A2(new_n721), .A3(new_n928), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n952), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(G387));
  INV_X1    g0783(.A(new_n940), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n673), .B1(new_n950), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n950), .B2(new_n984), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n742), .A2(G326), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G322), .A2(new_n769), .B1(new_n765), .B2(G303), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n771), .A2(new_n961), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(new_n772), .C2(new_n750), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT48), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n767), .B2(new_n746), .C1(new_n758), .C2(new_n737), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT49), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n319), .B(new_n987), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n993), .B2(new_n992), .C1(new_n242), .C2(new_n732), .ZN(new_n995));
  INV_X1    g0795(.A(new_n737), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G77), .A2(new_n996), .B1(new_n742), .B2(G150), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n215), .B2(new_n750), .C1(new_n753), .C2(new_n756), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n806), .A2(new_n568), .ZN(new_n999));
  INV_X1    g0799(.A(G159), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n999), .B1(new_n1000), .B2(new_n748), .C1(new_n378), .C2(new_n752), .ZN(new_n1001));
  OR4_X1    g0801(.A1(new_n249), .A2(new_n998), .A3(new_n1001), .A4(new_n953), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n995), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n729), .B1(new_n1003), .B2(new_n722), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n669), .A2(new_n206), .A3(new_n319), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(G107), .B2(new_n206), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT107), .Z(new_n1007));
  INV_X1    g0807(.A(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n379), .B2(new_n215), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n378), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1009), .A2(G45), .A3(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n670), .B(new_n1011), .C1(new_n753), .C2(new_n237), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n714), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n230), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1013), .B1(G45), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n723), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1004), .B(new_n1016), .C1(new_n658), .C2(new_n779), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n986), .B(new_n1017), .C1(new_n725), .C2(new_n984), .ZN(G393));
  OAI22_X1  g0818(.A1(new_n737), .A2(new_n767), .B1(new_n741), .B2(new_n762), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT111), .Z(new_n1020));
  OAI22_X1  g0820(.A1(new_n750), .A2(new_n815), .B1(new_n748), .B2(new_n772), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n249), .B1(new_n756), .B2(new_n758), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n734), .B1(new_n760), .B2(new_n752), .C1(new_n242), .C2(new_n746), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1020), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n750), .A2(new_n1000), .B1(new_n748), .B2(new_n426), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT108), .Z(new_n1028));
  AND2_X1   g0828(.A1(new_n1028), .A2(KEYINPUT51), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1028), .A2(KEYINPUT51), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n249), .B(new_n814), .C1(G68), .C2(new_n996), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n215), .A2(new_n752), .B1(new_n756), .B2(new_n378), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT109), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(KEYINPUT109), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n806), .A2(G77), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1029), .A2(new_n1030), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n742), .A2(G143), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1026), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT112), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n722), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n728), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n923), .A2(new_n779), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n243), .A2(new_n714), .B1(G97), .B2(new_n671), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1043), .C1(new_n723), .C2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n947), .B(new_n665), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1045), .B1(new_n1046), .B2(new_n726), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n949), .A2(new_n673), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1046), .B1(new_n712), .B2(new_n940), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(G390));
  OAI211_X1 g0850(.A(G330), .B(new_n886), .C1(new_n891), .C2(new_n894), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT114), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n900), .A2(new_n1053), .A3(G330), .A4(new_n886), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n877), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n710), .B2(new_n885), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n710), .A2(new_n1055), .A3(new_n885), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n791), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1059), .A2(new_n900), .A3(G330), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n874), .A2(KEYINPUT113), .A3(new_n876), .ZN(new_n1061));
  AOI21_X1  g0861(.A(KEYINPUT113), .B1(new_n874), .B2(new_n876), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1058), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n786), .A2(new_n449), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1065), .B(new_n655), .C1(new_n683), .C2(new_n686), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n871), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1057), .A2(new_n872), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n464), .A2(G330), .A3(new_n900), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n881), .A2(new_n639), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(KEYINPUT39), .B1(new_n868), .B2(new_n869), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n862), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n878), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n858), .A2(new_n825), .A3(new_n845), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1073), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1067), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1078), .A2(new_n897), .A3(new_n1074), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1079), .A3(new_n1058), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1078), .A2(new_n897), .A3(new_n1074), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n860), .B2(new_n1075), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1080), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n673), .B1(new_n1072), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1084), .B2(new_n1072), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n726), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n737), .A2(new_n735), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n803), .B1(new_n242), .B2(new_n750), .C1(new_n758), .C2(new_n741), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G77), .C2(new_n806), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n283), .A2(new_n756), .B1(new_n752), .B2(new_n240), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1091), .A2(KEYINPUT115), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(KEYINPUT115), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(new_n767), .C2(new_n748), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT116), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n319), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1090), .B(new_n1096), .C1(new_n1095), .C2(new_n1094), .ZN(new_n1097));
  INV_X1    g0897(.A(G125), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n741), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(G128), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n748), .A2(new_n1100), .B1(new_n752), .B2(new_n967), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT53), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n737), .B2(new_n426), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n996), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n750), .A2(new_n804), .B1(new_n732), .B2(new_n215), .ZN(new_n1106));
  XOR2_X1   g0906(.A(KEYINPUT54), .B(G143), .Z(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n765), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n249), .B1(new_n806), .B2(G159), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1105), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1097), .B1(new_n1099), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n729), .B1(new_n1111), .B2(new_n722), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n379), .B2(new_n822), .C1(new_n861), .C2(new_n720), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1086), .A2(new_n1087), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(G378));
  NAND3_X1  g0915(.A1(new_n896), .A2(G330), .A3(new_n901), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT119), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n896), .A2(KEYINPUT119), .A3(G330), .A4(new_n901), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n435), .A2(new_n453), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n430), .A2(new_n826), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT55), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1124), .A2(KEYINPUT56), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT56), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1118), .A2(new_n1119), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n902), .A2(new_n1128), .A3(KEYINPUT119), .A4(G330), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n880), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1130), .A2(new_n880), .A3(new_n1131), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n726), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n971), .B1(G97), .B2(new_n771), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n242), .B2(new_n748), .ZN(new_n1139));
  AOI211_X1 g0939(.A(G41), .B(new_n319), .C1(new_n996), .C2(G77), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1141), .A2(KEYINPUT117), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(KEYINPUT117), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n732), .A2(new_n751), .B1(new_n741), .B2(new_n767), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n568), .B2(new_n765), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1139), .B(new_n1146), .C1(G107), .C2(new_n972), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT58), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n748), .A2(new_n1098), .B1(new_n752), .B2(new_n804), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n972), .A2(G128), .B1(new_n765), .B2(G137), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1107), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n737), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1149), .B(new_n1152), .C1(G150), .C2(new_n806), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT59), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G41), .B1(new_n742), .B2(G124), .ZN(new_n1155));
  AOI21_X1  g0955(.A(G33), .B1(new_n733), .B2(G159), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n215), .B1(new_n247), .B2(G41), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n722), .B1(new_n1148), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n728), .B1(G50), .B2(new_n822), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT118), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(new_n1129), .C2(new_n720), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1137), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1071), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1083), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1077), .A2(new_n1079), .A3(new_n1058), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1165), .B1(new_n1168), .B2(new_n1069), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT120), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1057), .A2(new_n872), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1071), .B1(new_n1084), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT120), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1171), .A2(new_n1176), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n672), .B1(new_n1177), .B2(KEYINPUT57), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1175), .A2(KEYINPUT120), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1170), .B(new_n1071), .C1(new_n1084), .C2(new_n1174), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT57), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1130), .A2(new_n880), .A3(new_n1131), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT121), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n880), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1183), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1181), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1164), .B1(new_n1178), .B2(new_n1188), .ZN(G375));
  INV_X1    g0989(.A(new_n1072), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n939), .B(KEYINPUT122), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT123), .Z(new_n1194));
  NAND2_X1  g0994(.A1(new_n1063), .A2(new_n719), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n737), .A2(new_n283), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n750), .A2(new_n767), .B1(new_n756), .B2(new_n240), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(G303), .C2(new_n742), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n748), .A2(new_n758), .B1(new_n752), .B2(new_n242), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G77), .B2(new_n733), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1198), .A2(new_n249), .A3(new_n999), .A4(new_n1200), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT124), .Z(new_n1202));
  NOR2_X1   g1002(.A1(new_n737), .A2(new_n1000), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n748), .A2(new_n804), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT125), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n750), .A2(new_n967), .B1(new_n741), .B2(new_n1100), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G150), .B2(new_n765), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n249), .B1(new_n806), .B2(G50), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n771), .A2(new_n1107), .B1(new_n733), .B2(G58), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1202), .B1(new_n1203), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n729), .B1(new_n1211), .B2(new_n722), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1195), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n753), .B2(new_n821), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1174), .B2(new_n726), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1194), .A2(new_n1215), .ZN(G381));
  NOR2_X1   g1016(.A1(G375), .A2(G378), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(G407));
  INV_X1    g1020(.A(new_n1217), .ZN(new_n1221));
  OAI211_X1 g1021(.A(G407), .B(G213), .C1(G343), .C2(new_n1221), .ZN(G409));
  NOR2_X1   g1022(.A1(new_n982), .A2(G390), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  XOR2_X1   g1024(.A(G393), .B(G396), .Z(new_n1225));
  NAND2_X1  g1025(.A1(new_n982), .A2(G390), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1225), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT121), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n726), .B1(new_n1231), .B2(new_n1184), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1136), .B(new_n1191), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1232), .A2(new_n1114), .A3(new_n1233), .A4(new_n1163), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n651), .A2(G213), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(G375), .A2(G378), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1179), .A2(new_n1180), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n673), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1231), .B2(new_n1184), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1114), .B1(new_n1245), .B2(new_n1164), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT126), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT60), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n673), .B1(new_n1192), .B2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n1190), .C1(new_n1249), .C2(new_n1192), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(G384), .A2(new_n1251), .A3(new_n1215), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G384), .B1(new_n1251), .B2(new_n1215), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n651), .A2(G213), .A3(G2897), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1239), .A2(new_n1248), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1236), .A2(new_n1237), .A3(new_n1263), .A4(new_n1255), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1261), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1239), .A2(new_n1248), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1263), .B1(new_n1266), .B2(new_n1255), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1230), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(KEYINPUT63), .A3(new_n1255), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1236), .A2(new_n1237), .A3(new_n1255), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1236), .A2(new_n1237), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1270), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1269), .A2(new_n1273), .A3(new_n1262), .A4(new_n1229), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1268), .A2(new_n1274), .ZN(G405));
  OAI21_X1  g1075(.A(KEYINPUT127), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT127), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1255), .A2(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1221), .A2(new_n1276), .A3(new_n1237), .A4(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1277), .B(new_n1255), .C1(new_n1217), .C2(new_n1246), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(new_n1229), .ZN(G402));
endmodule


