

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n595), .A2(n570), .ZN(n829) );
  XNOR2_X1 U553 ( .A(G2104), .B(KEYINPUT66), .ZN(n559) );
  NAND2_X1 U554 ( .A1(G8), .A2(n681), .ZN(n690) );
  INV_X1 U555 ( .A(G2105), .ZN(n560) );
  XNOR2_X1 U556 ( .A(n531), .B(KEYINPUT15), .ZN(n1015) );
  OR2_X1 U557 ( .A1(n729), .A2(n728), .ZN(n518) );
  BUF_X2 U558 ( .A(n926), .Z(n519) );
  NOR2_X1 U559 ( .A1(n560), .A2(n559), .ZN(n926) );
  NOR2_X2 U560 ( .A1(G2104), .A2(G2105), .ZN(n555) );
  AND2_X1 U561 ( .A1(n552), .A2(n547), .ZN(n546) );
  OR2_X1 U562 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U563 ( .A1(G1966), .A2(n690), .ZN(n707) );
  INV_X1 U564 ( .A(n681), .ZN(n678) );
  BUF_X2 U565 ( .A(n649), .Z(n681) );
  NAND2_X1 U566 ( .A1(n639), .A2(n759), .ZN(n649) );
  BUF_X1 U567 ( .A(n632), .Z(n556) );
  AND2_X1 U568 ( .A1(n560), .A2(G101), .ZN(n533) );
  BUF_X1 U569 ( .A(n789), .Z(G160) );
  XNOR2_X1 U570 ( .A(n638), .B(KEYINPUT65), .ZN(n789) );
  NOR2_X1 U571 ( .A1(n729), .A2(n728), .ZN(n741) );
  NOR2_X1 U572 ( .A1(n649), .A2(n975), .ZN(n640) );
  NAND2_X1 U573 ( .A1(n1015), .A2(n655), .ZN(n548) );
  INV_X1 U574 ( .A(KEYINPUT104), .ZN(n537) );
  AND2_X1 U575 ( .A1(n540), .A2(KEYINPUT104), .ZN(n538) );
  XNOR2_X1 U576 ( .A(n646), .B(KEYINPUT77), .ZN(n532) );
  NOR2_X1 U577 ( .A1(n1010), .A2(n655), .ZN(n544) );
  NOR2_X1 U578 ( .A1(n661), .A2(n660), .ZN(n672) );
  XNOR2_X1 U579 ( .A(KEYINPUT100), .B(KEYINPUT30), .ZN(n683) );
  XNOR2_X1 U580 ( .A(n703), .B(n702), .ZN(n730) );
  XNOR2_X1 U581 ( .A(KEYINPUT102), .B(KEYINPUT32), .ZN(n702) );
  NAND2_X1 U582 ( .A1(KEYINPUT33), .A2(n537), .ZN(n536) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n827) );
  NOR2_X1 U584 ( .A1(n740), .A2(n742), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n521), .A2(n648), .ZN(n531) );
  NOR2_X1 U586 ( .A1(n647), .A2(n532), .ZN(n521) );
  AND2_X1 U587 ( .A1(n528), .A2(n774), .ZN(n522) );
  OR2_X1 U588 ( .A1(n690), .A2(n726), .ZN(n523) );
  AND2_X1 U589 ( .A1(n523), .A2(n536), .ZN(n524) );
  INV_X1 U590 ( .A(KEYINPUT33), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n545), .A2(n544), .ZN(n543) );
  NAND2_X1 U592 ( .A1(n525), .A2(n787), .ZN(n788) );
  NAND2_X1 U593 ( .A1(n529), .A2(n526), .ZN(n525) );
  AND2_X1 U594 ( .A1(n527), .A2(n522), .ZN(n526) );
  NAND2_X1 U595 ( .A1(n741), .A2(n742), .ZN(n527) );
  NAND2_X1 U596 ( .A1(n740), .A2(n742), .ZN(n528) );
  NAND2_X1 U597 ( .A1(n518), .A2(n530), .ZN(n529) );
  NAND2_X1 U598 ( .A1(n559), .A2(n533), .ZN(n628) );
  AND2_X1 U599 ( .A1(n559), .A2(n560), .ZN(n626) );
  XNOR2_X1 U600 ( .A(n724), .B(n542), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n541), .A2(n538), .ZN(n535) );
  NOR2_X1 U602 ( .A1(n539), .A2(n534), .ZN(n727) );
  NAND2_X1 U603 ( .A1(n535), .A2(n524), .ZN(n534) );
  NOR2_X1 U604 ( .A1(n541), .A2(KEYINPUT104), .ZN(n539) );
  INV_X1 U605 ( .A(KEYINPUT64), .ZN(n542) );
  NOR2_X1 U606 ( .A1(n643), .A2(n1010), .ZN(n654) );
  NAND2_X1 U607 ( .A1(n546), .A2(n543), .ZN(n554) );
  INV_X1 U608 ( .A(n643), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n551), .A2(n550), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n1010), .A2(n655), .ZN(n550) );
  INV_X1 U612 ( .A(n1015), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n643), .A2(n553), .ZN(n552) );
  NOR2_X1 U614 ( .A1(n1015), .A2(KEYINPUT98), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n656), .A2(n554), .ZN(n658) );
  AND2_X1 U616 ( .A1(n649), .A2(G1341), .ZN(n641) );
  INV_X1 U617 ( .A(KEYINPUT98), .ZN(n655) );
  INV_X1 U618 ( .A(KEYINPUT99), .ZN(n657) );
  NOR2_X1 U619 ( .A1(n672), .A2(n1012), .ZN(n673) );
  NOR2_X1 U620 ( .A1(n688), .A2(n687), .ZN(n689) );
  INV_X1 U621 ( .A(KEYINPUT23), .ZN(n627) );
  INV_X1 U622 ( .A(KEYINPUT106), .ZN(n742) );
  XNOR2_X1 U623 ( .A(KEYINPUT76), .B(KEYINPUT13), .ZN(n620) );
  XNOR2_X1 U624 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X1 U625 ( .A1(G651), .A2(n595), .ZN(n832) );
  XOR2_X1 U626 ( .A(KEYINPUT17), .B(n555), .Z(n632) );
  NAND2_X1 U627 ( .A1(n556), .A2(G138), .ZN(n558) );
  NAND2_X1 U628 ( .A1(n626), .A2(G102), .ZN(n557) );
  NAND2_X1 U629 ( .A1(n558), .A2(n557), .ZN(n565) );
  AND2_X1 U630 ( .A1(G2104), .A2(G2105), .ZN(n924) );
  NAND2_X1 U631 ( .A1(G114), .A2(n924), .ZN(n562) );
  NAND2_X1 U632 ( .A1(G126), .A2(n519), .ZN(n561) );
  NAND2_X1 U633 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U634 ( .A(KEYINPUT93), .B(n563), .Z(n564) );
  NOR2_X1 U635 ( .A1(n565), .A2(n564), .ZN(G164) );
  INV_X1 U636 ( .A(G651), .ZN(n570) );
  NOR2_X1 U637 ( .A1(G543), .A2(n570), .ZN(n567) );
  XNOR2_X1 U638 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n566) );
  XNOR2_X1 U639 ( .A(n567), .B(n566), .ZN(n828) );
  NAND2_X1 U640 ( .A1(G64), .A2(n828), .ZN(n569) );
  XOR2_X1 U641 ( .A(G543), .B(KEYINPUT0), .Z(n595) );
  NAND2_X1 U642 ( .A1(G52), .A2(n832), .ZN(n568) );
  NAND2_X1 U643 ( .A1(n569), .A2(n568), .ZN(n575) );
  NAND2_X1 U644 ( .A1(G77), .A2(n829), .ZN(n572) );
  NAND2_X1 U645 ( .A1(G90), .A2(n827), .ZN(n571) );
  NAND2_X1 U646 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U647 ( .A(KEYINPUT9), .B(n573), .Z(n574) );
  NOR2_X1 U648 ( .A1(n575), .A2(n574), .ZN(G171) );
  NAND2_X1 U649 ( .A1(n827), .A2(G89), .ZN(n576) );
  XNOR2_X1 U650 ( .A(n576), .B(KEYINPUT4), .ZN(n578) );
  NAND2_X1 U651 ( .A1(G76), .A2(n829), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U653 ( .A(n579), .B(KEYINPUT5), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G63), .A2(n828), .ZN(n581) );
  NAND2_X1 U655 ( .A1(G51), .A2(n832), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U657 ( .A(KEYINPUT6), .B(n582), .Z(n583) );
  NAND2_X1 U658 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U659 ( .A(n585), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U660 ( .A1(n832), .A2(G50), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G62), .A2(n828), .ZN(n587) );
  NAND2_X1 U662 ( .A1(G75), .A2(n829), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n827), .A2(G88), .ZN(n588) );
  XOR2_X1 U665 ( .A(KEYINPUT86), .B(n588), .Z(n589) );
  NOR2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U668 ( .A(KEYINPUT87), .B(n593), .Z(G303) );
  XNOR2_X1 U669 ( .A(G168), .B(KEYINPUT8), .ZN(n594) );
  XNOR2_X1 U670 ( .A(n594), .B(KEYINPUT79), .ZN(G286) );
  NAND2_X1 U671 ( .A1(G49), .A2(n832), .ZN(n597) );
  NAND2_X1 U672 ( .A1(G87), .A2(n595), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U674 ( .A1(n828), .A2(n598), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G74), .A2(G651), .ZN(n599) );
  XOR2_X1 U676 ( .A(KEYINPUT85), .B(n599), .Z(n600) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(G288) );
  NAND2_X1 U678 ( .A1(G61), .A2(n828), .ZN(n603) );
  NAND2_X1 U679 ( .A1(G86), .A2(n827), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n829), .A2(G73), .ZN(n604) );
  XOR2_X1 U682 ( .A(KEYINPUT2), .B(n604), .Z(n605) );
  NOR2_X1 U683 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n832), .A2(G48), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(G305) );
  AND2_X1 U686 ( .A1(n828), .A2(G60), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G72), .A2(n829), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G85), .A2(n827), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n832), .A2(G47), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(G290) );
  NAND2_X1 U693 ( .A1(n828), .A2(G56), .ZN(n615) );
  XOR2_X1 U694 ( .A(KEYINPUT14), .B(n615), .Z(n623) );
  NAND2_X1 U695 ( .A1(n829), .A2(G68), .ZN(n616) );
  XNOR2_X1 U696 ( .A(KEYINPUT75), .B(n616), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n827), .A2(G81), .ZN(n617) );
  XOR2_X1 U698 ( .A(n617), .B(KEYINPUT12), .Z(n618) );
  NOR2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n621) );
  NOR2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n832), .A2(G43), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n1010) );
  XNOR2_X1 U703 ( .A(n628), .B(n627), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n926), .A2(G125), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n631), .B(KEYINPUT67), .ZN(n637) );
  NAND2_X1 U707 ( .A1(G137), .A2(n632), .ZN(n634) );
  NAND2_X1 U708 ( .A1(G113), .A2(n924), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U710 ( .A(KEYINPUT68), .B(n635), .Z(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n789), .A2(G40), .ZN(n758) );
  XNOR2_X1 U713 ( .A(n758), .B(KEYINPUT95), .ZN(n639) );
  NOR2_X1 U714 ( .A1(G164), .A2(G1384), .ZN(n759) );
  INV_X1 U715 ( .A(G1996), .ZN(n975) );
  XNOR2_X1 U716 ( .A(n640), .B(KEYINPUT26), .ZN(n642) );
  NAND2_X1 U717 ( .A1(G54), .A2(n832), .ZN(n648) );
  NAND2_X1 U718 ( .A1(G66), .A2(n828), .ZN(n645) );
  NAND2_X1 U719 ( .A1(G79), .A2(n829), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U721 ( .A1(G92), .A2(n827), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n654), .A2(n1015), .ZN(n653) );
  NOR2_X1 U723 ( .A1(n678), .A2(G1348), .ZN(n651) );
  NOR2_X1 U724 ( .A1(G2067), .A2(n681), .ZN(n650) );
  NOR2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n658), .B(n657), .ZN(n671) );
  NAND2_X1 U728 ( .A1(n678), .A2(G2072), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n659), .B(KEYINPUT27), .ZN(n661) );
  INV_X1 U730 ( .A(G1956), .ZN(n1026) );
  NOR2_X1 U731 ( .A1(n1026), .A2(n678), .ZN(n660) );
  NAND2_X1 U732 ( .A1(G78), .A2(n829), .ZN(n663) );
  NAND2_X1 U733 ( .A1(G91), .A2(n827), .ZN(n662) );
  NAND2_X1 U734 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U735 ( .A(KEYINPUT70), .B(n664), .ZN(n668) );
  NAND2_X1 U736 ( .A1(G65), .A2(n828), .ZN(n666) );
  NAND2_X1 U737 ( .A1(G53), .A2(n832), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U740 ( .A(KEYINPUT71), .B(n669), .Z(n1012) );
  NAND2_X1 U741 ( .A1(n672), .A2(n1012), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n675) );
  XOR2_X1 U743 ( .A(n673), .B(KEYINPUT28), .Z(n674) );
  NAND2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n677) );
  INV_X1 U745 ( .A(KEYINPUT29), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(n713) );
  XNOR2_X1 U747 ( .A(G1961), .B(KEYINPUT97), .ZN(n1047) );
  NAND2_X1 U748 ( .A1(n681), .A2(n1047), .ZN(n680) );
  XNOR2_X1 U749 ( .A(KEYINPUT25), .B(G2078), .ZN(n974) );
  NAND2_X1 U750 ( .A1(n678), .A2(n974), .ZN(n679) );
  NAND2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n686) );
  NAND2_X1 U752 ( .A1(n686), .A2(G171), .ZN(n711) );
  NAND2_X1 U753 ( .A1(n713), .A2(n711), .ZN(n696) );
  NOR2_X1 U754 ( .A1(n681), .A2(G2084), .ZN(n704) );
  NOR2_X1 U755 ( .A1(n707), .A2(n704), .ZN(n682) );
  NAND2_X1 U756 ( .A1(n682), .A2(G8), .ZN(n684) );
  XNOR2_X1 U757 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X1 U758 ( .A1(G168), .A2(n685), .ZN(n688) );
  NOR2_X1 U759 ( .A1(G171), .A2(n686), .ZN(n687) );
  XOR2_X1 U760 ( .A(KEYINPUT31), .B(n689), .Z(n708) );
  NOR2_X1 U761 ( .A1(G1971), .A2(n690), .ZN(n692) );
  NOR2_X1 U762 ( .A1(G2090), .A2(n681), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U764 ( .A(KEYINPUT101), .B(n693), .Z(n694) );
  NAND2_X1 U765 ( .A1(n694), .A2(G303), .ZN(n697) );
  AND2_X1 U766 ( .A1(n708), .A2(n697), .ZN(n695) );
  NAND2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n701) );
  INV_X1 U768 ( .A(n697), .ZN(n698) );
  OR2_X1 U769 ( .A1(n698), .A2(G286), .ZN(n699) );
  AND2_X1 U770 ( .A1(n699), .A2(G8), .ZN(n700) );
  NAND2_X1 U771 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U772 ( .A1(G8), .A2(n704), .ZN(n705) );
  XOR2_X1 U773 ( .A(KEYINPUT96), .B(n705), .Z(n706) );
  NOR2_X1 U774 ( .A1(n707), .A2(n706), .ZN(n710) );
  INV_X1 U775 ( .A(n710), .ZN(n709) );
  OR2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n715) );
  AND2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  AND2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n731) );
  NAND2_X1 U780 ( .A1(G288), .A2(G1976), .ZN(n716) );
  XOR2_X1 U781 ( .A(KEYINPUT103), .B(n716), .Z(n1002) );
  INV_X1 U782 ( .A(n1002), .ZN(n717) );
  OR2_X1 U783 ( .A1(n717), .A2(n690), .ZN(n721) );
  INV_X1 U784 ( .A(n721), .ZN(n718) );
  AND2_X1 U785 ( .A1(n731), .A2(n718), .ZN(n719) );
  NAND2_X1 U786 ( .A1(n730), .A2(n719), .ZN(n723) );
  NOR2_X1 U787 ( .A1(G1976), .A2(G288), .ZN(n725) );
  NOR2_X1 U788 ( .A1(G1971), .A2(G303), .ZN(n720) );
  NOR2_X1 U789 ( .A1(n725), .A2(n720), .ZN(n999) );
  OR2_X1 U790 ( .A1(n721), .A2(n999), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U792 ( .A1(n725), .A2(KEYINPUT33), .ZN(n726) );
  XNOR2_X1 U793 ( .A(n727), .B(KEYINPUT105), .ZN(n729) );
  XOR2_X1 U794 ( .A(G1981), .B(G305), .Z(n1004) );
  INV_X1 U795 ( .A(n1004), .ZN(n728) );
  NAND2_X1 U796 ( .A1(n730), .A2(n731), .ZN(n734) );
  NOR2_X1 U797 ( .A1(G2090), .A2(G303), .ZN(n732) );
  NAND2_X1 U798 ( .A1(G8), .A2(n732), .ZN(n733) );
  NAND2_X1 U799 ( .A1(n734), .A2(n733), .ZN(n735) );
  AND2_X1 U800 ( .A1(n735), .A2(n690), .ZN(n739) );
  NOR2_X1 U801 ( .A1(G1981), .A2(G305), .ZN(n736) );
  XOR2_X1 U802 ( .A(n736), .B(KEYINPUT24), .Z(n737) );
  NOR2_X1 U803 ( .A1(n690), .A2(n737), .ZN(n738) );
  OR2_X1 U804 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U805 ( .A1(G107), .A2(n924), .ZN(n744) );
  NAND2_X1 U806 ( .A1(G95), .A2(n626), .ZN(n743) );
  NAND2_X1 U807 ( .A1(n744), .A2(n743), .ZN(n748) );
  NAND2_X1 U808 ( .A1(G119), .A2(n519), .ZN(n746) );
  NAND2_X1 U809 ( .A1(G131), .A2(n556), .ZN(n745) );
  NAND2_X1 U810 ( .A1(n746), .A2(n745), .ZN(n747) );
  OR2_X1 U811 ( .A1(n748), .A2(n747), .ZN(n901) );
  AND2_X1 U812 ( .A1(n901), .A2(G1991), .ZN(n757) );
  NAND2_X1 U813 ( .A1(G117), .A2(n924), .ZN(n750) );
  NAND2_X1 U814 ( .A1(G129), .A2(n519), .ZN(n749) );
  NAND2_X1 U815 ( .A1(n750), .A2(n749), .ZN(n753) );
  NAND2_X1 U816 ( .A1(n626), .A2(G105), .ZN(n751) );
  XOR2_X1 U817 ( .A(KEYINPUT38), .B(n751), .Z(n752) );
  NOR2_X1 U818 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U819 ( .A1(n556), .A2(G141), .ZN(n754) );
  NAND2_X1 U820 ( .A1(n755), .A2(n754), .ZN(n905) );
  AND2_X1 U821 ( .A1(G1996), .A2(n905), .ZN(n756) );
  NOR2_X1 U822 ( .A1(n757), .A2(n756), .ZN(n960) );
  NOR2_X1 U823 ( .A1(n759), .A2(n758), .ZN(n785) );
  INV_X1 U824 ( .A(n785), .ZN(n760) );
  NOR2_X1 U825 ( .A1(n960), .A2(n760), .ZN(n777) );
  XNOR2_X1 U826 ( .A(G1986), .B(G290), .ZN(n1001) );
  AND2_X1 U827 ( .A1(n1001), .A2(n785), .ZN(n772) );
  NAND2_X1 U828 ( .A1(G104), .A2(n626), .ZN(n762) );
  NAND2_X1 U829 ( .A1(G140), .A2(n556), .ZN(n761) );
  NAND2_X1 U830 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U831 ( .A(KEYINPUT34), .B(n763), .ZN(n768) );
  NAND2_X1 U832 ( .A1(G116), .A2(n924), .ZN(n765) );
  NAND2_X1 U833 ( .A1(G128), .A2(n519), .ZN(n764) );
  NAND2_X1 U834 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U835 ( .A(KEYINPUT35), .B(n766), .Z(n767) );
  NOR2_X1 U836 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U837 ( .A(KEYINPUT36), .B(n769), .Z(n919) );
  XOR2_X1 U838 ( .A(G2067), .B(KEYINPUT37), .Z(n782) );
  AND2_X1 U839 ( .A1(n919), .A2(n782), .ZN(n969) );
  NAND2_X1 U840 ( .A1(n785), .A2(n969), .ZN(n770) );
  XNOR2_X1 U841 ( .A(KEYINPUT94), .B(n770), .ZN(n780) );
  INV_X1 U842 ( .A(n780), .ZN(n771) );
  OR2_X1 U843 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U844 ( .A1(n777), .A2(n773), .ZN(n774) );
  NOR2_X1 U845 ( .A1(G1996), .A2(n905), .ZN(n962) );
  NOR2_X1 U846 ( .A1(G1986), .A2(G290), .ZN(n775) );
  NOR2_X1 U847 ( .A1(G1991), .A2(n901), .ZN(n958) );
  NOR2_X1 U848 ( .A1(n775), .A2(n958), .ZN(n776) );
  NOR2_X1 U849 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U850 ( .A1(n962), .A2(n778), .ZN(n779) );
  XNOR2_X1 U851 ( .A(n779), .B(KEYINPUT39), .ZN(n781) );
  NAND2_X1 U852 ( .A1(n781), .A2(n780), .ZN(n784) );
  NOR2_X1 U853 ( .A1(n782), .A2(n919), .ZN(n783) );
  XNOR2_X1 U854 ( .A(n783), .B(KEYINPUT107), .ZN(n948) );
  NAND2_X1 U855 ( .A1(n784), .A2(n948), .ZN(n786) );
  NAND2_X1 U856 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U857 ( .A(n788), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U858 ( .A(G2438), .B(G2454), .Z(n791) );
  XNOR2_X1 U859 ( .A(G2435), .B(G2430), .ZN(n790) );
  XNOR2_X1 U860 ( .A(n791), .B(n790), .ZN(n792) );
  XOR2_X1 U861 ( .A(n792), .B(G2427), .Z(n794) );
  XNOR2_X1 U862 ( .A(G1348), .B(G1341), .ZN(n793) );
  XNOR2_X1 U863 ( .A(n794), .B(n793), .ZN(n798) );
  XOR2_X1 U864 ( .A(G2443), .B(G2446), .Z(n796) );
  XNOR2_X1 U865 ( .A(KEYINPUT108), .B(G2451), .ZN(n795) );
  XNOR2_X1 U866 ( .A(n796), .B(n795), .ZN(n797) );
  XOR2_X1 U867 ( .A(n798), .B(n797), .Z(n799) );
  AND2_X1 U868 ( .A1(G14), .A2(n799), .ZN(G401) );
  AND2_X1 U869 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U870 ( .A(G120), .ZN(G236) );
  INV_X1 U871 ( .A(G108), .ZN(G238) );
  INV_X1 U872 ( .A(G132), .ZN(G219) );
  INV_X1 U873 ( .A(G82), .ZN(G220) );
  NAND2_X1 U874 ( .A1(G7), .A2(G661), .ZN(n800) );
  XNOR2_X1 U875 ( .A(n800), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U876 ( .A(G567), .ZN(n860) );
  NOR2_X1 U877 ( .A1(G223), .A2(n860), .ZN(n802) );
  XNOR2_X1 U878 ( .A(KEYINPUT74), .B(KEYINPUT11), .ZN(n801) );
  XNOR2_X1 U879 ( .A(n802), .B(n801), .ZN(G234) );
  INV_X1 U880 ( .A(G860), .ZN(n808) );
  OR2_X1 U881 ( .A1(n1010), .A2(n808), .ZN(G153) );
  NAND2_X1 U882 ( .A1(G171), .A2(G868), .ZN(n804) );
  INV_X1 U883 ( .A(G868), .ZN(n844) );
  NAND2_X1 U884 ( .A1(n1015), .A2(n844), .ZN(n803) );
  NAND2_X1 U885 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U886 ( .A(KEYINPUT78), .B(n805), .Z(G284) );
  XOR2_X1 U887 ( .A(n1012), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U888 ( .A1(G299), .A2(G868), .ZN(n807) );
  NOR2_X1 U889 ( .A1(G286), .A2(n844), .ZN(n806) );
  NOR2_X1 U890 ( .A1(n807), .A2(n806), .ZN(G297) );
  NAND2_X1 U891 ( .A1(n808), .A2(G559), .ZN(n809) );
  NAND2_X1 U892 ( .A1(n809), .A2(n1015), .ZN(n810) );
  XNOR2_X1 U893 ( .A(n810), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U894 ( .A1(G868), .A2(n1010), .ZN(n811) );
  XNOR2_X1 U895 ( .A(KEYINPUT80), .B(n811), .ZN(n814) );
  NAND2_X1 U896 ( .A1(G868), .A2(n1015), .ZN(n812) );
  NOR2_X1 U897 ( .A1(G559), .A2(n812), .ZN(n813) );
  NOR2_X1 U898 ( .A1(n814), .A2(n813), .ZN(G282) );
  NAND2_X1 U899 ( .A1(G111), .A2(n924), .ZN(n816) );
  NAND2_X1 U900 ( .A1(G99), .A2(n626), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n816), .A2(n815), .ZN(n822) );
  NAND2_X1 U902 ( .A1(G123), .A2(n519), .ZN(n817) );
  XNOR2_X1 U903 ( .A(n817), .B(KEYINPUT18), .ZN(n820) );
  NAND2_X1 U904 ( .A1(G135), .A2(n556), .ZN(n818) );
  XOR2_X1 U905 ( .A(KEYINPUT81), .B(n818), .Z(n819) );
  NAND2_X1 U906 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U907 ( .A1(n822), .A2(n821), .ZN(n957) );
  XNOR2_X1 U908 ( .A(n957), .B(G2096), .ZN(n824) );
  INV_X1 U909 ( .A(G2100), .ZN(n823) );
  NAND2_X1 U910 ( .A1(n824), .A2(n823), .ZN(G156) );
  INV_X1 U911 ( .A(G303), .ZN(G166) );
  NAND2_X1 U912 ( .A1(G559), .A2(n1015), .ZN(n825) );
  XOR2_X1 U913 ( .A(n1010), .B(n825), .Z(n869) );
  XNOR2_X1 U914 ( .A(G166), .B(KEYINPUT19), .ZN(n826) );
  XNOR2_X1 U915 ( .A(n826), .B(G288), .ZN(n842) );
  NAND2_X1 U916 ( .A1(G93), .A2(n827), .ZN(n837) );
  NAND2_X1 U917 ( .A1(G67), .A2(n828), .ZN(n831) );
  NAND2_X1 U918 ( .A1(G80), .A2(n829), .ZN(n830) );
  NAND2_X1 U919 ( .A1(n831), .A2(n830), .ZN(n835) );
  NAND2_X1 U920 ( .A1(G55), .A2(n832), .ZN(n833) );
  XNOR2_X1 U921 ( .A(KEYINPUT83), .B(n833), .ZN(n834) );
  NOR2_X1 U922 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U923 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U924 ( .A(n838), .B(KEYINPUT84), .ZN(n872) );
  XNOR2_X1 U925 ( .A(n872), .B(G290), .ZN(n839) );
  XNOR2_X1 U926 ( .A(n839), .B(G305), .ZN(n840) );
  XOR2_X1 U927 ( .A(G299), .B(n840), .Z(n841) );
  XNOR2_X1 U928 ( .A(n842), .B(n841), .ZN(n935) );
  XNOR2_X1 U929 ( .A(n869), .B(n935), .ZN(n843) );
  NAND2_X1 U930 ( .A1(n843), .A2(G868), .ZN(n846) );
  NAND2_X1 U931 ( .A1(n844), .A2(n872), .ZN(n845) );
  NAND2_X1 U932 ( .A1(n846), .A2(n845), .ZN(G295) );
  NAND2_X1 U933 ( .A1(G2078), .A2(G2084), .ZN(n848) );
  XOR2_X1 U934 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n847) );
  XNOR2_X1 U935 ( .A(n848), .B(n847), .ZN(n849) );
  NAND2_X1 U936 ( .A1(G2090), .A2(n849), .ZN(n850) );
  XNOR2_X1 U937 ( .A(KEYINPUT21), .B(n850), .ZN(n851) );
  NAND2_X1 U938 ( .A1(n851), .A2(G2072), .ZN(G158) );
  XOR2_X1 U939 ( .A(KEYINPUT89), .B(G44), .Z(n852) );
  XNOR2_X1 U940 ( .A(KEYINPUT3), .B(n852), .ZN(G218) );
  XNOR2_X1 U941 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  NOR2_X1 U942 ( .A1(G220), .A2(G219), .ZN(n853) );
  XOR2_X1 U943 ( .A(KEYINPUT22), .B(n853), .Z(n854) );
  NOR2_X1 U944 ( .A1(G218), .A2(n854), .ZN(n855) );
  XNOR2_X1 U945 ( .A(KEYINPUT90), .B(n855), .ZN(n856) );
  NAND2_X1 U946 ( .A1(n856), .A2(G96), .ZN(n873) );
  NAND2_X1 U947 ( .A1(G2106), .A2(n873), .ZN(n857) );
  XNOR2_X1 U948 ( .A(n857), .B(KEYINPUT91), .ZN(n862) );
  NOR2_X1 U949 ( .A1(G236), .A2(G237), .ZN(n858) );
  NAND2_X1 U950 ( .A1(G69), .A2(n858), .ZN(n859) );
  NOR2_X1 U951 ( .A1(G238), .A2(n859), .ZN(n875) );
  NOR2_X1 U952 ( .A1(n860), .A2(n875), .ZN(n861) );
  NOR2_X1 U953 ( .A1(n862), .A2(n861), .ZN(G319) );
  INV_X1 U954 ( .A(G319), .ZN(n942) );
  NAND2_X1 U955 ( .A1(G661), .A2(G483), .ZN(n863) );
  XNOR2_X1 U956 ( .A(KEYINPUT92), .B(n863), .ZN(n864) );
  NOR2_X1 U957 ( .A1(n942), .A2(n864), .ZN(n868) );
  NAND2_X1 U958 ( .A1(n868), .A2(G36), .ZN(G176) );
  INV_X1 U959 ( .A(G223), .ZN(n865) );
  NAND2_X1 U960 ( .A1(G2106), .A2(n865), .ZN(G217) );
  AND2_X1 U961 ( .A1(G15), .A2(G2), .ZN(n866) );
  NAND2_X1 U962 ( .A1(G661), .A2(n866), .ZN(G259) );
  NAND2_X1 U963 ( .A1(G3), .A2(G1), .ZN(n867) );
  NAND2_X1 U964 ( .A1(n868), .A2(n867), .ZN(G188) );
  XNOR2_X1 U965 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  XOR2_X1 U967 ( .A(n869), .B(KEYINPUT82), .Z(n870) );
  NOR2_X1 U968 ( .A1(G860), .A2(n870), .ZN(n871) );
  XOR2_X1 U969 ( .A(n872), .B(n871), .Z(G145) );
  INV_X1 U970 ( .A(G96), .ZN(G221) );
  INV_X1 U971 ( .A(n873), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(G261) );
  INV_X1 U973 ( .A(G261), .ZN(G325) );
  XOR2_X1 U974 ( .A(G2100), .B(G2096), .Z(n877) );
  XNOR2_X1 U975 ( .A(KEYINPUT42), .B(G2678), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(n881) );
  XOR2_X1 U977 ( .A(KEYINPUT43), .B(G2072), .Z(n879) );
  XNOR2_X1 U978 ( .A(G2067), .B(G2090), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U980 ( .A(n881), .B(n880), .Z(n883) );
  XNOR2_X1 U981 ( .A(G2078), .B(G2084), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(G227) );
  XNOR2_X1 U983 ( .A(G1956), .B(G2474), .ZN(n893) );
  XOR2_X1 U984 ( .A(G1981), .B(G1966), .Z(n885) );
  XNOR2_X1 U985 ( .A(G1986), .B(G1961), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n889) );
  XOR2_X1 U987 ( .A(G1976), .B(G1971), .Z(n887) );
  XNOR2_X1 U988 ( .A(G1996), .B(G1991), .ZN(n886) );
  XNOR2_X1 U989 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U990 ( .A(n889), .B(n888), .Z(n891) );
  XNOR2_X1 U991 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(G229) );
  NAND2_X1 U994 ( .A1(G112), .A2(n924), .ZN(n895) );
  NAND2_X1 U995 ( .A1(G136), .A2(n556), .ZN(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n900) );
  NAND2_X1 U997 ( .A1(n519), .A2(G124), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n896), .B(KEYINPUT44), .ZN(n898) );
  NAND2_X1 U999 ( .A1(G100), .A2(n626), .ZN(n897) );
  NAND2_X1 U1000 ( .A1(n898), .A2(n897), .ZN(n899) );
  NOR2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(G162) );
  XOR2_X1 U1002 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n903) );
  XOR2_X1 U1003 ( .A(n901), .B(KEYINPUT114), .Z(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1005 ( .A(n904), .B(n957), .Z(n907) );
  XOR2_X1 U1006 ( .A(n905), .B(G162), .Z(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(n556), .A2(G142), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n908), .B(KEYINPUT112), .ZN(n910) );
  NAND2_X1 U1010 ( .A1(G106), .A2(n626), .ZN(n909) );
  NAND2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n911), .B(KEYINPUT45), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(G118), .A2(n924), .ZN(n912) );
  NAND2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(G130), .A2(n519), .ZN(n914) );
  XNOR2_X1 U1016 ( .A(KEYINPUT111), .B(n914), .ZN(n915) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1018 ( .A(n918), .B(n917), .Z(n921) );
  XNOR2_X1 U1019 ( .A(G160), .B(n919), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(n921), .B(n920), .ZN(n933) );
  NAND2_X1 U1021 ( .A1(G103), .A2(n626), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(G139), .A2(n556), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n931) );
  NAND2_X1 U1024 ( .A1(n924), .A2(G115), .ZN(n925) );
  XOR2_X1 U1025 ( .A(KEYINPUT113), .B(n925), .Z(n928) );
  NAND2_X1 U1026 ( .A1(n519), .A2(G127), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1028 ( .A(KEYINPUT47), .B(n929), .Z(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n950) );
  XNOR2_X1 U1030 ( .A(n950), .B(G164), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n933), .B(n932), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(G37), .A2(n934), .ZN(G395) );
  XNOR2_X1 U1033 ( .A(n1010), .B(n935), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(G171), .B(n1015), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(n937), .B(n936), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n938), .B(G286), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(G37), .A2(n939), .ZN(G397) );
  XNOR2_X1 U1038 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(G227), .A2(G229), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(n941), .B(n940), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(G401), .A2(n942), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(KEYINPUT115), .B(n943), .ZN(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(G395), .A2(G397), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(G225) );
  INV_X1 U1046 ( .A(G225), .ZN(G308) );
  INV_X1 U1047 ( .A(KEYINPUT55), .ZN(n994) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n971) );
  XNOR2_X1 U1049 ( .A(G2084), .B(G160), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(G2072), .B(n950), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(G164), .B(G2078), .ZN(n951) );
  NAND2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1054 ( .A(KEYINPUT117), .B(n953), .Z(n954) );
  XNOR2_X1 U1055 ( .A(KEYINPUT50), .B(n954), .ZN(n955) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n967) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n965) );
  XOR2_X1 U1059 ( .A(G2090), .B(G162), .Z(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(n963), .B(KEYINPUT51), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n971), .B(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n994), .A2(n972), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n973), .A2(G29), .ZN(n1058) );
  XNOR2_X1 U1068 ( .A(G2090), .B(G35), .ZN(n989) );
  XNOR2_X1 U1069 ( .A(n974), .B(G27), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n975), .B(G32), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(G2067), .B(G26), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G2072), .B(G33), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n980), .B(KEYINPUT119), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT120), .B(n983), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n984), .A2(G28), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G25), .B(G1991), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(KEYINPUT53), .B(n987), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n992) );
  XOR2_X1 U1083 ( .A(G2084), .B(KEYINPUT54), .Z(n990) );
  XNOR2_X1 U1084 ( .A(G34), .B(n990), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n994), .B(n993), .ZN(n996) );
  INV_X1 U1087 ( .A(G29), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(G11), .A2(n997), .ZN(n1056) );
  XNOR2_X1 U1090 ( .A(G16), .B(KEYINPUT56), .ZN(n1024) );
  NAND2_X1 U1091 ( .A1(G1971), .A2(G303), .ZN(n998) );
  NAND2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G168), .B(G1966), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(n1006), .B(KEYINPUT121), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(n1007), .B(KEYINPUT57), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1022) );
  XNOR2_X1 U1100 ( .A(G1341), .B(KEYINPUT123), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(n1011), .B(n1010), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(n1012), .B(G1956), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(G1348), .B(n1015), .Z(n1017) );
  XOR2_X1 U1105 ( .A(G171), .B(G1961), .Z(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(KEYINPUT122), .B(n1018), .Z(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1054) );
  INV_X1 U1111 ( .A(G16), .ZN(n1052) );
  XNOR2_X1 U1112 ( .A(KEYINPUT127), .B(G1966), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(n1025), .B(G21), .ZN(n1046) );
  XNOR2_X1 U1114 ( .A(n1026), .B(G20), .ZN(n1034) );
  XOR2_X1 U1115 ( .A(G1981), .B(G6), .Z(n1029) );
  XOR2_X1 U1116 ( .A(G19), .B(KEYINPUT124), .Z(n1027) );
  XNOR2_X1 U1117 ( .A(G1341), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1032) );
  XOR2_X1 U1119 ( .A(KEYINPUT59), .B(G1348), .Z(n1030) );
  XNOR2_X1 U1120 ( .A(G4), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1121 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1122 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1123 ( .A(n1035), .B(KEYINPUT126), .ZN(n1037) );
  XOR2_X1 U1124 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n1036) );
  XNOR2_X1 U1125 ( .A(n1037), .B(n1036), .ZN(n1044) );
  XNOR2_X1 U1126 ( .A(G1971), .B(G22), .ZN(n1039) );
  XNOR2_X1 U1127 ( .A(G23), .B(G1976), .ZN(n1038) );
  NOR2_X1 U1128 ( .A1(n1039), .A2(n1038), .ZN(n1041) );
  XOR2_X1 U1129 ( .A(G1986), .B(G24), .Z(n1040) );
  NAND2_X1 U1130 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1131 ( .A(KEYINPUT58), .B(n1042), .ZN(n1043) );
  NOR2_X1 U1132 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NAND2_X1 U1133 ( .A1(n1046), .A2(n1045), .ZN(n1049) );
  XOR2_X1 U1134 ( .A(G5), .B(n1047), .Z(n1048) );
  NOR2_X1 U1135 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XNOR2_X1 U1136 ( .A(KEYINPUT61), .B(n1050), .ZN(n1051) );
  NAND2_X1 U1137 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  NAND2_X1 U1138 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  NOR2_X1 U1139 ( .A1(n1056), .A2(n1055), .ZN(n1057) );
  NAND2_X1 U1140 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
  XOR2_X1 U1141 ( .A(KEYINPUT62), .B(n1059), .Z(G311) );
  INV_X1 U1142 ( .A(G311), .ZN(G150) );
  INV_X1 U1143 ( .A(G171), .ZN(G301) );
endmodule

