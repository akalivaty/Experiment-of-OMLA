//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(G122), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G122), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  XNOR2_X1  g008(.A(G128), .B(G143), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n193), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n189), .A2(KEYINPUT14), .A3(G122), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n188), .A2(new_n190), .ZN(new_n199));
  OAI211_X1 g013(.A(G107), .B(new_n198), .C1(new_n199), .C2(KEYINPUT14), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n197), .B(new_n200), .C1(new_n194), .C2(new_n196), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT9), .B(G234), .ZN(new_n202));
  INV_X1    g016(.A(G217), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n202), .A2(new_n203), .A3(G953), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT87), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n191), .B1(new_n188), .B2(new_n190), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n193), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n206), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(new_n192), .A3(KEYINPUT87), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT88), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  OAI22_X1  g025(.A1(new_n210), .A2(KEYINPUT13), .B1(new_n211), .B2(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(KEYINPUT13), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(G134), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(new_n196), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT13), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT88), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n213), .B(new_n218), .C1(G128), .C2(new_n211), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n195), .B1(new_n219), .B2(G134), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n207), .B(new_n209), .C1(new_n216), .C2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n221), .A2(KEYINPUT89), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(KEYINPUT89), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n201), .B(new_n204), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT90), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n221), .B(KEYINPUT89), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT90), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n201), .A4(new_n204), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n201), .B1(new_n222), .B2(new_n223), .ZN(new_n229));
  INV_X1    g043(.A(new_n204), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n225), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G902), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT15), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G478), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n235), .B1(new_n232), .B2(new_n233), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G475), .ZN(new_n240));
  XNOR2_X1  g054(.A(G113), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(G104), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G140), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G125), .ZN(new_n246));
  INV_X1    g060(.A(G125), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G140), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT76), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT76), .ZN(new_n252));
  INV_X1    g066(.A(G146), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT75), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n246), .A2(new_n248), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n247), .A2(KEYINPUT75), .A3(G140), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(G146), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT18), .A2(G131), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G237), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(G214), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(KEYINPUT83), .B2(new_n211), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT83), .B(G143), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n259), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n262), .A2(new_n263), .A3(G214), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n211), .A2(KEYINPUT83), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n211), .A2(KEYINPUT83), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n265), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n272), .B2(new_n265), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n261), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT85), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n267), .A2(KEYINPUT84), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n274), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n261), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n268), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n267), .A2(G131), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT17), .ZN(new_n285));
  INV_X1    g099(.A(G131), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n272), .A2(new_n286), .A3(new_n265), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n256), .A2(KEYINPUT16), .A3(new_n257), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT16), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n246), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n253), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n253), .B1(new_n289), .B2(new_n291), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n286), .B1(new_n272), .B2(new_n265), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT17), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n288), .A2(new_n292), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n244), .B1(new_n283), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n268), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n281), .B1(new_n280), .B2(new_n261), .ZN(new_n301));
  AOI211_X1 g115(.A(KEYINPUT85), .B(new_n260), .C1(new_n279), .C2(new_n274), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n243), .A3(new_n297), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n240), .B1(new_n305), .B2(new_n233), .ZN(new_n306));
  NOR2_X1   g120(.A1(G475), .A2(G902), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n283), .A2(new_n244), .A3(new_n298), .ZN(new_n308));
  INV_X1    g122(.A(new_n287), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n294), .B1(new_n309), .B2(new_n295), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT19), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n251), .A2(new_n252), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n256), .A2(KEYINPUT19), .A3(new_n257), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n253), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n313), .A2(KEYINPUT86), .A3(new_n253), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n311), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n243), .B1(new_n303), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n307), .B1(new_n308), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT20), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n244), .B1(new_n283), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n304), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT20), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n307), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n306), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(G234), .A2(G237), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G952), .A3(new_n263), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT91), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT21), .B(G898), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT92), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(G902), .A3(G953), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n239), .A2(new_n329), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G110), .B(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n263), .A2(G227), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n338), .B(new_n339), .Z(new_n340));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n242), .B2(G107), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n191), .A2(KEYINPUT3), .A3(G104), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G101), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n242), .A2(G107), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT79), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n242), .A3(G107), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n344), .A2(new_n345), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n346), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n242), .A2(G107), .ZN(new_n352));
  OAI21_X1  g166(.A(G101), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G143), .B(G146), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT1), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G128), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT67), .ZN(new_n360));
  INV_X1    g174(.A(G128), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n211), .A2(G146), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n253), .A2(G143), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(KEYINPUT1), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n253), .A2(G143), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n211), .A2(G146), .ZN(new_n368));
  AOI21_X1  g182(.A(G128), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n358), .A2(new_n253), .A3(G143), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n369), .A2(KEYINPUT67), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n359), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n350), .A3(new_n353), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n356), .A2(new_n372), .B1(new_n374), .B2(new_n355), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n286), .A2(KEYINPUT66), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT11), .B1(new_n194), .B2(G137), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT11), .ZN(new_n378));
  INV_X1    g192(.A(G137), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G134), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT65), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n379), .B2(G134), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n194), .A2(KEYINPUT65), .A3(G137), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n376), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n194), .A2(KEYINPUT65), .A3(G137), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT65), .B1(new_n194), .B2(G137), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n377), .A2(new_n380), .ZN(new_n390));
  INV_X1    g204(.A(new_n376), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  INV_X1    g209(.A(new_n344), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n347), .A2(new_n349), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n395), .B(G101), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT0), .A2(G128), .ZN(new_n399));
  OR2_X1    g213(.A1(KEYINPUT0), .A2(G128), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n399), .B(new_n400), .C1(new_n362), .C2(new_n363), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT0), .A4(G128), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n396), .A2(new_n397), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(new_n345), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n350), .A2(KEYINPUT4), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n398), .B(new_n403), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n375), .A2(new_n394), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n394), .B1(new_n375), .B2(new_n407), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n340), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n357), .A2(new_n358), .A3(G128), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT67), .B1(new_n369), .B2(new_n370), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n365), .B(new_n360), .C1(new_n357), .C2(G128), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n354), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n394), .B1(new_n416), .B2(new_n374), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(KEYINPUT80), .A2(KEYINPUT12), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n340), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n419), .A2(new_n421), .A3(new_n408), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n411), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G469), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n233), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n233), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n419), .A2(new_n408), .A3(new_n421), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n340), .ZN(new_n430));
  OR3_X1    g244(.A1(new_n409), .A2(new_n410), .A3(new_n340), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n431), .A3(G469), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n426), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G221), .B1(new_n202), .B2(G902), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G214), .B1(G237), .B2(G902), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n415), .A2(new_n247), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n247), .B2(new_n403), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n263), .A2(G224), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT7), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n354), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT2), .B(G113), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G116), .B(G119), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G119), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n450), .A3(G116), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G113), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n446), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n442), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT8), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT81), .B1(new_n449), .B2(new_n452), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n452), .B1(KEYINPUT5), .B2(new_n445), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT81), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n446), .A3(new_n460), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n454), .B(new_n456), .C1(new_n461), .C2(new_n442), .ZN(new_n462));
  INV_X1    g276(.A(new_n440), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n437), .B(new_n463), .C1(new_n247), .C2(new_n403), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n441), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n442), .A2(new_n457), .A3(new_n460), .A4(new_n446), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n398), .B1(new_n405), .B2(new_n406), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n447), .A2(new_n443), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n446), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n446), .A3(KEYINPUT68), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n455), .B(new_n466), .C1(new_n467), .C2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n465), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n466), .B1(new_n467), .B2(new_n473), .ZN(new_n476));
  INV_X1    g290(.A(new_n455), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(KEYINPUT6), .A3(new_n474), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n439), .B(KEYINPUT82), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n438), .B(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n476), .A2(new_n482), .A3(new_n477), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G210), .B1(G237), .B2(G902), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n475), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n485), .B1(new_n475), .B2(new_n484), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n436), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n337), .A2(new_n435), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(G472), .A2(G902), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n381), .A2(new_n385), .A3(new_n376), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n391), .B1(new_n389), .B2(new_n390), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n403), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT69), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n390), .A2(new_n383), .A3(new_n384), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n286), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n194), .A2(G137), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n379), .A2(G134), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n497), .A2(new_n498), .A3(new_n286), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n372), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT69), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n393), .A2(new_n503), .A3(new_n403), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n494), .A2(new_n502), .A3(new_n473), .A4(new_n504), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n506));
  NAND3_X1  g320(.A1(new_n262), .A2(new_n263), .A3(G210), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(G101), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT64), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n401), .A2(new_n514), .A3(new_n402), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n401), .A2(new_n402), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT64), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n393), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n499), .B1(new_n495), .B2(new_n286), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n415), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n513), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n494), .A2(new_n502), .A3(KEYINPUT30), .A4(new_n504), .ZN(new_n522));
  INV_X1    g336(.A(new_n473), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n512), .A2(new_n524), .A3(KEYINPUT71), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT71), .B1(new_n512), .B2(new_n524), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n510), .B(KEYINPUT72), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n523), .B1(new_n518), .B2(new_n520), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(new_n505), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n473), .A2(new_n493), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT28), .B1(new_n533), .B2(new_n502), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n529), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n512), .A2(new_n524), .A3(new_n527), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n490), .B1(new_n528), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT32), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n490), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(new_n539), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n528), .B2(new_n537), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT73), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT29), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n524), .A2(new_n505), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n510), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n532), .A2(new_n534), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n545), .B(new_n547), .C1(new_n548), .C2(new_n529), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n494), .A2(new_n502), .A3(new_n504), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n523), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n530), .B1(new_n551), .B2(new_n505), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n534), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n510), .A2(new_n545), .ZN(new_n554));
  AOI21_X1  g368(.A(G902), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G472), .ZN(new_n557));
  INV_X1    g371(.A(new_n537), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n512), .A2(new_n524), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT71), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n512), .A2(new_n524), .A3(KEYINPUT71), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(KEYINPUT31), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT73), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n542), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n540), .A2(new_n544), .A3(new_n557), .A4(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT24), .B(G110), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT74), .ZN(new_n569));
  XNOR2_X1  g383(.A(G119), .B(G128), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT23), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n450), .B2(G128), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n361), .A2(KEYINPUT23), .A3(G119), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n572), .B(new_n573), .C1(G119), .C2(new_n361), .ZN(new_n574));
  OAI22_X1  g388(.A1(new_n569), .A2(new_n570), .B1(G110), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n294), .A3(new_n254), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT74), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n568), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n568), .A2(new_n577), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n570), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n574), .A2(G110), .ZN(new_n581));
  INV_X1    g395(.A(new_n292), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n293), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT77), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n576), .A2(new_n583), .A3(new_n588), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n233), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT25), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n203), .B1(G234), .B2(new_n233), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n590), .A2(new_n591), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n597), .A2(G902), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n489), .A2(new_n567), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  AOI21_X1  g419(.A(new_n243), .B1(new_n303), .B2(new_n297), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n233), .B1(new_n308), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(G475), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n323), .A2(new_n328), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n232), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n610), .B1(new_n229), .B2(new_n230), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n224), .ZN(new_n613));
  INV_X1    g427(.A(G478), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(G902), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n232), .A2(new_n233), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n614), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n608), .A2(new_n609), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT93), .ZN(new_n620));
  INV_X1    g434(.A(new_n436), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n475), .A2(new_n484), .ZN(new_n622));
  INV_X1    g436(.A(new_n485), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n475), .A2(new_n484), .A3(new_n485), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n619), .A2(new_n620), .A3(new_n336), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n616), .A2(new_n618), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n327), .B1(new_n326), .B2(new_n307), .ZN(new_n629));
  INV_X1    g443(.A(new_n307), .ZN(new_n630));
  AOI211_X1 g444(.A(KEYINPUT20), .B(new_n630), .C1(new_n325), .C2(new_n304), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n608), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n336), .B(new_n436), .C1(new_n486), .C2(new_n487), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT93), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n541), .B1(new_n558), .B2(new_n563), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n233), .B1(new_n528), .B2(new_n537), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n638), .B2(G472), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n435), .A2(new_n602), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n636), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  INV_X1    g457(.A(new_n238), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n236), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n329), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n336), .B(KEYINPUT94), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n436), .B(new_n647), .C1(new_n486), .C2(new_n487), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(new_n639), .A3(new_n640), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  INV_X1    g466(.A(new_n337), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n584), .A2(KEYINPUT95), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT95), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n576), .A2(new_n583), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(KEYINPUT36), .B2(new_n589), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n589), .A2(KEYINPUT36), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n654), .A2(new_n659), .A3(new_n656), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n600), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n598), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n488), .ZN(new_n665));
  INV_X1    g479(.A(new_n435), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n653), .A2(new_n665), .A3(new_n639), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  OR2_X1    g483(.A1(new_n335), .A2(G900), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n332), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n646), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n567), .A2(new_n666), .A3(new_n665), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NAND2_X1  g488(.A1(new_n544), .A2(new_n566), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n525), .A2(new_n526), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n551), .A2(new_n505), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n529), .ZN(new_n678));
  AOI21_X1  g492(.A(G902), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(G472), .ZN(new_n680));
  OAI22_X1  g494(.A1(new_n637), .A2(KEYINPUT32), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT96), .B1(new_n675), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n561), .A2(new_n562), .A3(new_n678), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n680), .B1(new_n683), .B2(new_n233), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n538), .B2(new_n539), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT96), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n685), .A2(new_n686), .A3(new_n544), .A4(new_n566), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n239), .A2(new_n329), .A3(new_n621), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n664), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT97), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n624), .A2(new_n625), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT38), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n671), .B(new_n696), .Z(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n666), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AND4_X1   g515(.A1(new_n688), .A2(new_n691), .A3(new_n695), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n211), .ZN(G45));
  NOR2_X1   g517(.A1(new_n633), .A2(new_n671), .ZN(new_n704));
  AND4_X1   g518(.A1(new_n567), .A2(new_n666), .A3(new_n665), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n253), .ZN(G48));
  AOI21_X1  g520(.A(new_n565), .B1(new_n564), .B2(new_n542), .ZN(new_n707));
  INV_X1    g521(.A(new_n542), .ZN(new_n708));
  AOI211_X1 g522(.A(KEYINPUT73), .B(new_n708), .C1(new_n558), .C2(new_n563), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n538), .A2(new_n539), .B1(new_n556), .B2(G472), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n602), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(KEYINPUT99), .A2(G469), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n424), .B2(new_n233), .ZN(new_n714));
  INV_X1    g528(.A(new_n713), .ZN(new_n715));
  AOI211_X1 g529(.A(G902), .B(new_n715), .C1(new_n411), .C2(new_n423), .ZN(new_n716));
  INV_X1    g530(.A(new_n434), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n712), .A2(new_n636), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n567), .A2(new_n603), .A3(new_n649), .A4(new_n718), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT100), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  NAND2_X1  g538(.A1(new_n718), .A2(new_n626), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n239), .A2(new_n663), .A3(new_n329), .A4(new_n336), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(new_n567), .A3(KEYINPUT101), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT101), .B1(new_n727), .B2(new_n567), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT102), .B(G119), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G21));
  NAND2_X1  g546(.A1(new_n638), .A2(G472), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n529), .B1(new_n552), .B2(new_n534), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n536), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n490), .B1(new_n528), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  AND4_X1   g551(.A1(new_n645), .A2(new_n692), .A3(new_n632), .A4(new_n436), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n718), .A2(new_n647), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(new_n603), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  INV_X1    g555(.A(new_n671), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n619), .A2(new_n626), .A3(new_n742), .A4(new_n718), .ZN(new_n743));
  AOI21_X1  g557(.A(G902), .B1(new_n558), .B2(new_n563), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n736), .B(new_n663), .C1(new_n744), .C2(new_n680), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT103), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n733), .A2(new_n747), .A3(new_n663), .A4(new_n736), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n743), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n247), .ZN(G27));
  NOR2_X1   g564(.A1(new_n717), .A2(new_n621), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n624), .A2(new_n625), .A3(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n426), .A2(new_n428), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n430), .A2(KEYINPUT104), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n430), .A2(KEYINPUT104), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n431), .A4(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n752), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n712), .A2(new_n704), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n602), .B1(new_n711), .B2(new_n543), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(KEYINPUT42), .A3(new_n704), .A4(new_n757), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  NAND4_X1  g578(.A1(new_n567), .A2(new_n603), .A3(new_n672), .A4(new_n757), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  INV_X1    g580(.A(KEYINPUT106), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n754), .A2(KEYINPUT45), .A3(new_n431), .A4(new_n755), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT45), .B1(new_n430), .B2(new_n431), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n425), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n427), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n771), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT105), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(KEYINPUT46), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n772), .A2(new_n426), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n434), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n767), .B1(new_n776), .B2(new_n697), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n775), .A2(KEYINPUT106), .A3(new_n434), .A4(new_n698), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT43), .B1(new_n329), .B2(KEYINPUT107), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n628), .A2(new_n329), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n639), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n782), .A3(new_n663), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n624), .A2(new_n436), .A3(new_n625), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n783), .B2(new_n784), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n777), .A2(new_n778), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(KEYINPUT108), .B(G137), .Z(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(G39));
  NAND2_X1  g604(.A1(new_n619), .A2(new_n742), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n567), .A2(new_n791), .A3(new_n603), .A4(new_n786), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n775), .A2(KEYINPUT47), .A3(new_n434), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT47), .B1(new_n775), .B2(new_n434), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  AOI21_X1  g610(.A(KEYINPUT116), .B1(new_n263), .B2(G952), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n263), .A2(KEYINPUT116), .A3(G952), .ZN(new_n798));
  INV_X1    g612(.A(new_n332), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n781), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(new_n603), .A3(new_n737), .ZN(new_n801));
  INV_X1    g615(.A(new_n725), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n797), .B(new_n798), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n714), .A2(new_n716), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n717), .A3(new_n786), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n800), .A2(new_n761), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n808));
  OR2_X1    g622(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n806), .A2(new_n603), .A3(new_n799), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n688), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n633), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n807), .A2(new_n808), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n811), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n694), .A2(new_n621), .A3(new_n718), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT115), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n801), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT50), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n813), .A2(new_n632), .A3(new_n628), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n745), .A2(KEYINPUT103), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n745), .A2(KEYINPUT103), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n800), .B(new_n806), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n821), .A2(KEYINPUT51), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n786), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n801), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n793), .A2(new_n794), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n804), .A2(new_n717), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n816), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n829), .A2(KEYINPUT114), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n830), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n829), .A2(KEYINPUT114), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n827), .B(new_n801), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n822), .A3(new_n825), .A4(new_n821), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n756), .A2(new_n753), .ZN(new_n840));
  INV_X1    g654(.A(new_n752), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n619), .A2(new_n840), .A3(new_n742), .A4(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n824), .B2(new_n823), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT110), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n239), .B2(new_n632), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n645), .A2(KEYINPUT110), .A3(new_n329), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n633), .ZN(new_n847));
  INV_X1    g661(.A(new_n648), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n639), .A3(new_n640), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n843), .A2(new_n604), .A3(new_n667), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n239), .A2(new_n329), .A3(new_n742), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n664), .A3(new_n786), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n567), .A3(new_n666), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n765), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT112), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n849), .A2(new_n604), .A3(new_n667), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n765), .A2(new_n853), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n843), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n760), .B2(new_n762), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n855), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT113), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT100), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n722), .B(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n719), .B(new_n740), .C1(new_n728), .C2(new_n729), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n728), .A2(new_n729), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n627), .A2(new_n635), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n567), .A2(new_n603), .A3(new_n718), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n740), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n723), .A2(new_n868), .A3(new_n872), .A4(KEYINPUT113), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n717), .B(new_n671), .C1(new_n624), .C2(new_n625), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n689), .A2(new_n664), .A3(new_n875), .A4(new_n840), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n682), .B2(new_n687), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n705), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n567), .A2(new_n666), .A3(new_n665), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n749), .B1(new_n879), .B2(new_n672), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT52), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n862), .A2(new_n874), .A3(new_n885), .ZN(new_n886));
  XOR2_X1   g700(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n887));
  INV_X1    g701(.A(new_n743), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n824), .B2(new_n823), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n673), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n890), .A2(new_n877), .A3(new_n882), .A4(new_n705), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT52), .B1(new_n878), .B2(new_n880), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n849), .A2(new_n604), .A3(new_n667), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n704), .A2(new_n757), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n748), .B2(new_n746), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n894), .A2(new_n854), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n730), .A2(new_n871), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n723), .A4(new_n763), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n887), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n886), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n893), .A2(new_n899), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n860), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n887), .B2(new_n903), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n902), .B1(new_n905), .B2(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n839), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT118), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n839), .A2(new_n909), .A3(new_n906), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n908), .B(new_n910), .C1(G952), .C2(G953), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n603), .A2(new_n751), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT109), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n780), .B1(KEYINPUT49), .B2(new_n805), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(KEYINPUT49), .B2(new_n805), .ZN(new_n915));
  OR4_X1    g729(.A1(new_n688), .A2(new_n913), .A3(new_n915), .A4(new_n695), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n916), .ZN(G75));
  NOR2_X1   g731(.A1(new_n263), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n886), .A2(new_n900), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n233), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT56), .B1(new_n921), .B2(G210), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n479), .A2(new_n483), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n481), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT55), .Z(new_n925));
  OAI21_X1  g739(.A(new_n919), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n901), .A2(KEYINPUT119), .A3(G902), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT119), .B1(new_n901), .B2(G902), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n623), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n925), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n926), .B1(new_n931), .B2(new_n933), .ZN(G51));
  NAND2_X1  g748(.A1(new_n768), .A2(new_n770), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n927), .A2(new_n929), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n427), .B(KEYINPUT57), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT121), .B1(new_n901), .B2(KEYINPUT54), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n939), .B(new_n940), .C1(new_n886), .C2(new_n900), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT120), .B1(new_n901), .B2(KEYINPUT54), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n886), .A2(new_n900), .A3(new_n944), .A4(new_n940), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n937), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n936), .B1(new_n947), .B2(new_n424), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT122), .B1(new_n948), .B2(new_n918), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n943), .B(new_n945), .C1(new_n938), .C2(new_n941), .ZN(new_n951));
  AOI22_X1  g765(.A1(new_n951), .A2(new_n937), .B1(new_n411), .B2(new_n423), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n950), .B(new_n919), .C1(new_n952), .C2(new_n936), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n949), .A2(new_n953), .ZN(G54));
  NAND4_X1  g768(.A1(new_n928), .A2(KEYINPUT58), .A3(new_n930), .A4(G475), .ZN(new_n955));
  INV_X1    g769(.A(new_n326), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n955), .A2(KEYINPUT123), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n919), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT123), .B1(new_n955), .B2(new_n956), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G60));
  NAND2_X1  g774(.A1(new_n611), .A2(new_n613), .ZN(new_n961));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT59), .Z(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n906), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n919), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n961), .A2(new_n963), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n951), .B2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n920), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n919), .B1(new_n970), .B2(new_n599), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n661), .B2(new_n970), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g787(.A(new_n263), .B1(new_n334), .B2(G224), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n898), .A2(new_n723), .A3(new_n856), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT124), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n974), .B1(new_n977), .B2(new_n263), .ZN(new_n978));
  INV_X1    g792(.A(G898), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n923), .B1(new_n979), .B2(G953), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n978), .B(new_n980), .ZN(G69));
  NAND2_X1  g795(.A1(new_n788), .A2(new_n795), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n699), .A2(new_n786), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n983), .A2(new_n847), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n982), .B1(new_n712), .B2(new_n984), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n702), .A2(new_n705), .A3(new_n890), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT62), .ZN(new_n987));
  AOI21_X1  g801(.A(G953), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n521), .A2(new_n522), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n313), .A2(new_n314), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n777), .A2(new_n738), .A3(new_n761), .A4(new_n778), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n890), .A2(new_n705), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n994), .A2(new_n763), .A3(new_n765), .A4(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(new_n982), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n263), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n263), .A2(G900), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT126), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  AOI22_X1  g815(.A1(new_n993), .A2(KEYINPUT125), .B1(new_n992), .B2(new_n1001), .ZN(new_n1002));
  OR3_X1    g816(.A1(new_n988), .A2(KEYINPUT125), .A3(new_n992), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n263), .B1(G227), .B2(G900), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1004), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1005), .A2(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  OAI21_X1  g823(.A(new_n1009), .B1(new_n997), .B2(new_n977), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1010), .A2(new_n524), .A3(new_n505), .A4(new_n510), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n676), .A2(new_n547), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1012), .A2(new_n1009), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n918), .B1(new_n905), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n985), .A2(new_n987), .A3(new_n976), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n1009), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n511), .A3(new_n546), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1011), .B(new_n1014), .C1(new_n1017), .C2(KEYINPUT127), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(KEYINPUT127), .B2(new_n1017), .ZN(G57));
endmodule


