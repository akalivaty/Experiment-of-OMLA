//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT0), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n192), .A3(new_n193), .A4(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT0), .A4(G128), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT65), .A2(G137), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT65), .A2(G137), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT11), .A2(G134), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT11), .A2(G134), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT11), .A2(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n203), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(new_n203), .B2(new_n206), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n198), .B(new_n199), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n189), .A2(G146), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n187), .A2(G143), .ZN(new_n215));
  OAI211_X1 g029(.A(G128), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n188), .B(new_n190), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n216), .A2(KEYINPUT67), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT67), .B1(new_n216), .B2(new_n217), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n221));
  INV_X1    g035(.A(G134), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G137), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT65), .B(G137), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(new_n222), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n221), .B1(new_n225), .B2(new_n207), .ZN(new_n226));
  OAI211_X1 g040(.A(KEYINPUT30), .B(new_n212), .C1(new_n220), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(G134), .B1(new_n200), .B2(new_n201), .ZN(new_n228));
  OAI21_X1  g042(.A(G131), .B1(new_n228), .B2(new_n223), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n229), .A2(new_n217), .A3(new_n216), .A4(new_n221), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n212), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT30), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT2), .B(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n236), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n234), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n227), .A2(new_n233), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n240), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n242), .B(new_n212), .C1(new_n220), .C2(new_n226), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n245));
  INV_X1    g059(.A(G237), .ZN(new_n246));
  INV_X1    g060(.A(G953), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(G210), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n245), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT26), .B(G101), .ZN(new_n250));
  XOR2_X1   g064(.A(new_n249), .B(new_n250), .Z(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT29), .B1(new_n244), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n243), .A2(KEYINPUT70), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT70), .B1(new_n243), .B2(new_n254), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n231), .A2(KEYINPUT69), .A3(new_n240), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n243), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n242), .B1(new_n212), .B2(new_n230), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT69), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT28), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n253), .B1(new_n263), .B2(new_n252), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n216), .A2(new_n217), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n216), .A2(KEYINPUT67), .A3(new_n217), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n226), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n192), .B1(new_n214), .B2(new_n215), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n197), .A2(new_n193), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n199), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n211), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n203), .A2(new_n206), .A3(new_n209), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(new_n242), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n270), .A2(new_n240), .A3(new_n276), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n257), .B1(new_n254), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n251), .A2(KEYINPUT29), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n264), .B(new_n265), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G472), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n241), .A2(new_n243), .A3(new_n251), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT31), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n277), .A2(new_n242), .B1(new_n260), .B2(KEYINPUT69), .ZN(new_n287));
  INV_X1    g101(.A(new_n261), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n254), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n279), .B2(KEYINPUT28), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n243), .A2(KEYINPUT70), .A3(new_n254), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n252), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT71), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n263), .A2(new_n296), .A3(new_n252), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n286), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n298), .A2(KEYINPUT32), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT32), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT31), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n285), .B(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n296), .B1(new_n263), .B2(new_n252), .ZN(new_n305));
  AOI211_X1 g119(.A(KEYINPUT71), .B(new_n251), .C1(new_n257), .C2(new_n262), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n302), .B1(new_n307), .B2(new_n299), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n284), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G217), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(G234), .B2(new_n265), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT22), .B(G137), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n247), .A2(G221), .A3(G234), .ZN(new_n314));
  XOR2_X1   g128(.A(new_n313), .B(new_n314), .Z(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(G140), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(new_n317), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n316), .B2(G140), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n322), .A2(KEYINPUT72), .A3(G125), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n319), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n318), .B1(new_n324), .B2(KEYINPUT16), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT74), .B1(new_n325), .B2(new_n187), .ZN(new_n326));
  INV_X1    g140(.A(new_n318), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n316), .A2(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n320), .A2(new_n316), .A3(G140), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n317), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT16), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(G146), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n319), .A2(new_n328), .A3(new_n187), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n337));
  INV_X1    g151(.A(G119), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(G128), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n340));
  INV_X1    g154(.A(G110), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(G128), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n339), .A2(new_n340), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n343), .A2(KEYINPUT73), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(KEYINPUT73), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n196), .A2(G119), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT24), .B(G110), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n344), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n326), .A2(new_n335), .A3(new_n336), .A4(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n347), .A2(new_n348), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n339), .A2(new_n342), .A3(new_n340), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(G110), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n325), .A2(new_n187), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n187), .B(new_n327), .C1(new_n331), .C2(new_n332), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n355), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n351), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n352), .B1(new_n351), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n315), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n315), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n351), .A2(new_n359), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(KEYINPUT75), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n265), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n367), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n362), .A2(new_n265), .A3(new_n365), .A4(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n312), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n362), .A2(new_n365), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n311), .A2(G902), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G214), .B1(G237), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(G104), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n378), .B2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G104), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(G107), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G101), .ZN(new_n385));
  AND2_X1   g199(.A1(KEYINPUT78), .A2(G101), .ZN(new_n386));
  NOR2_X1   g200(.A1(KEYINPUT78), .A2(G101), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(new_n383), .A3(new_n379), .A4(new_n382), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(KEYINPUT4), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(new_n391), .A3(G101), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n240), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n338), .A3(G116), .ZN(new_n395));
  OAI211_X1 g209(.A(G113), .B(new_n395), .C1(new_n235), .C2(new_n394), .ZN(new_n396));
  INV_X1    g210(.A(new_n383), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n378), .A2(G107), .ZN(new_n398));
  OAI21_X1  g212(.A(G101), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n396), .A2(new_n239), .A3(new_n399), .A4(new_n389), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G122), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n393), .A2(new_n402), .A3(new_n400), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(KEYINPUT6), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n401), .A2(new_n407), .A3(new_n403), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n198), .A2(G125), .A3(new_n199), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n216), .A2(new_n316), .A3(new_n217), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n247), .A2(G224), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n406), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n406), .A2(KEYINPUT80), .A3(new_n408), .A4(new_n413), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n402), .B(KEYINPUT8), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT81), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n400), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n396), .A2(new_n239), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n389), .A2(new_n399), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n421), .A3(new_n424), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n420), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n429));
  OAI211_X1 g243(.A(KEYINPUT7), .B(new_n412), .C1(new_n411), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n412), .A2(new_n429), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n412), .A2(KEYINPUT7), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n409), .A2(new_n410), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n405), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n265), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n418), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G210), .B1(G237), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n418), .A2(new_n438), .A3(new_n436), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(G475), .A2(G902), .ZN(new_n443));
  XOR2_X1   g257(.A(KEYINPUT85), .B(G104), .Z(new_n444));
  XNOR2_X1  g258(.A(G113), .B(G122), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n246), .A2(new_n247), .A3(G214), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(KEYINPUT83), .B2(new_n189), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT83), .B(G143), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n449), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT18), .A3(G131), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n336), .B1(new_n331), .B2(new_n187), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n450), .A2(new_n448), .ZN(new_n454));
  NAND2_X1  g268(.A1(KEYINPUT18), .A2(G131), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n333), .A2(G146), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n451), .A2(KEYINPUT17), .A3(G131), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n458), .A2(new_n357), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT84), .B1(new_n451), .B2(G131), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT17), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n454), .A2(new_n449), .A3(new_n463), .A4(new_n207), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n451), .A2(G131), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n461), .A2(new_n462), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n447), .B(new_n457), .C1(new_n460), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n465), .A3(new_n464), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT19), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n319), .A2(new_n328), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n187), .B(new_n470), .C1(new_n331), .C2(new_n469), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n468), .A2(new_n326), .A3(new_n335), .A4(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n457), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n446), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n443), .B1(new_n467), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n473), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n447), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n466), .A2(new_n357), .A3(new_n458), .A4(new_n459), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n446), .A3(new_n473), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n476), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n475), .B1(new_n481), .B2(KEYINPUT20), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n480), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n483), .A2(new_n476), .A3(new_n484), .A4(new_n443), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n446), .B1(new_n479), .B2(new_n473), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n265), .B1(new_n467), .B2(new_n486), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n482), .A2(new_n485), .B1(G475), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n189), .A2(G128), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n196), .A2(G143), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(new_n222), .ZN(new_n492));
  INV_X1    g306(.A(G116), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G122), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n493), .A2(G122), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n495), .A2(G107), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT14), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n494), .A2(KEYINPUT88), .A3(KEYINPUT14), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n494), .A2(KEYINPUT14), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(new_n496), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n381), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n491), .A2(new_n222), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n495), .A2(new_n496), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(new_n381), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n511), .B2(new_n497), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT13), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n489), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n189), .A2(KEYINPUT13), .A3(G128), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(KEYINPUT87), .A3(new_n515), .A4(new_n490), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n515), .A2(KEYINPUT87), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(G134), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT9), .B(G234), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n521), .A2(new_n310), .A3(G953), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n508), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  OAI22_X1  g337(.A1(new_n499), .A2(new_n507), .B1(new_n512), .B2(new_n519), .ZN(new_n524));
  INV_X1    g338(.A(new_n522), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(G902), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G478), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(KEYINPUT15), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n527), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(G234), .A2(G237), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(G952), .A3(new_n247), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n265), .B1(G234), .B2(G237), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G953), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT21), .B(G898), .Z(new_n535));
  OAI21_X1  g349(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(new_n536), .B(KEYINPUT89), .Z(new_n537));
  AND2_X1   g351(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  AND4_X1   g352(.A1(new_n377), .A2(new_n442), .A3(new_n488), .A4(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G221), .ZN(new_n540));
  INV_X1    g354(.A(new_n521), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n541), .B2(new_n265), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT77), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n392), .A2(new_n198), .A3(new_n199), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n390), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n389), .A2(new_n399), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n546), .B(KEYINPUT10), .C1(new_n218), .C2(new_n219), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n210), .A2(new_n211), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n389), .A2(new_n217), .A3(new_n399), .A4(new_n216), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT10), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n545), .A2(new_n547), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n424), .A2(new_n266), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n549), .ZN(new_n554));
  INV_X1    g368(.A(new_n548), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n554), .A2(KEYINPUT12), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT12), .B1(new_n554), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G110), .B(G140), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n247), .A2(G227), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n544), .A2(new_n390), .B1(new_n550), .B2(new_n549), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n547), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n555), .ZN(new_n565));
  INV_X1    g379(.A(new_n561), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n552), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n562), .A2(new_n567), .A3(G469), .ZN(new_n568));
  NAND2_X1  g382(.A1(G469), .A2(G902), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n552), .B(new_n566), .C1(new_n556), .C2(new_n557), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT79), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n554), .A2(new_n555), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n554), .A2(KEYINPUT12), .A3(new_n555), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n578), .A2(KEYINPUT79), .A3(new_n566), .A4(new_n552), .ZN(new_n579));
  INV_X1    g393(.A(new_n552), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n548), .B1(new_n563), .B2(new_n547), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n561), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n573), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G469), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n265), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n543), .B1(new_n570), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n309), .A2(new_n376), .A3(new_n539), .A4(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n388), .B(KEYINPUT90), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT91), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n587), .B(new_n589), .ZN(G3));
  OAI21_X1  g404(.A(G472), .B1(new_n298), .B2(G902), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n591), .A2(KEYINPUT92), .B1(new_n299), .B2(new_n307), .ZN(new_n592));
  INV_X1    g406(.A(G472), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n307), .B2(new_n265), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n586), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n375), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n592), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT93), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n440), .A2(new_n600), .A3(new_n441), .ZN(new_n601));
  INV_X1    g415(.A(new_n377), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n439), .B(new_n435), .C1(new_n416), .C2(new_n417), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(KEYINPUT93), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n522), .B1(new_n508), .B2(new_n520), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n524), .A2(new_n525), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT33), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n523), .A2(new_n609), .A3(new_n526), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n608), .A2(G478), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n527), .A2(new_n528), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n528), .A2(new_n265), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT94), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT94), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n611), .A2(new_n618), .A3(new_n613), .A4(new_n615), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n485), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT86), .B1(new_n467), .B2(new_n474), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n622), .A2(new_n484), .B1(new_n483), .B2(new_n443), .ZN(new_n623));
  INV_X1    g437(.A(G475), .ZN(new_n624));
  INV_X1    g438(.A(new_n466), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n458), .A2(new_n357), .A3(new_n459), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n473), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n447), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n628), .B2(new_n480), .ZN(new_n629));
  OAI22_X1  g443(.A1(new_n621), .A2(new_n623), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n620), .A2(new_n630), .A3(new_n537), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n599), .A2(new_n605), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n629), .B2(new_n624), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n487), .A2(KEYINPUT95), .A3(G475), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n475), .A2(new_n484), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n483), .A2(KEYINPUT20), .A3(new_n443), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n537), .B(KEYINPUT96), .Z(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n640), .A2(new_n530), .A3(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n643), .A2(new_n601), .A3(new_n604), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n599), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT35), .B(G107), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n364), .A2(KEYINPUT97), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT97), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n351), .A2(new_n359), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n652), .B1(KEYINPUT36), .B2(new_n363), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n363), .A2(KEYINPUT36), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n649), .A2(new_n654), .A3(new_n651), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n653), .A2(new_n373), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n371), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n597), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n592), .A2(new_n539), .A3(new_n596), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  NOR2_X1   g475(.A1(new_n247), .A2(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n533), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(KEYINPUT98), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(KEYINPUT98), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n532), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT99), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n640), .A2(new_n530), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n605), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n309), .A3(new_n658), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XOR2_X1   g486(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n667), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n586), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT102), .Z(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT40), .Z(new_n677));
  INV_X1    g491(.A(new_n657), .ZN(new_n678));
  OAI21_X1  g492(.A(KEYINPUT32), .B1(new_n298), .B2(new_n300), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n307), .A2(new_n302), .A3(new_n299), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(G902), .B1(new_n280), .B2(new_n252), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n244), .A2(new_n251), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n593), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT100), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n687));
  AOI211_X1 g501(.A(new_n687), .B(new_n684), .C1(new_n679), .C2(new_n680), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n442), .B(KEYINPUT38), .ZN(new_n690));
  INV_X1    g504(.A(new_n530), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n690), .A2(new_n377), .A3(new_n630), .A4(new_n691), .ZN(new_n692));
  NOR4_X1   g506(.A1(new_n677), .A2(new_n678), .A3(new_n689), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n189), .ZN(G45));
  INV_X1    g508(.A(new_n605), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n620), .A2(new_n630), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n667), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n309), .A2(new_n695), .A3(new_n658), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NOR2_X1   g513(.A1(new_n605), .A2(new_n631), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n583), .A2(new_n584), .A3(new_n265), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n584), .B1(new_n583), .B2(new_n265), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n701), .A2(new_n702), .A3(new_n542), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n309), .A2(new_n700), .A3(new_n376), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND4_X1  g520(.A1(new_n309), .A2(new_n644), .A3(new_n376), .A4(new_n703), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NAND3_X1  g522(.A1(new_n601), .A2(new_n703), .A3(new_n604), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n488), .B(new_n538), .C1(new_n371), .C2(new_n656), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n309), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT103), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n711), .B1(new_n681), .B2(new_n284), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n710), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  AOI21_X1  g533(.A(new_n438), .B1(new_n418), .B2(new_n436), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n720), .A2(new_n603), .A3(KEYINPUT93), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n630), .A2(new_n691), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n377), .B1(new_n441), .B2(new_n600), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n281), .A2(new_n252), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n300), .B1(new_n725), .B2(new_n304), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n594), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n701), .A2(new_n702), .ZN(new_n728));
  INV_X1    g542(.A(new_n542), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n642), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n724), .A2(new_n727), .A3(new_n376), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  NOR3_X1   g547(.A1(new_n594), .A2(new_n657), .A3(new_n726), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n710), .A3(new_n697), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT104), .B(G125), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G27));
  NAND3_X1  g551(.A1(new_n440), .A2(new_n377), .A3(new_n441), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n569), .B(KEYINPUT105), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n568), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n729), .B1(new_n701), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n309), .A2(new_n376), .A3(new_n697), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n375), .B1(new_n681), .B2(new_n284), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(KEYINPUT42), .A3(new_n697), .A4(new_n742), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  NAND4_X1  g563(.A1(new_n309), .A2(new_n376), .A3(new_n668), .A4(new_n742), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  NAND2_X1  g565(.A1(new_n562), .A2(new_n567), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n562), .A2(new_n567), .A3(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n761));
  INV_X1    g575(.A(new_n756), .ZN(new_n762));
  INV_X1    g576(.A(new_n739), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n759), .A2(new_n585), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n729), .A3(new_n674), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT107), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n592), .A2(new_n596), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n620), .A2(new_n488), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT43), .B1(new_n488), .B2(KEYINPUT108), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n771), .A3(new_n678), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n738), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n773), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n767), .A2(new_n774), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  NAND2_X1  g592(.A1(new_n765), .A2(new_n729), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT47), .Z(new_n780));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n679), .A2(new_n680), .B1(G472), .B2(new_n283), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n782), .A2(new_n375), .A3(new_n697), .A4(new_n775), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n781), .B1(new_n780), .B2(new_n783), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NOR3_X1   g602(.A1(new_n769), .A2(new_n543), .A3(new_n602), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n728), .B(KEYINPUT49), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n790), .A3(new_n376), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n690), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n689), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT112), .B1(new_n671), .B2(new_n735), .ZN(new_n794));
  INV_X1    g608(.A(new_n698), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n605), .A2(new_n667), .A3(new_n722), .A4(new_n741), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n797), .B(new_n657), .C1(new_n686), .C2(new_n688), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n671), .A2(new_n735), .A3(KEYINPUT112), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(KEYINPUT52), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n698), .A2(new_n671), .A3(new_n735), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n798), .ZN(new_n802));
  XOR2_X1   g616(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT53), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n734), .A2(new_n697), .A3(new_n742), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n691), .A2(new_n667), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n738), .A2(new_n808), .A3(new_n640), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n309), .A2(new_n658), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n750), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT110), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n750), .A2(new_n810), .A3(new_n807), .A4(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n812), .A2(new_n748), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n716), .B1(new_n715), .B2(new_n710), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n782), .A2(new_n709), .A3(KEYINPUT103), .A4(new_n711), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n377), .B(new_n641), .C1(new_n720), .C2(new_n603), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n488), .A2(new_n691), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n819), .B1(new_n696), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n592), .A2(new_n821), .A3(new_n596), .A4(new_n598), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n704), .A2(new_n707), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n587), .A2(new_n659), .A3(new_n732), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n818), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT111), .B1(new_n815), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n812), .A2(new_n748), .A3(new_n814), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n704), .A2(new_n707), .A3(new_n822), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n587), .A2(new_n659), .A3(new_n732), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n718), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n827), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n806), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n801), .A2(KEYINPUT52), .A3(new_n798), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(new_n801), .B2(new_n798), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n750), .A2(new_n807), .A3(new_n810), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n838), .A2(new_n813), .B1(new_n745), .B2(new_n747), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n825), .A2(new_n839), .A3(KEYINPUT111), .A4(new_n812), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n831), .B1(new_n827), .B2(new_n830), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n833), .B(KEYINPUT54), .C1(new_n834), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n827), .A2(new_n830), .A3(new_n834), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n800), .A2(new_n805), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g661(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n848));
  OAI211_X1 g662(.A(new_n847), .B(new_n848), .C1(new_n842), .C2(KEYINPUT53), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n843), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n532), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n771), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n852), .A2(new_n376), .A3(new_n727), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n690), .A2(new_n377), .A3(new_n730), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT50), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n730), .A2(new_n738), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n852), .A2(new_n734), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n689), .A2(new_n376), .A3(new_n851), .A4(new_n857), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n859), .A2(new_n630), .A3(new_n620), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n728), .A2(new_n543), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n780), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n853), .A2(new_n775), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT51), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n852), .A2(new_n746), .A3(new_n857), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT48), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n247), .A2(G952), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n853), .B2(new_n710), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n868), .B(new_n870), .C1(new_n696), .C2(new_n859), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n843), .A2(new_n849), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT115), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n863), .A2(KEYINPUT116), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n863), .A2(KEYINPUT116), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n864), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n861), .A2(KEYINPUT51), .A3(new_n877), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n850), .A2(new_n872), .A3(new_n874), .A4(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(G952), .A2(G953), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n793), .B1(new_n879), .B2(new_n880), .ZN(G75));
  AND2_X1   g695(.A1(new_n845), .A2(new_n846), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n826), .A2(new_n832), .B1(new_n836), .B2(new_n835), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n882), .B1(new_n883), .B2(new_n834), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n265), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(G210), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n406), .A2(new_n408), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(new_n413), .Z(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT55), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n886), .A2(new_n887), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n886), .B2(new_n887), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n247), .A2(G952), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(G51));
  NAND2_X1  g708(.A1(new_n883), .A2(new_n834), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n896), .A3(new_n848), .A4(new_n847), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n849), .A2(KEYINPUT117), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n847), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n901));
  INV_X1    g715(.A(new_n848), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT118), .B1(new_n884), .B2(new_n848), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n739), .B(KEYINPUT57), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n583), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n885), .A2(new_n762), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n893), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND3_X1  g724(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n480), .A3(new_n478), .ZN(new_n912));
  INV_X1    g726(.A(new_n893), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .A4(new_n483), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G60));
  XNOR2_X1  g729(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n615), .B(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n874), .B2(new_n850), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n608), .A2(new_n610), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n913), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n917), .B1(new_n608), .B2(new_n610), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n905), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT120), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n905), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n920), .B1(new_n923), .B2(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT121), .Z(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT60), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n884), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n655), .A3(new_n653), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n931), .B(new_n913), .C1(new_n372), .C2(new_n930), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G66));
  AOI21_X1  g748(.A(new_n247), .B1(new_n535), .B2(G224), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n830), .B2(new_n247), .ZN(new_n936));
  INV_X1    g750(.A(G898), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n888), .B1(new_n937), .B2(G953), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n936), .B(new_n938), .ZN(G69));
  NAND2_X1  g753(.A1(G227), .A2(G900), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(G953), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n227), .A2(new_n233), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT122), .Z(new_n943));
  OAI21_X1  g757(.A(new_n470), .B1(new_n331), .B2(new_n469), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n796), .A2(new_n799), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n693), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT62), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n738), .B1(new_n696), .B2(new_n820), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n676), .A2(new_n746), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n777), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT123), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n948), .A2(new_n787), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n945), .B1(new_n954), .B2(G953), .ZN(new_n955));
  INV_X1    g769(.A(new_n946), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n777), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n748), .B(new_n750), .C1(new_n785), .C2(new_n786), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n767), .A2(new_n746), .A3(new_n724), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n959), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n662), .B1(new_n969), .B2(new_n247), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n941), .B(new_n955), .C1(new_n970), .C2(new_n945), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n959), .A2(new_n964), .A3(new_n967), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n967), .B1(new_n959), .B2(new_n964), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n247), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n662), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(G953), .B(new_n940), .C1(new_n976), .C2(new_n945), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n971), .A2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n969), .B2(new_n830), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n244), .A2(new_n251), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n980), .B1(new_n953), .B2(new_n830), .ZN(new_n984));
  INV_X1    g798(.A(new_n683), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n893), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n833), .B1(new_n842), .B2(new_n834), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n683), .A2(new_n980), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n987), .A2(new_n982), .A3(new_n988), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT127), .Z(new_n990));
  AND3_X1   g804(.A1(new_n983), .A2(new_n986), .A3(new_n990), .ZN(G57));
endmodule


