//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G134), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT65), .B1(new_n191), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(new_n189), .A3(G134), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(KEYINPUT66), .A3(G137), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n190), .A2(new_n192), .A3(new_n194), .A4(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n199), .B(new_n201), .C1(KEYINPUT1), .C2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n200), .A2(G146), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n198), .A2(G143), .ZN(new_n206));
  OAI211_X1 g020(.A(G128), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT11), .B1(new_n191), .B2(G137), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n189), .A3(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT64), .A2(G131), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT64), .A2(G131), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n191), .A2(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n197), .A2(new_n203), .A3(new_n207), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT69), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n208), .A2(new_n210), .B1(new_n191), .B2(G137), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n214), .A2(new_n219), .B1(new_n196), .B2(G131), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n207), .A2(new_n203), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n225));
  INV_X1    g039(.A(G116), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT68), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G116), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n229), .A3(G119), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G116), .ZN(new_n232));
  INV_X1    g046(.A(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT2), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT2), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n230), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n230), .B2(new_n232), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n225), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n199), .A2(new_n201), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G143), .B(G146), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G128), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n211), .B2(new_n215), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n230), .A2(new_n232), .ZN(new_n252));
  INV_X1    g066(.A(new_n237), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n238), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n241), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n224), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n217), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT30), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT67), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n262), .A3(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n218), .A2(new_n223), .A3(KEYINPUT30), .A4(new_n251), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n254), .A2(new_n238), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n257), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n269));
  XOR2_X1   g083(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n270));
  NOR2_X1   g084(.A1(G237), .A2(G953), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G210), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n270), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT26), .B(G101), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n273), .B(new_n274), .Z(new_n275));
  NAND4_X1  g089(.A1(new_n268), .A2(KEYINPUT72), .A3(new_n269), .A4(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n262), .B1(new_n258), .B2(new_n259), .ZN(new_n277));
  AOI211_X1 g091(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n251), .C2(new_n217), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n266), .B(new_n265), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n217), .A2(KEYINPUT69), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n221), .B1(new_n220), .B2(new_n222), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n256), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n279), .A2(new_n269), .A3(new_n284), .A4(new_n275), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n276), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n279), .A2(new_n284), .A3(new_n275), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT31), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n258), .A2(new_n266), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n224), .B2(new_n256), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT28), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n241), .A2(new_n255), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(new_n258), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n294), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n290), .B1(new_n300), .B2(new_n275), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n187), .B1(new_n288), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT32), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n187), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(new_n303), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n288), .B2(new_n301), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT76), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n268), .B2(new_n275), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n298), .A2(new_n275), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n294), .A2(new_n295), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n309), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n218), .A2(new_n223), .A3(new_n251), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n282), .A2(new_n283), .B1(new_n315), .B2(new_n297), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT75), .B1(new_n316), .B2(new_n296), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n315), .A2(new_n297), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n318), .B(KEYINPUT28), .C1(new_n319), .C2(new_n257), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n312), .A2(new_n310), .ZN(new_n322));
  AOI21_X1  g136(.A(G902), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n292), .A2(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT28), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n275), .A3(new_n326), .A4(new_n298), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n279), .A2(new_n284), .ZN(new_n328));
  INV_X1    g142(.A(new_n275), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n327), .A2(new_n330), .A3(KEYINPUT74), .A4(new_n310), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n314), .A2(new_n323), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G472), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n325), .A2(new_n326), .A3(new_n298), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n334), .A2(new_n329), .B1(KEYINPUT31), .B2(new_n289), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n276), .A2(new_n287), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n306), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n304), .A2(new_n308), .A3(new_n333), .A4(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT9), .B(G234), .ZN(new_n341));
  OAI21_X1  g155(.A(G221), .B1(new_n341), .B2(G902), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT84), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G110), .B(G140), .ZN(new_n345));
  INV_X1    g159(.A(G227), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G953), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G104), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT86), .B1(new_n350), .B2(G107), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n352));
  INV_X1    g166(.A(G107), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(G104), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(G107), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G101), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(new_n350), .B2(G107), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n353), .A3(G104), .ZN(new_n360));
  INV_X1    g174(.A(G101), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n358), .A2(new_n360), .A3(new_n361), .A4(new_n355), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n207), .A2(new_n203), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT10), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n222), .A2(new_n366), .A3(new_n362), .A4(new_n357), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n248), .A2(new_n250), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n358), .A2(new_n360), .A3(new_n355), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G101), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT85), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n370), .A2(KEYINPUT85), .A3(new_n371), .A4(G101), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n371), .B1(new_n370), .B2(G101), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n246), .B1(new_n377), .B2(new_n362), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n368), .A2(new_n369), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT87), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n365), .A2(new_n367), .B1(new_n376), .B2(new_n378), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n369), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n382), .A2(new_n369), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n349), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n357), .A2(new_n362), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(new_n222), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n363), .A2(new_n364), .ZN(new_n390));
  OAI22_X1  g204(.A1(new_n389), .A2(new_n390), .B1(new_n248), .B2(new_n250), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT12), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n348), .B1(new_n381), .B2(new_n384), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n393), .B2(KEYINPUT88), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n380), .A2(KEYINPUT87), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n383), .B1(new_n382), .B2(new_n369), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n349), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT88), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n387), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n400), .A2(G469), .A3(G902), .ZN(new_n401));
  INV_X1    g215(.A(G469), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT12), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n391), .B(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n385), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n348), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n393), .A2(new_n386), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G902), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n402), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n344), .B1(new_n401), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G214), .B1(G237), .B2(G902), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G210), .B1(G237), .B2(G902), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n230), .A2(KEYINPUT5), .A3(new_n232), .ZN(new_n416));
  OAI21_X1  g230(.A(G113), .B1(new_n232), .B2(KEYINPUT5), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n388), .A2(new_n238), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n376), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n377), .A2(new_n362), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n266), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n420), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G122), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n425), .B(new_n420), .C1(new_n421), .C2(new_n423), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n424), .A2(new_n430), .A3(new_n426), .ZN(new_n431));
  AOI21_X1  g245(.A(G125), .B1(new_n207), .B2(new_n203), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n432), .A2(new_n433), .B1(G125), .B2(new_n246), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT89), .B1(new_n222), .B2(G125), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G224), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(G953), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n436), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n429), .A2(new_n431), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n409), .ZN(new_n441));
  INV_X1    g255(.A(new_n438), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT7), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G125), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n364), .A2(new_n433), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n246), .A2(G125), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n432), .A2(new_n433), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n434), .A2(new_n435), .A3(new_n444), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n443), .B1(new_n442), .B2(KEYINPUT7), .ZN(new_n454));
  INV_X1    g268(.A(new_n232), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT68), .B(G116), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n456), .B2(G119), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n416), .A2(new_n418), .B1(new_n457), .B2(new_n237), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n417), .A2(KEYINPUT90), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT90), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(G113), .C1(new_n232), .C2(KEYINPUT5), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n416), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n357), .A2(new_n238), .A3(new_n362), .ZN(new_n463));
  OAI22_X1  g277(.A1(new_n458), .A2(new_n388), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n425), .B(KEYINPUT8), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n454), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n453), .A2(new_n466), .A3(KEYINPUT92), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n428), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT92), .B1(new_n453), .B2(new_n466), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n415), .B1(new_n441), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n469), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n428), .A3(new_n467), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n473), .A2(new_n409), .A3(new_n414), .A4(new_n440), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n413), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  INV_X1    g291(.A(G217), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n341), .A2(new_n478), .A3(G953), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n227), .A2(new_n229), .A3(G122), .ZN(new_n481));
  OR2_X1    g295(.A1(new_n226), .A2(G122), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT98), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT98), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n485), .A3(new_n482), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n353), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT99), .B1(new_n202), .B2(G143), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT99), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n200), .A3(G128), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n200), .A2(G128), .ZN(new_n492));
  OAI21_X1  g306(.A(G134), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(new_n490), .ZN(new_n494));
  INV_X1    g308(.A(new_n492), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n191), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT14), .A4(G122), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n497), .A2(G107), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n481), .A2(new_n499), .A3(new_n482), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n493), .A2(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n496), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n481), .A2(new_n485), .A3(new_n482), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n485), .B1(new_n481), .B2(new_n482), .ZN(new_n504));
  OAI21_X1  g318(.A(G107), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n505), .B2(new_n487), .ZN(new_n506));
  OAI211_X1 g320(.A(KEYINPUT100), .B(new_n495), .C1(new_n491), .C2(KEYINPUT13), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT100), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT13), .B1(new_n488), .B2(new_n490), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n508), .B1(new_n509), .B2(new_n492), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n491), .A2(KEYINPUT13), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G134), .ZN(new_n513));
  AOI221_X4 g327(.A(new_n480), .B1(new_n487), .B2(new_n501), .C1(new_n506), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n506), .A2(new_n513), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n501), .A2(new_n487), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n479), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n409), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT101), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT101), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n520), .B(new_n409), .C1(new_n514), .C2(new_n517), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n477), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n477), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G953), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n409), .B(new_n525), .C1(G234), .C2(G237), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT21), .B(G898), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(KEYINPUT102), .A2(G952), .ZN(new_n529));
  NAND2_X1  g343(.A1(KEYINPUT102), .A2(G952), .ZN(new_n530));
  AOI21_X1  g344(.A(G953), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G234), .ZN(new_n532));
  INV_X1    g346(.A(G237), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n522), .A2(new_n524), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT96), .B(G104), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n271), .A2(G214), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n200), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n271), .A2(G143), .A3(G214), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n214), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT94), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n542), .A2(new_n548), .A3(new_n214), .A4(new_n543), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G140), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G125), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n446), .A2(G140), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT19), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT19), .B1(new_n552), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n198), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n556), .A2(KEYINPUT95), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT79), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n552), .A2(new_n553), .A3(new_n558), .A4(KEYINPUT16), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT16), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT79), .B1(new_n552), .B2(KEYINPUT16), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G146), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n556), .A2(KEYINPUT95), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n550), .A2(new_n557), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT93), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n552), .A2(new_n553), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G146), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n567), .A2(G146), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n552), .A2(new_n553), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n198), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT93), .A3(new_n568), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n544), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT18), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(new_n249), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n544), .A2(KEYINPUT18), .A3(G131), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n540), .B1(new_n565), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n198), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT80), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT16), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n586), .B(KEYINPUT79), .C1(KEYINPUT16), .C2(new_n552), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n198), .B1(new_n587), .B2(new_n559), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n563), .A2(new_n584), .A3(new_n583), .ZN(new_n590));
  INV_X1    g404(.A(new_n547), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n589), .A2(new_n590), .B1(KEYINPUT17), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n546), .A2(new_n593), .A3(new_n547), .A4(new_n549), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n582), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n581), .B1(new_n595), .B2(new_n540), .ZN(new_n596));
  NOR2_X1   g410(.A1(G475), .A2(G902), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(KEYINPUT97), .B(new_n537), .C1(new_n596), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n591), .A2(KEYINPUT17), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n585), .A2(new_n588), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n562), .A2(KEYINPUT80), .A3(G146), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n594), .B(new_n600), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n603), .A2(new_n580), .A3(new_n540), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n540), .B1(new_n603), .B2(new_n580), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n409), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G475), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n603), .A2(new_n580), .A3(new_n540), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n565), .A2(new_n580), .ZN(new_n609));
  INV_X1    g423(.A(new_n540), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n598), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT20), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI211_X1 g428(.A(KEYINPUT97), .B(new_n598), .C1(new_n608), .C2(new_n611), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n599), .B(new_n607), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n475), .A2(new_n536), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n411), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n478), .B1(G234), .B2(new_n409), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT25), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n231), .A2(G128), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n231), .A2(G128), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(KEYINPUT23), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G110), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT78), .ZN(new_n628));
  OR3_X1    g442(.A1(new_n231), .A2(KEYINPUT77), .A3(G128), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT77), .B1(new_n231), .B2(G128), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n630), .A3(new_n623), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT24), .B(G110), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n589), .A2(new_n590), .A3(new_n628), .A4(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n631), .A2(KEYINPUT81), .A3(new_n632), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(G110), .B2(new_n626), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT81), .B1(new_n631), .B2(new_n632), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n563), .B(new_n573), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT22), .B(G137), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n525), .A2(G221), .A3(G234), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT82), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n634), .A2(new_n638), .A3(new_n642), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n622), .B1(new_n646), .B2(G902), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n644), .A2(KEYINPUT25), .A3(new_n409), .A4(new_n645), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n621), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n646), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n621), .A2(new_n409), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT83), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n340), .A2(new_n619), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G101), .ZN(G3));
  INV_X1    g470(.A(G472), .ZN(new_n657));
  AOI21_X1  g471(.A(G902), .B1(new_n335), .B2(new_n336), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n302), .B(new_n654), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n411), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n515), .A2(new_n516), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n480), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n506), .A2(new_n513), .B1(new_n487), .B2(new_n501), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n479), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT33), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n476), .A2(G902), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n517), .A2(KEYINPUT103), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n663), .B2(new_n479), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n668), .A2(new_n670), .A3(KEYINPUT33), .A4(new_n664), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n664), .A2(KEYINPUT33), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n674), .A2(KEYINPUT104), .A3(new_n668), .A4(new_n670), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n665), .B(new_n667), .C1(new_n673), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n662), .A2(new_n664), .ZN(new_n677));
  AOI21_X1  g491(.A(G478), .B1(new_n677), .B2(new_n409), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n616), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n535), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n475), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n660), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT34), .B(G104), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G6));
  INV_X1    g499(.A(new_n477), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n520), .B1(new_n677), .B2(new_n409), .ZN(new_n687));
  INV_X1    g501(.A(new_n521), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n523), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n617), .A2(new_n475), .A3(new_n680), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n660), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT35), .B(G107), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G9));
  AOI21_X1  g508(.A(new_n657), .B1(new_n337), .B2(new_n409), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n305), .B1(new_n335), .B2(new_n336), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n643), .A2(KEYINPUT36), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n639), .B(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n698), .A2(new_n652), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n649), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n695), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n619), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT37), .B(G110), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT105), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n702), .B(new_n704), .ZN(G12));
  NOR2_X1   g519(.A1(new_n522), .A2(new_n524), .ZN(new_n706));
  INV_X1    g520(.A(new_n534), .ZN(new_n707));
  INV_X1    g521(.A(G900), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n707), .B1(new_n708), .B2(new_n526), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n706), .A2(new_n616), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n385), .A2(new_n386), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n348), .ZN(new_n712));
  OAI211_X1 g526(.A(KEYINPUT88), .B(new_n349), .C1(new_n395), .C2(new_n396), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n404), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n393), .A2(KEYINPUT88), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n402), .A3(new_n409), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n402), .A2(new_n409), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n405), .A2(new_n348), .B1(new_n386), .B2(new_n393), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n718), .B1(new_n719), .B2(G469), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n343), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n710), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n649), .A2(new_n699), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n340), .A2(new_n722), .A3(new_n475), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  AND2_X1   g539(.A1(new_n471), .A2(new_n474), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT38), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n617), .A2(new_n706), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n412), .A3(new_n700), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n316), .A2(new_n275), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n268), .B2(new_n275), .ZN(new_n732));
  OAI21_X1  g546(.A(G472), .B1(new_n732), .B2(G902), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n304), .A2(new_n308), .A3(new_n339), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g551(.A(new_n709), .B(KEYINPUT39), .Z(new_n738));
  NAND2_X1  g552(.A1(new_n721), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(KEYINPUT40), .Z(new_n740));
  NAND3_X1  g554(.A1(new_n730), .A2(KEYINPUT106), .A3(new_n734), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G143), .ZN(G45));
  INV_X1    g557(.A(new_n709), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n616), .B(new_n744), .C1(new_n676), .C2(new_n678), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n411), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n340), .A3(new_n475), .A4(new_n723), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G146), .ZN(G48));
  NAND2_X1  g562(.A1(new_n717), .A2(new_n344), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n716), .A2(new_n409), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n402), .B1(new_n750), .B2(KEYINPUT107), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n716), .A2(new_n752), .A3(new_n409), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n749), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n340), .A2(new_n682), .A3(new_n654), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT41), .B(G113), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G15));
  NAND4_X1  g571(.A1(new_n340), .A2(new_n654), .A3(new_n691), .A4(new_n754), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G116), .ZN(G18));
  OAI21_X1  g573(.A(KEYINPUT107), .B1(new_n400), .B2(G902), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(G469), .A3(new_n753), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n689), .A2(new_n680), .A3(new_n523), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n616), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n394), .A2(new_n399), .ZN(new_n764));
  AOI21_X1  g578(.A(G902), .B1(new_n764), .B2(new_n712), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n343), .B1(new_n765), .B2(new_n402), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n761), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(new_n340), .A3(new_n475), .A4(new_n723), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G119), .ZN(G21));
  XOR2_X1   g583(.A(new_n187), .B(KEYINPUT108), .Z(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n276), .A2(new_n287), .B1(KEYINPUT31), .B2(new_n289), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n321), .A2(new_n298), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n329), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n771), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n649), .A2(new_n653), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n695), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n475), .A2(new_n616), .A3(new_n680), .A4(new_n690), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n754), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT109), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n285), .A2(new_n286), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n285), .A2(new_n286), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n290), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n275), .B1(new_n321), .B2(new_n298), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n770), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(new_n654), .C1(new_n657), .C2(new_n658), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n778), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n754), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n781), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G122), .ZN(G24));
  NOR3_X1   g606(.A1(new_n695), .A2(new_n775), .A3(new_n700), .ZN(new_n793));
  INV_X1    g607(.A(new_n745), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n754), .A3(new_n794), .A4(new_n475), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G125), .ZN(G27));
  NAND2_X1  g610(.A1(new_n340), .A2(new_n654), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n745), .A2(KEYINPUT42), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n471), .A2(new_n412), .A3(new_n474), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n721), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n745), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n304), .A2(new_n333), .A3(new_n307), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n803), .A2(KEYINPUT110), .A3(new_n654), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT110), .B1(new_n803), .B2(new_n654), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n801), .B1(new_n806), .B2(KEYINPUT42), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G131), .ZN(G33));
  INV_X1    g622(.A(new_n800), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n340), .A3(new_n654), .A4(new_n710), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G134), .ZN(G36));
  INV_X1    g625(.A(KEYINPUT45), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n402), .B1(new_n408), .B2(new_n812), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n813), .A2(KEYINPUT111), .B1(KEYINPUT45), .B2(new_n719), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n408), .A2(new_n812), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(G469), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n718), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n717), .B1(new_n819), .B2(KEYINPUT46), .ZN(new_n820));
  INV_X1    g634(.A(new_n718), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n815), .A2(KEYINPUT111), .A3(G469), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n719), .A2(KEYINPUT45), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n813), .A2(KEYINPUT111), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT46), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n344), .B(new_n738), .C1(new_n820), .C2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n799), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT44), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT43), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n665), .B1(new_n673), .B2(new_n675), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n678), .B1(new_n834), .B2(new_n666), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n616), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  OAI211_X1 g653(.A(KEYINPUT112), .B(KEYINPUT43), .C1(new_n835), .C2(new_n616), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n695), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n700), .B1(new_n842), .B2(new_n302), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n839), .B1(new_n838), .B2(new_n840), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n832), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n845), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(KEYINPUT44), .A3(new_n841), .A4(new_n843), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n831), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G137), .ZN(G39));
  NOR4_X1   g664(.A1(new_n340), .A2(new_n654), .A3(new_n745), .A4(new_n830), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n826), .A2(new_n827), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n814), .A2(new_n818), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(KEYINPUT46), .A3(new_n821), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n852), .A2(new_n717), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(KEYINPUT47), .A3(new_n344), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT47), .B1(new_n855), .B2(new_n344), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n851), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(G140), .ZN(G42));
  NAND4_X1  g674(.A1(new_n838), .A2(new_n707), .A3(new_n777), .A4(new_n840), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n754), .A2(new_n475), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n863), .A2(new_n531), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n754), .A2(new_n707), .A3(new_n799), .ZN(new_n865));
  INV_X1    g679(.A(new_n734), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n654), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n840), .A3(new_n838), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n804), .A2(new_n805), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT48), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n871), .B1(new_n869), .B2(new_n870), .ZN(new_n873));
  OAI221_X1 g687(.A(new_n864), .B1(new_n679), .B2(new_n867), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n855), .A2(new_n344), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT47), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n761), .A2(new_n717), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n877), .B(new_n856), .C1(new_n344), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n861), .A2(new_n830), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT118), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n793), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n835), .A2(new_n617), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n883), .A2(new_n868), .B1(new_n867), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT50), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n727), .A2(new_n413), .A3(new_n754), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n861), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n886), .B1(new_n861), .B2(new_n887), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT51), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n882), .A2(new_n893), .A3(new_n890), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n874), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n655), .A2(new_n683), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT114), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT114), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n655), .A2(new_n683), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT115), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n689), .A2(new_n901), .A3(new_n523), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT115), .B1(new_n522), .B2(new_n524), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n616), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n535), .B(new_n413), .C1(new_n471), .C2(new_n474), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n660), .A2(new_n906), .B1(new_n619), .B2(new_n701), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(new_n768), .A3(new_n755), .A4(new_n758), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n900), .A2(new_n909), .A3(new_n791), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n616), .A2(new_n709), .ZN(new_n911));
  AND4_X1   g725(.A1(new_n799), .A2(new_n911), .A3(new_n903), .A4(new_n902), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n340), .A2(new_n721), .A3(new_n912), .A4(new_n723), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n809), .A2(new_n793), .A3(new_n794), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n810), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n807), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n724), .A2(new_n795), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT116), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n700), .A2(new_n744), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT117), .B1(new_n411), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n728), .A2(new_n475), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT117), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n721), .A2(new_n923), .A3(new_n700), .A4(new_n744), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n921), .A2(new_n734), .A3(new_n922), .A4(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(KEYINPUT52), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT116), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n724), .A2(new_n927), .A3(new_n795), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n919), .A2(new_n926), .A3(new_n747), .A4(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n747), .A2(new_n925), .A3(new_n724), .A4(new_n795), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT52), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT53), .B1(new_n917), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n789), .B1(new_n788), .B2(new_n754), .ZN(new_n935));
  AND4_X1   g749(.A1(new_n789), .A2(new_n777), .A3(new_n754), .A4(new_n779), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n908), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n938), .A2(new_n807), .A3(new_n900), .A4(new_n915), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n930), .B(KEYINPUT52), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT53), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT54), .B1(new_n934), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n939), .B2(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n660), .A2(new_n906), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n755), .A2(new_n702), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n768), .A2(new_n758), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n947), .A3(new_n791), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n655), .A2(new_n683), .A3(new_n898), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n898), .B1(new_n655), .B2(new_n683), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n806), .A2(KEYINPUT42), .ZN(new_n953));
  INV_X1    g767(.A(new_n801), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n915), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n933), .A2(new_n952), .A3(KEYINPUT53), .A4(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT54), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n944), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n895), .A2(new_n943), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(G952), .A2(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n776), .A2(new_n343), .A3(new_n413), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n866), .A2(new_n727), .A3(new_n836), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n878), .A2(KEYINPUT49), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n878), .A2(KEYINPUT49), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n961), .A2(new_n966), .ZN(G75));
  NOR2_X1   g781(.A1(new_n525), .A2(G952), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n409), .B1(new_n944), .B2(new_n956), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT56), .B1(new_n970), .B2(G210), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n429), .A2(new_n431), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(new_n439), .Z(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT55), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n969), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  AOI211_X1 g790(.A(KEYINPUT56), .B(new_n974), .C1(new_n970), .C2(G210), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G51));
  XNOR2_X1  g792(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n718), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n944), .A2(new_n956), .A3(new_n957), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n957), .B1(new_n944), .B2(new_n956), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n716), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n853), .B(KEYINPUT120), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n970), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n968), .B1(new_n984), .B2(new_n986), .ZN(G54));
  INV_X1    g801(.A(new_n596), .ZN(new_n988));
  AND2_X1   g802(.A1(KEYINPUT58), .A2(G475), .ZN(new_n989));
  AOI211_X1 g803(.A(KEYINPUT121), .B(new_n988), .C1(new_n970), .C2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT121), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n944), .A2(new_n956), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(G902), .A3(new_n989), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n991), .B1(new_n993), .B2(new_n596), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n992), .A2(G902), .A3(new_n988), .A4(new_n989), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n969), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n990), .A2(new_n994), .A3(new_n996), .ZN(G60));
  NAND2_X1  g811(.A1(new_n943), .A2(new_n958), .ZN(new_n998));
  NAND2_X1  g812(.A1(G478), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT59), .Z(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n834), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n834), .A2(new_n1001), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n981), .B2(new_n982), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n969), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1002), .A2(new_n1005), .ZN(G63));
  NAND2_X1  g820(.A1(G217), .A2(G902), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT60), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n992), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT122), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1010), .A2(new_n1011), .A3(new_n646), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1008), .B1(new_n944), .B2(new_n956), .ZN(new_n1013));
  OAI21_X1  g827(.A(KEYINPUT122), .B1(new_n1013), .B2(new_n650), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n968), .B1(new_n1013), .B2(new_n698), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(KEYINPUT61), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT61), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n992), .A2(new_n698), .A3(new_n1009), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n969), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1013), .A2(new_n650), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1016), .A2(new_n1021), .ZN(G66));
  OAI21_X1  g836(.A(G953), .B1(new_n527), .B2(new_n437), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1023), .B1(new_n952), .B2(G953), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n972), .B1(G898), .B2(new_n525), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(G69));
  OAI21_X1  g840(.A(G953), .B1(new_n346), .B2(new_n708), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT125), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n264), .A2(new_n265), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT123), .Z(new_n1030));
  OR2_X1    g844(.A1(new_n554), .A2(new_n555), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1030), .B(new_n1031), .Z(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT62), .ZN(new_n1034));
  INV_X1    g848(.A(new_n747), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1035), .B1(new_n918), .B2(KEYINPUT116), .ZN(new_n1036));
  AND2_X1   g850(.A1(new_n1036), .A2(new_n928), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1034), .B1(new_n1037), .B2(new_n742), .ZN(new_n1038));
  INV_X1    g852(.A(new_n835), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n904), .B1(new_n616), .B2(new_n1039), .ZN(new_n1040));
  OR4_X1    g854(.A1(new_n797), .A2(new_n1040), .A3(new_n739), .A4(new_n830), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n859), .A2(new_n849), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g857(.A1(new_n742), .A2(new_n1036), .A3(new_n1034), .A4(new_n928), .ZN(new_n1044));
  XNOR2_X1  g858(.A(new_n1044), .B(KEYINPUT124), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1033), .B1(new_n1046), .B2(new_n525), .ZN(new_n1047));
  AND2_X1   g861(.A1(new_n859), .A2(new_n849), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n807), .A2(new_n810), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1036), .A2(new_n928), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n922), .B1(new_n804), .B2(new_n805), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n829), .A2(new_n1051), .ZN(new_n1052));
  NOR3_X1   g866(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1054), .A2(new_n525), .ZN(new_n1055));
  NOR2_X1   g869(.A1(new_n525), .A2(G900), .ZN(new_n1056));
  INV_X1    g870(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n1032), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1028), .B1(new_n1047), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g873(.A(G953), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1060));
  OAI21_X1  g874(.A(new_n1033), .B1(new_n1060), .B2(new_n1056), .ZN(new_n1061));
  INV_X1    g875(.A(new_n1028), .ZN(new_n1062));
  AOI21_X1  g876(.A(G953), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1063));
  OAI211_X1 g877(.A(new_n1061), .B(new_n1062), .C1(new_n1063), .C2(new_n1033), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1059), .A2(new_n1064), .ZN(G72));
  XOR2_X1   g879(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1066));
  NOR2_X1   g880(.A1(new_n657), .A2(new_n409), .ZN(new_n1067));
  XNOR2_X1  g881(.A(new_n1066), .B(new_n1067), .ZN(new_n1068));
  OAI21_X1  g882(.A(new_n1068), .B1(new_n1054), .B2(new_n910), .ZN(new_n1069));
  XNOR2_X1  g883(.A(new_n328), .B(KEYINPUT127), .ZN(new_n1070));
  NOR2_X1   g884(.A1(new_n1070), .A2(new_n275), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g886(.A1(new_n330), .A2(new_n289), .ZN(new_n1073));
  OAI211_X1 g887(.A(new_n1068), .B(new_n1073), .C1(new_n934), .C2(new_n942), .ZN(new_n1074));
  NAND3_X1  g888(.A1(new_n1072), .A2(new_n969), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n1070), .A2(new_n275), .ZN(new_n1076));
  NAND3_X1  g890(.A1(new_n1043), .A2(new_n1045), .A3(new_n952), .ZN(new_n1077));
  AOI21_X1  g891(.A(new_n1076), .B1(new_n1077), .B2(new_n1068), .ZN(new_n1078));
  NOR2_X1   g892(.A1(new_n1075), .A2(new_n1078), .ZN(G57));
endmodule


