

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582;

  XNOR2_X1 U324 ( .A(n425), .B(n424), .ZN(n426) );
  NOR2_X1 U325 ( .A1(n518), .A2(n445), .ZN(n567) );
  XNOR2_X1 U326 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n446) );
  XNOR2_X1 U327 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U328 ( .A(n573), .B(KEYINPUT41), .Z(n551) );
  XNOR2_X1 U329 ( .A(KEYINPUT31), .B(KEYINPUT74), .ZN(n292) );
  XNOR2_X1 U330 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n424) );
  INV_X1 U331 ( .A(KEYINPUT48), .ZN(n428) );
  XNOR2_X1 U332 ( .A(n428), .B(KEYINPUT64), .ZN(n429) );
  INV_X1 U333 ( .A(KEYINPUT65), .ZN(n359) );
  XNOR2_X1 U334 ( .A(n430), .B(n429), .ZN(n529) );
  XNOR2_X1 U335 ( .A(n391), .B(n292), .ZN(n392) );
  XNOR2_X1 U336 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U337 ( .A(n393), .B(n392), .ZN(n399) );
  XNOR2_X1 U338 ( .A(n447), .B(n446), .ZN(n448) );
  NOR2_X1 U339 ( .A1(n534), .A2(n448), .ZN(n564) );
  XNOR2_X1 U340 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U341 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n294) );
  XNOR2_X1 U343 ( .A(KEYINPUT17), .B(KEYINPUT88), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U345 ( .A(KEYINPUT19), .B(n295), .Z(n434) );
  XOR2_X1 U346 ( .A(KEYINPUT66), .B(G99GAT), .Z(n297) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U349 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n299) );
  XNOR2_X1 U350 ( .A(G183GAT), .B(G176GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U352 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U353 ( .A(G71GAT), .B(G15GAT), .Z(n303) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(n304), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n434), .B(n307), .ZN(n312) );
  XOR2_X1 U359 ( .A(KEYINPUT0), .B(G120GAT), .Z(n309) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(G127GAT), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n311) );
  XOR2_X1 U362 ( .A(G134GAT), .B(KEYINPUT85), .Z(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n343) );
  XNOR2_X1 U364 ( .A(n312), .B(n343), .ZN(n534) );
  XOR2_X1 U365 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT23), .B(KEYINPUT91), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n328) );
  XOR2_X1 U368 ( .A(G204GAT), .B(G211GAT), .Z(n316) );
  XNOR2_X1 U369 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n433) );
  XOR2_X1 U371 ( .A(n433), .B(KEYINPUT22), .Z(n318) );
  NAND2_X1 U372 ( .A1(G228GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U374 ( .A(n319), .B(G218GAT), .Z(n321) );
  XOR2_X1 U375 ( .A(G141GAT), .B(G22GAT), .Z(n405) );
  XNOR2_X1 U376 ( .A(G50GAT), .B(n405), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n324) );
  XOR2_X1 U378 ( .A(G155GAT), .B(KEYINPUT3), .Z(n323) );
  XNOR2_X1 U379 ( .A(KEYINPUT2), .B(KEYINPUT90), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n340) );
  XOR2_X1 U381 ( .A(n324), .B(n340), .Z(n326) );
  XOR2_X1 U382 ( .A(G162GAT), .B(G106GAT), .Z(n350) );
  XOR2_X1 U383 ( .A(G148GAT), .B(G78GAT), .Z(n397) );
  XNOR2_X1 U384 ( .A(n350), .B(n397), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n328), .B(n327), .ZN(n465) );
  XOR2_X1 U387 ( .A(G57GAT), .B(KEYINPUT5), .Z(n330) );
  XNOR2_X1 U388 ( .A(G1GAT), .B(KEYINPUT92), .ZN(n329) );
  XNOR2_X1 U389 ( .A(n330), .B(n329), .ZN(n338) );
  NAND2_X1 U390 ( .A1(G225GAT), .A2(G233GAT), .ZN(n336) );
  XOR2_X1 U391 ( .A(KEYINPUT4), .B(G148GAT), .Z(n332) );
  XNOR2_X1 U392 ( .A(G29GAT), .B(G141GAT), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U394 ( .A(G162GAT), .B(G85GAT), .Z(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U398 ( .A(n339), .B(KEYINPUT6), .Z(n342) );
  XNOR2_X1 U399 ( .A(n340), .B(KEYINPUT1), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n518) );
  XOR2_X1 U402 ( .A(KEYINPUT8), .B(G50GAT), .Z(n346) );
  XNOR2_X1 U403 ( .A(G43GAT), .B(G29GAT), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U405 ( .A(KEYINPUT7), .B(n347), .ZN(n414) );
  XOR2_X1 U406 ( .A(KEYINPUT67), .B(KEYINPUT77), .Z(n349) );
  XNOR2_X1 U407 ( .A(G134GAT), .B(KEYINPUT68), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U409 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n352) );
  XOR2_X1 U410 ( .A(G99GAT), .B(G85GAT), .Z(n384) );
  XNOR2_X1 U411 ( .A(n350), .B(n384), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n356) );
  AND2_X1 U414 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n362) );
  XOR2_X1 U416 ( .A(G92GAT), .B(G218GAT), .Z(n358) );
  XNOR2_X1 U417 ( .A(G36GAT), .B(G190GAT), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n435) );
  XNOR2_X1 U419 ( .A(n435), .B(KEYINPUT10), .ZN(n360) );
  XOR2_X1 U420 ( .A(n414), .B(n363), .Z(n558) );
  XNOR2_X1 U421 ( .A(n558), .B(KEYINPUT78), .ZN(n453) );
  XNOR2_X1 U422 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n453), .B(n364), .ZN(n488) );
  XOR2_X1 U424 ( .A(G15GAT), .B(G1GAT), .Z(n402) );
  XNOR2_X1 U425 ( .A(G71GAT), .B(G57GAT), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n365), .B(KEYINPUT13), .ZN(n390) );
  XOR2_X1 U427 ( .A(n402), .B(n390), .Z(n367) );
  NAND2_X1 U428 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n382) );
  XOR2_X1 U430 ( .A(KEYINPUT81), .B(KEYINPUT15), .Z(n369) );
  XNOR2_X1 U431 ( .A(KEYINPUT82), .B(KEYINPUT14), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U433 ( .A(KEYINPUT12), .B(G64GAT), .Z(n371) );
  XNOR2_X1 U434 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n380) );
  XOR2_X1 U437 ( .A(KEYINPUT83), .B(G155GAT), .Z(n375) );
  XNOR2_X1 U438 ( .A(G127GAT), .B(G78GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U440 ( .A(G183GAT), .B(KEYINPUT79), .Z(n438) );
  XOR2_X1 U441 ( .A(n376), .B(n438), .Z(n378) );
  XNOR2_X1 U442 ( .A(G22GAT), .B(G211GAT), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n576) );
  NOR2_X1 U446 ( .A1(n488), .A2(n576), .ZN(n383) );
  XNOR2_X1 U447 ( .A(KEYINPUT45), .B(n383), .ZN(n418) );
  XOR2_X1 U448 ( .A(G176GAT), .B(G64GAT), .Z(n431) );
  XOR2_X1 U449 ( .A(n431), .B(n384), .Z(n386) );
  NAND2_X1 U450 ( .A1(G230GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n393) );
  XOR2_X1 U452 ( .A(KEYINPUT33), .B(KEYINPUT76), .Z(n388) );
  XNOR2_X1 U453 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U456 ( .A(G92GAT), .B(G106GAT), .Z(n395) );
  XNOR2_X1 U457 ( .A(G120GAT), .B(G204GAT), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n573) );
  XOR2_X1 U461 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n401) );
  XNOR2_X1 U462 ( .A(G197GAT), .B(KEYINPUT72), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n413) );
  XOR2_X1 U464 ( .A(G113GAT), .B(G36GAT), .Z(n404) );
  XOR2_X1 U465 ( .A(G169GAT), .B(G8GAT), .Z(n432) );
  XNOR2_X1 U466 ( .A(n402), .B(n432), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n406) );
  XOR2_X1 U468 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U469 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n408) );
  NAND2_X1 U470 ( .A1(G229GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U472 ( .A(KEYINPUT71), .B(n409), .ZN(n410) );
  XNOR2_X1 U473 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n568) );
  XNOR2_X1 U476 ( .A(KEYINPUT73), .B(n568), .ZN(n560) );
  INV_X1 U477 ( .A(n560), .ZN(n416) );
  AND2_X1 U478 ( .A1(n573), .A2(n416), .ZN(n417) );
  AND2_X1 U479 ( .A1(n418), .A2(n417), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n419), .B(KEYINPUT113), .ZN(n427) );
  INV_X1 U481 ( .A(n576), .ZN(n563) );
  NOR2_X1 U482 ( .A1(n551), .A2(n568), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n420), .B(KEYINPUT46), .ZN(n421) );
  NOR2_X1 U484 ( .A1(n563), .A2(n421), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n422), .B(KEYINPUT111), .ZN(n423) );
  NOR2_X1 U486 ( .A1(n558), .A2(n423), .ZN(n425) );
  NAND2_X1 U487 ( .A1(n427), .A2(n426), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n442) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U491 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U492 ( .A1(G226GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n520) );
  XOR2_X1 U495 ( .A(KEYINPUT120), .B(n520), .Z(n443) );
  NOR2_X1 U496 ( .A1(n529), .A2(n443), .ZN(n444) );
  XOR2_X1 U497 ( .A(KEYINPUT54), .B(n444), .Z(n445) );
  NAND2_X1 U498 ( .A1(n465), .A2(n567), .ZN(n447) );
  INV_X1 U499 ( .A(n551), .ZN(n537) );
  NAND2_X1 U500 ( .A1(n564), .A2(n537), .ZN(n452) );
  XOR2_X1 U501 ( .A(G176GAT), .B(KEYINPUT123), .Z(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(G1349GAT) );
  NAND2_X1 U505 ( .A1(n564), .A2(n453), .ZN(n457) );
  XOR2_X1 U506 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n455) );
  INV_X1 U507 ( .A(G190GAT), .ZN(n454) );
  NAND2_X1 U508 ( .A1(n560), .A2(n573), .ZN(n493) );
  XNOR2_X1 U509 ( .A(n520), .B(KEYINPUT27), .ZN(n467) );
  NAND2_X1 U510 ( .A1(n467), .A2(n518), .ZN(n458) );
  XOR2_X1 U511 ( .A(KEYINPUT93), .B(n458), .Z(n530) );
  XNOR2_X1 U512 ( .A(KEYINPUT28), .B(n465), .ZN(n532) );
  NAND2_X1 U513 ( .A1(n532), .A2(n534), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n530), .A2(n459), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT94), .ZN(n473) );
  XOR2_X1 U516 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n464) );
  INV_X1 U517 ( .A(n534), .ZN(n522) );
  NAND2_X1 U518 ( .A1(n522), .A2(n520), .ZN(n461) );
  XOR2_X1 U519 ( .A(KEYINPUT95), .B(n461), .Z(n462) );
  NAND2_X1 U520 ( .A1(n462), .A2(n465), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n464), .B(n463), .ZN(n469) );
  NOR2_X1 U522 ( .A1(n465), .A2(n522), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n466), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U524 ( .A1(n566), .A2(n467), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U526 ( .A(KEYINPUT97), .B(n470), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n471), .A2(n518), .ZN(n472) );
  NOR2_X1 U528 ( .A1(n473), .A2(n472), .ZN(n489) );
  NOR2_X1 U529 ( .A1(n453), .A2(n576), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT16), .B(n474), .Z(n475) );
  XNOR2_X1 U531 ( .A(n475), .B(KEYINPUT84), .ZN(n476) );
  OR2_X1 U532 ( .A1(n489), .A2(n476), .ZN(n505) );
  NOR2_X1 U533 ( .A1(n493), .A2(n505), .ZN(n486) );
  NAND2_X1 U534 ( .A1(n518), .A2(n486), .ZN(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(n477), .ZN(n478) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n478), .ZN(G1324GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n480) );
  NAND2_X1 U538 ( .A1(n486), .A2(n520), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U540 ( .A(G8GAT), .B(n481), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n483) );
  NAND2_X1 U542 ( .A1(n486), .A2(n522), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(n485) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT100), .Z(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  INV_X1 U546 ( .A(n532), .ZN(n526) );
  NAND2_X1 U547 ( .A1(n526), .A2(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .Z(n496) );
  XOR2_X1 U550 ( .A(KEYINPUT37), .B(KEYINPUT104), .Z(n492) );
  NOR2_X1 U551 ( .A1(n488), .A2(n489), .ZN(n490) );
  NAND2_X1 U552 ( .A1(n490), .A2(n576), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(n517) );
  NOR2_X1 U554 ( .A1(n493), .A2(n517), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(KEYINPUT38), .ZN(n502) );
  NAND2_X1 U556 ( .A1(n518), .A2(n502), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U558 ( .A(KEYINPUT102), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n502), .A2(n520), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n500) );
  NAND2_X1 U562 ( .A1(n522), .A2(n502), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n504) );
  NAND2_X1 U566 ( .A1(n526), .A2(n502), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n508) );
  NAND2_X1 U569 ( .A1(n568), .A2(n537), .ZN(n516) );
  OR2_X1 U570 ( .A1(n505), .A2(n516), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(KEYINPUT107), .ZN(n513) );
  NAND2_X1 U572 ( .A1(n518), .A2(n513), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n510) );
  NAND2_X1 U575 ( .A1(n513), .A2(n520), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n511), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n522), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U581 ( .A1(n513), .A2(n526), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n518), .A2(n525), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n525), .A2(n520), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n522), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(KEYINPUT110), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  XOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT115), .Z(n536) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT114), .ZN(n549) );
  NAND2_X1 U597 ( .A1(n532), .A2(n549), .ZN(n533) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n545), .A2(n560), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n539) );
  NAND2_X1 U602 ( .A1(n545), .A2(n537), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(n540), .ZN(G1341GAT) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n544) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n542) );
  NAND2_X1 U607 ( .A1(n545), .A2(n563), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n547) );
  NAND2_X1 U611 ( .A1(n545), .A2(n453), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U613 ( .A(G134GAT), .B(n548), .Z(G1343GAT) );
  NAND2_X1 U614 ( .A1(n566), .A2(n549), .ZN(n556) );
  NOR2_X1 U615 ( .A1(n568), .A2(n556), .ZN(n550) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n550), .Z(G1344GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n556), .ZN(n553) );
  XNOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U621 ( .A1(n576), .A2(n556), .ZN(n555) );
  XOR2_X1 U622 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  INV_X1 U623 ( .A(n556), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n560), .A2(n564), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n579) );
  NOR2_X1 U632 ( .A1(n579), .A2(n568), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n573), .A2(n579), .ZN(n575) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n579), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(n577), .Z(n578) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n488), .A2(n579), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

