

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(G164), .A2(G1384), .ZN(n704) );
  BUF_X2 U550 ( .A(n864), .Z(n513) );
  XOR2_X1 U551 ( .A(KEYINPUT17), .B(n532), .Z(n864) );
  NOR2_X1 U552 ( .A1(G168), .A2(n743), .ZN(n744) );
  AND2_X1 U553 ( .A1(n767), .A2(n989), .ZN(n768) );
  XOR2_X1 U554 ( .A(n732), .B(KEYINPUT29), .Z(n514) );
  NOR2_X1 U555 ( .A1(n751), .A2(n739), .ZN(n740) );
  INV_X1 U556 ( .A(KEYINPUT28), .ZN(n710) );
  NAND2_X1 U557 ( .A1(n762), .A2(G8), .ZN(n763) );
  XNOR2_X1 U558 ( .A(n763), .B(KEYINPUT32), .ZN(n764) );
  AND2_X1 U559 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U560 ( .A1(G8), .A2(n756), .ZN(n784) );
  NOR2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  NOR2_X1 U562 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U563 ( .A1(G651), .A2(n622), .ZN(n641) );
  BUF_X1 U564 ( .A(n675), .Z(G160) );
  XOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .Z(n622) );
  NAND2_X1 U566 ( .A1(G51), .A2(n641), .ZN(n517) );
  INV_X1 U567 ( .A(G651), .ZN(n520) );
  NOR2_X1 U568 ( .A1(G543), .A2(n520), .ZN(n515) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n515), .Z(n637) );
  NAND2_X1 U570 ( .A1(G63), .A2(n637), .ZN(n516) );
  NAND2_X1 U571 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U572 ( .A(KEYINPUT6), .B(n518), .ZN(n525) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n633) );
  NAND2_X1 U574 ( .A1(n633), .A2(G89), .ZN(n519) );
  XNOR2_X1 U575 ( .A(n519), .B(KEYINPUT4), .ZN(n522) );
  NOR2_X1 U576 ( .A1(n622), .A2(n520), .ZN(n634) );
  NAND2_X1 U577 ( .A1(G76), .A2(n634), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U579 ( .A(n523), .B(KEYINPUT5), .Z(n524) );
  NOR2_X1 U580 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U581 ( .A(KEYINPUT72), .B(n526), .Z(n527) );
  XNOR2_X1 U582 ( .A(KEYINPUT7), .B(n527), .ZN(G168) );
  INV_X1 U583 ( .A(G2105), .ZN(n528) );
  NOR2_X2 U584 ( .A1(G2104), .A2(n528), .ZN(n867) );
  NAND2_X1 U585 ( .A1(n867), .A2(G125), .ZN(n531) );
  AND2_X1 U586 ( .A1(n528), .A2(G2104), .ZN(n863) );
  NAND2_X1 U587 ( .A1(G101), .A2(n863), .ZN(n529) );
  XOR2_X1 U588 ( .A(KEYINPUT23), .B(n529), .Z(n530) );
  NAND2_X1 U589 ( .A1(n531), .A2(n530), .ZN(n536) );
  NAND2_X1 U590 ( .A1(G137), .A2(n513), .ZN(n534) );
  AND2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n869) );
  NAND2_X1 U592 ( .A1(G113), .A2(n869), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n675) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U596 ( .A1(G99), .A2(n863), .ZN(n538) );
  NAND2_X1 U597 ( .A1(G111), .A2(n869), .ZN(n537) );
  NAND2_X1 U598 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U599 ( .A(KEYINPUT77), .B(n539), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n867), .A2(G123), .ZN(n540) );
  XNOR2_X1 U601 ( .A(n540), .B(KEYINPUT18), .ZN(n542) );
  NAND2_X1 U602 ( .A1(G135), .A2(n513), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U604 ( .A(KEYINPUT76), .B(n543), .Z(n544) );
  NAND2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n902) );
  XNOR2_X1 U606 ( .A(G2096), .B(n902), .ZN(n546) );
  OR2_X1 U607 ( .A1(G2100), .A2(n546), .ZN(G156) );
  INV_X1 U608 ( .A(G108), .ZN(G238) );
  NAND2_X1 U609 ( .A1(G52), .A2(n641), .ZN(n548) );
  NAND2_X1 U610 ( .A1(G64), .A2(n637), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G90), .A2(n633), .ZN(n550) );
  NAND2_X1 U613 ( .A1(G77), .A2(n634), .ZN(n549) );
  NAND2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(n551), .Z(n552) );
  NOR2_X1 U616 ( .A1(n553), .A2(n552), .ZN(G171) );
  NAND2_X1 U617 ( .A1(n633), .A2(G88), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(KEYINPUT82), .ZN(n556) );
  NAND2_X1 U619 ( .A1(G62), .A2(n637), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G75), .A2(n634), .ZN(n558) );
  NAND2_X1 U622 ( .A1(G50), .A2(n641), .ZN(n557) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n560), .A2(n559), .ZN(G166) );
  AND2_X1 U625 ( .A1(G102), .A2(n863), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G126), .A2(n867), .ZN(n562) );
  NAND2_X1 U627 ( .A1(G114), .A2(n869), .ZN(n561) );
  AND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U629 ( .A1(G138), .A2(n864), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(G164) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U634 ( .A(G567), .ZN(n670) );
  NOR2_X1 U635 ( .A1(n670), .A2(G223), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT11), .ZN(G234) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n570) );
  NAND2_X1 U638 ( .A1(G56), .A2(n637), .ZN(n569) );
  XNOR2_X1 U639 ( .A(n570), .B(n569), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n634), .A2(G68), .ZN(n571) );
  XNOR2_X1 U641 ( .A(KEYINPUT71), .B(n571), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n633), .A2(G81), .ZN(n572) );
  XOR2_X1 U643 ( .A(KEYINPUT12), .B(n572), .Z(n573) );
  NOR2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U645 ( .A(n575), .B(KEYINPUT13), .ZN(n576) );
  NOR2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n641), .A2(G43), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n975) );
  INV_X1 U649 ( .A(G860), .ZN(n601) );
  OR2_X1 U650 ( .A1(n975), .A2(n601), .ZN(G153) );
  INV_X1 U651 ( .A(G171), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G79), .A2(n634), .ZN(n581) );
  NAND2_X1 U654 ( .A1(G66), .A2(n637), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G92), .A2(n633), .ZN(n583) );
  NAND2_X1 U657 ( .A1(G54), .A2(n641), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U660 ( .A(KEYINPUT15), .B(n586), .Z(n983) );
  OR2_X1 U661 ( .A1(n983), .A2(G868), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(G284) );
  XOR2_X1 U663 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U664 ( .A1(G91), .A2(n633), .ZN(n589) );
  XNOR2_X1 U665 ( .A(n589), .B(KEYINPUT66), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G53), .A2(n641), .ZN(n590) );
  XOR2_X1 U667 ( .A(KEYINPUT67), .B(n590), .Z(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G78), .A2(n634), .ZN(n594) );
  NAND2_X1 U670 ( .A1(G65), .A2(n637), .ZN(n593) );
  NAND2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n986) );
  XOR2_X1 U673 ( .A(n986), .B(KEYINPUT68), .Z(G299) );
  INV_X1 U674 ( .A(G868), .ZN(n653) );
  NOR2_X1 U675 ( .A1(G286), .A2(n653), .ZN(n597) );
  XOR2_X1 U676 ( .A(KEYINPUT73), .B(n597), .Z(n599) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U679 ( .A(KEYINPUT74), .B(n600), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n602), .A2(n983), .ZN(n603) );
  XNOR2_X1 U682 ( .A(n603), .B(KEYINPUT16), .ZN(n604) );
  XOR2_X1 U683 ( .A(KEYINPUT75), .B(n604), .Z(G148) );
  NOR2_X1 U684 ( .A1(G868), .A2(n975), .ZN(n607) );
  NAND2_X1 U685 ( .A1(G868), .A2(n983), .ZN(n605) );
  NOR2_X1 U686 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U687 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G559), .A2(n983), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n608), .B(n975), .ZN(n650) );
  NOR2_X1 U690 ( .A1(n650), .A2(G860), .ZN(n617) );
  NAND2_X1 U691 ( .A1(G80), .A2(n634), .ZN(n610) );
  NAND2_X1 U692 ( .A1(G67), .A2(n637), .ZN(n609) );
  NAND2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U694 ( .A1(G93), .A2(n633), .ZN(n611) );
  XNOR2_X1 U695 ( .A(KEYINPUT79), .B(n611), .ZN(n612) );
  NOR2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n641), .A2(G55), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n652) );
  XOR2_X1 U699 ( .A(n652), .B(KEYINPUT78), .Z(n616) );
  XNOR2_X1 U700 ( .A(n617), .B(n616), .ZN(G145) );
  NAND2_X1 U701 ( .A1(G49), .A2(n641), .ZN(n619) );
  NAND2_X1 U702 ( .A1(G74), .A2(G651), .ZN(n618) );
  NAND2_X1 U703 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U704 ( .A1(n637), .A2(n620), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n621), .B(KEYINPUT80), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G87), .A2(n622), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U708 ( .A1(G73), .A2(n634), .ZN(n625) );
  XNOR2_X1 U709 ( .A(n625), .B(KEYINPUT2), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G86), .A2(n633), .ZN(n627) );
  NAND2_X1 U711 ( .A1(G48), .A2(n641), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U713 ( .A1(G61), .A2(n637), .ZN(n628) );
  XNOR2_X1 U714 ( .A(KEYINPUT81), .B(n628), .ZN(n629) );
  NOR2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U717 ( .A1(G85), .A2(n633), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G72), .A2(n634), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U720 ( .A1(G60), .A2(n637), .ZN(n638) );
  XNOR2_X1 U721 ( .A(KEYINPUT65), .B(n638), .ZN(n639) );
  NOR2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n641), .A2(G47), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(G290) );
  XNOR2_X1 U725 ( .A(G299), .B(G288), .ZN(n649) );
  XNOR2_X1 U726 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n645) );
  XNOR2_X1 U727 ( .A(G305), .B(G166), .ZN(n644) );
  XNOR2_X1 U728 ( .A(n645), .B(n644), .ZN(n646) );
  XOR2_X1 U729 ( .A(n646), .B(G290), .Z(n647) );
  XNOR2_X1 U730 ( .A(n652), .B(n647), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n649), .B(n648), .ZN(n887) );
  XNOR2_X1 U732 ( .A(n650), .B(n887), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n651), .A2(G868), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U736 ( .A(KEYINPUT84), .B(n656), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n657) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n658), .ZN(n660) );
  XOR2_X1 U740 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n659) );
  XNOR2_X1 U741 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U742 ( .A1(G2072), .A2(n661), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U744 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  NAND2_X1 U745 ( .A1(G132), .A2(G82), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n662), .B(KEYINPUT86), .ZN(n663) );
  XNOR2_X1 U747 ( .A(n663), .B(KEYINPUT22), .ZN(n664) );
  NOR2_X1 U748 ( .A1(G218), .A2(n664), .ZN(n665) );
  NAND2_X1 U749 ( .A1(G96), .A2(n665), .ZN(n812) );
  NAND2_X1 U750 ( .A1(G2106), .A2(n812), .ZN(n666) );
  XNOR2_X1 U751 ( .A(n666), .B(KEYINPUT87), .ZN(n672) );
  NAND2_X1 U752 ( .A1(G120), .A2(G69), .ZN(n667) );
  NOR2_X1 U753 ( .A1(G237), .A2(n667), .ZN(n668) );
  XOR2_X1 U754 ( .A(KEYINPUT88), .B(n668), .Z(n669) );
  NOR2_X1 U755 ( .A1(G238), .A2(n669), .ZN(n814) );
  NOR2_X1 U756 ( .A1(n670), .A2(n814), .ZN(n671) );
  NOR2_X1 U757 ( .A1(n672), .A2(n671), .ZN(G319) );
  INV_X1 U758 ( .A(G319), .ZN(n892) );
  NAND2_X1 U759 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U760 ( .A1(n892), .A2(n673), .ZN(n674) );
  XOR2_X1 U761 ( .A(KEYINPUT89), .B(n674), .Z(n811) );
  NAND2_X1 U762 ( .A1(n811), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U764 ( .A(G1986), .B(G290), .ZN(n988) );
  NAND2_X1 U765 ( .A1(n675), .A2(G40), .ZN(n703) );
  NOR2_X1 U766 ( .A1(n704), .A2(n703), .ZN(n803) );
  NAND2_X1 U767 ( .A1(n988), .A2(n803), .ZN(n793) );
  XNOR2_X1 U768 ( .A(KEYINPUT37), .B(G2067), .ZN(n801) );
  NAND2_X1 U769 ( .A1(G104), .A2(n863), .ZN(n677) );
  NAND2_X1 U770 ( .A1(G140), .A2(n513), .ZN(n676) );
  NAND2_X1 U771 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n678), .ZN(n683) );
  NAND2_X1 U773 ( .A1(G116), .A2(n869), .ZN(n680) );
  NAND2_X1 U774 ( .A1(G128), .A2(n867), .ZN(n679) );
  NAND2_X1 U775 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U776 ( .A(KEYINPUT35), .B(n681), .Z(n682) );
  NOR2_X1 U777 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U778 ( .A(KEYINPUT36), .B(n684), .ZN(n883) );
  NOR2_X1 U779 ( .A1(n801), .A2(n883), .ZN(n912) );
  NAND2_X1 U780 ( .A1(n803), .A2(n912), .ZN(n799) );
  NAND2_X1 U781 ( .A1(G95), .A2(n863), .ZN(n686) );
  NAND2_X1 U782 ( .A1(G131), .A2(n513), .ZN(n685) );
  NAND2_X1 U783 ( .A1(n686), .A2(n685), .ZN(n690) );
  NAND2_X1 U784 ( .A1(G107), .A2(n869), .ZN(n688) );
  NAND2_X1 U785 ( .A1(G119), .A2(n867), .ZN(n687) );
  NAND2_X1 U786 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U787 ( .A1(n690), .A2(n689), .ZN(n878) );
  INV_X1 U788 ( .A(G1991), .ZN(n953) );
  NOR2_X1 U789 ( .A1(n878), .A2(n953), .ZN(n699) );
  NAND2_X1 U790 ( .A1(G117), .A2(n869), .ZN(n692) );
  NAND2_X1 U791 ( .A1(G129), .A2(n867), .ZN(n691) );
  NAND2_X1 U792 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n863), .A2(G105), .ZN(n693) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n693), .Z(n694) );
  NOR2_X1 U795 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U796 ( .A1(n513), .A2(G141), .ZN(n696) );
  NAND2_X1 U797 ( .A1(n697), .A2(n696), .ZN(n879) );
  AND2_X1 U798 ( .A1(n879), .A2(G1996), .ZN(n698) );
  NOR2_X1 U799 ( .A1(n699), .A2(n698), .ZN(n898) );
  INV_X1 U800 ( .A(n803), .ZN(n700) );
  NOR2_X1 U801 ( .A1(n898), .A2(n700), .ZN(n796) );
  INV_X1 U802 ( .A(n796), .ZN(n701) );
  NAND2_X1 U803 ( .A1(n799), .A2(n701), .ZN(n702) );
  XNOR2_X1 U804 ( .A(n702), .B(KEYINPUT90), .ZN(n791) );
  INV_X1 U805 ( .A(n703), .ZN(n705) );
  NAND2_X2 U806 ( .A1(n705), .A2(n704), .ZN(n756) );
  NOR2_X1 U807 ( .A1(G2084), .A2(n756), .ZN(n739) );
  NAND2_X1 U808 ( .A1(G8), .A2(n739), .ZN(n754) );
  XOR2_X1 U809 ( .A(KEYINPUT92), .B(n756), .Z(n733) );
  NAND2_X1 U810 ( .A1(G2072), .A2(n733), .ZN(n706) );
  XNOR2_X1 U811 ( .A(n706), .B(KEYINPUT27), .ZN(n709) );
  XNOR2_X1 U812 ( .A(KEYINPUT93), .B(G1956), .ZN(n931) );
  NOR2_X1 U813 ( .A1(n733), .A2(n931), .ZN(n707) );
  XNOR2_X1 U814 ( .A(n707), .B(KEYINPUT94), .ZN(n708) );
  NOR2_X1 U815 ( .A1(n709), .A2(n708), .ZN(n712) );
  NOR2_X1 U816 ( .A1(n986), .A2(n712), .ZN(n711) );
  XNOR2_X1 U817 ( .A(n711), .B(n710), .ZN(n731) );
  NAND2_X1 U818 ( .A1(n986), .A2(n712), .ZN(n729) );
  INV_X1 U819 ( .A(n756), .ZN(n735) );
  AND2_X1 U820 ( .A1(n735), .A2(G1996), .ZN(n715) );
  XNOR2_X1 U821 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n713) );
  XNOR2_X1 U822 ( .A(n713), .B(KEYINPUT64), .ZN(n714) );
  XNOR2_X1 U823 ( .A(n715), .B(n714), .ZN(n717) );
  NAND2_X1 U824 ( .A1(n756), .A2(G1341), .ZN(n716) );
  NAND2_X1 U825 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U826 ( .A1(n975), .A2(n718), .ZN(n720) );
  NOR2_X1 U827 ( .A1(n720), .A2(n983), .ZN(n719) );
  XNOR2_X1 U828 ( .A(n719), .B(KEYINPUT97), .ZN(n727) );
  NAND2_X1 U829 ( .A1(n720), .A2(n983), .ZN(n725) );
  NAND2_X1 U830 ( .A1(G2067), .A2(n733), .ZN(n722) );
  NAND2_X1 U831 ( .A1(G1348), .A2(n756), .ZN(n721) );
  NAND2_X1 U832 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U833 ( .A(KEYINPUT96), .B(n723), .ZN(n724) );
  NAND2_X1 U834 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U835 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U836 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U837 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U838 ( .A(G2078), .B(KEYINPUT25), .Z(n956) );
  INV_X1 U839 ( .A(n733), .ZN(n734) );
  NOR2_X1 U840 ( .A1(n956), .A2(n734), .ZN(n737) );
  NOR2_X1 U841 ( .A1(n735), .A2(G1961), .ZN(n736) );
  NOR2_X1 U842 ( .A1(n737), .A2(n736), .ZN(n745) );
  OR2_X1 U843 ( .A1(n745), .A2(G301), .ZN(n738) );
  NAND2_X1 U844 ( .A1(n514), .A2(n738), .ZN(n750) );
  NOR2_X1 U845 ( .A1(G1966), .A2(n784), .ZN(n751) );
  XNOR2_X1 U846 ( .A(KEYINPUT98), .B(n740), .ZN(n741) );
  NAND2_X1 U847 ( .A1(n741), .A2(G8), .ZN(n742) );
  XNOR2_X1 U848 ( .A(KEYINPUT30), .B(n742), .ZN(n743) );
  XNOR2_X1 U849 ( .A(n744), .B(KEYINPUT99), .ZN(n747) );
  NAND2_X1 U850 ( .A1(n745), .A2(G301), .ZN(n746) );
  NAND2_X1 U851 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U852 ( .A(KEYINPUT31), .B(n748), .ZN(n749) );
  NAND2_X1 U853 ( .A1(n750), .A2(n749), .ZN(n755) );
  XOR2_X1 U854 ( .A(n755), .B(KEYINPUT100), .Z(n752) );
  NOR2_X1 U855 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U856 ( .A1(n754), .A2(n753), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n755), .A2(G286), .ZN(n761) );
  NOR2_X1 U858 ( .A1(G1971), .A2(n784), .ZN(n758) );
  NOR2_X1 U859 ( .A1(G2090), .A2(n756), .ZN(n757) );
  NOR2_X1 U860 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U861 ( .A1(n759), .A2(G303), .ZN(n760) );
  NAND2_X1 U862 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U863 ( .A1(n765), .A2(n764), .ZN(n781) );
  NOR2_X1 U864 ( .A1(G1976), .A2(G288), .ZN(n774) );
  NOR2_X1 U865 ( .A1(G1971), .A2(G303), .ZN(n766) );
  NOR2_X1 U866 ( .A1(n774), .A2(n766), .ZN(n990) );
  NAND2_X1 U867 ( .A1(n781), .A2(n990), .ZN(n769) );
  INV_X1 U868 ( .A(n784), .ZN(n767) );
  NAND2_X1 U869 ( .A1(G1976), .A2(G288), .ZN(n989) );
  NOR2_X2 U870 ( .A1(KEYINPUT33), .A2(n770), .ZN(n771) );
  XNOR2_X1 U871 ( .A(n771), .B(KEYINPUT101), .ZN(n773) );
  XOR2_X1 U872 ( .A(KEYINPUT102), .B(G1981), .Z(n772) );
  XNOR2_X1 U873 ( .A(G305), .B(n772), .ZN(n977) );
  NAND2_X1 U874 ( .A1(n773), .A2(n977), .ZN(n777) );
  NAND2_X1 U875 ( .A1(KEYINPUT33), .A2(n774), .ZN(n775) );
  NOR2_X1 U876 ( .A1(n784), .A2(n775), .ZN(n776) );
  NOR2_X1 U877 ( .A1(n777), .A2(n776), .ZN(n789) );
  NOR2_X1 U878 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XOR2_X1 U879 ( .A(n778), .B(KEYINPUT24), .Z(n779) );
  NOR2_X1 U880 ( .A1(n784), .A2(n779), .ZN(n780) );
  XNOR2_X1 U881 ( .A(n780), .B(KEYINPUT91), .ZN(n787) );
  NOR2_X1 U882 ( .A1(G2090), .A2(G303), .ZN(n782) );
  NAND2_X1 U883 ( .A1(G8), .A2(n782), .ZN(n783) );
  NAND2_X1 U884 ( .A1(n781), .A2(n783), .ZN(n785) );
  NAND2_X1 U885 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U886 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n806) );
  NOR2_X1 U889 ( .A1(G1996), .A2(n879), .ZN(n905) );
  AND2_X1 U890 ( .A1(n953), .A2(n878), .ZN(n901) );
  NOR2_X1 U891 ( .A1(G1986), .A2(G290), .ZN(n794) );
  NOR2_X1 U892 ( .A1(n901), .A2(n794), .ZN(n795) );
  NOR2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U894 ( .A1(n905), .A2(n797), .ZN(n798) );
  XNOR2_X1 U895 ( .A(n798), .B(KEYINPUT39), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n801), .A2(n883), .ZN(n909) );
  NAND2_X1 U898 ( .A1(n802), .A2(n909), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U901 ( .A(KEYINPUT40), .B(n807), .ZN(G329) );
  INV_X1 U902 ( .A(G223), .ZN(n808) );
  NAND2_X1 U903 ( .A1(G2106), .A2(n808), .ZN(G217) );
  AND2_X1 U904 ( .A1(G15), .A2(G2), .ZN(n809) );
  NAND2_X1 U905 ( .A1(G661), .A2(n809), .ZN(G259) );
  NAND2_X1 U906 ( .A1(G3), .A2(G1), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(G188) );
  XOR2_X1 U908 ( .A(G69), .B(KEYINPUT104), .Z(G235) );
  INV_X1 U910 ( .A(G132), .ZN(G219) );
  INV_X1 U911 ( .A(G120), .ZN(G236) );
  INV_X1 U912 ( .A(G82), .ZN(G220) );
  INV_X1 U913 ( .A(n812), .ZN(n813) );
  NAND2_X1 U914 ( .A1(n814), .A2(n813), .ZN(G261) );
  INV_X1 U915 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U916 ( .A(G1348), .B(G2454), .ZN(n815) );
  XNOR2_X1 U917 ( .A(n815), .B(G2430), .ZN(n816) );
  XNOR2_X1 U918 ( .A(n816), .B(G1341), .ZN(n822) );
  XOR2_X1 U919 ( .A(G2443), .B(G2427), .Z(n818) );
  XNOR2_X1 U920 ( .A(G2438), .B(G2446), .ZN(n817) );
  XNOR2_X1 U921 ( .A(n818), .B(n817), .ZN(n820) );
  XOR2_X1 U922 ( .A(G2451), .B(G2435), .Z(n819) );
  XNOR2_X1 U923 ( .A(n820), .B(n819), .ZN(n821) );
  XNOR2_X1 U924 ( .A(n822), .B(n821), .ZN(n823) );
  NAND2_X1 U925 ( .A1(n823), .A2(G14), .ZN(n824) );
  XNOR2_X1 U926 ( .A(KEYINPUT103), .B(n824), .ZN(G401) );
  XOR2_X1 U927 ( .A(KEYINPUT105), .B(G1971), .Z(n826) );
  XNOR2_X1 U928 ( .A(G1986), .B(G1976), .ZN(n825) );
  XNOR2_X1 U929 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U930 ( .A(n827), .B(KEYINPUT41), .Z(n829) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n828) );
  XNOR2_X1 U932 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U933 ( .A(G1956), .B(G1961), .Z(n831) );
  XNOR2_X1 U934 ( .A(G1981), .B(G1966), .ZN(n830) );
  XNOR2_X1 U935 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U936 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U937 ( .A(G2474), .B(KEYINPUT106), .ZN(n834) );
  XNOR2_X1 U938 ( .A(n835), .B(n834), .ZN(G229) );
  XOR2_X1 U939 ( .A(G2100), .B(G2096), .Z(n837) );
  XNOR2_X1 U940 ( .A(KEYINPUT42), .B(G2678), .ZN(n836) );
  XNOR2_X1 U941 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U942 ( .A(KEYINPUT43), .B(G2090), .Z(n839) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U944 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U945 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U946 ( .A(G2084), .B(G2078), .ZN(n842) );
  XNOR2_X1 U947 ( .A(n843), .B(n842), .ZN(G227) );
  NAND2_X1 U948 ( .A1(G124), .A2(n867), .ZN(n844) );
  XNOR2_X1 U949 ( .A(n844), .B(KEYINPUT44), .ZN(n846) );
  NAND2_X1 U950 ( .A1(n863), .A2(G100), .ZN(n845) );
  NAND2_X1 U951 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U952 ( .A1(G136), .A2(n513), .ZN(n848) );
  NAND2_X1 U953 ( .A1(G112), .A2(n869), .ZN(n847) );
  NAND2_X1 U954 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U955 ( .A1(n850), .A2(n849), .ZN(G162) );
  XOR2_X1 U956 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n861) );
  NAND2_X1 U957 ( .A1(G118), .A2(n869), .ZN(n852) );
  NAND2_X1 U958 ( .A1(G130), .A2(n867), .ZN(n851) );
  NAND2_X1 U959 ( .A1(n852), .A2(n851), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G106), .A2(n863), .ZN(n854) );
  NAND2_X1 U961 ( .A1(G142), .A2(n513), .ZN(n853) );
  NAND2_X1 U962 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U963 ( .A(KEYINPUT107), .B(n855), .ZN(n856) );
  XNOR2_X1 U964 ( .A(KEYINPUT45), .B(n856), .ZN(n857) );
  NOR2_X1 U965 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U966 ( .A(n859), .B(KEYINPUT110), .ZN(n860) );
  XNOR2_X1 U967 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U968 ( .A(n902), .B(n862), .ZN(n877) );
  NAND2_X1 U969 ( .A1(G103), .A2(n863), .ZN(n866) );
  NAND2_X1 U970 ( .A1(G139), .A2(n513), .ZN(n865) );
  NAND2_X1 U971 ( .A1(n866), .A2(n865), .ZN(n875) );
  NAND2_X1 U972 ( .A1(n867), .A2(G127), .ZN(n868) );
  XNOR2_X1 U973 ( .A(n868), .B(KEYINPUT108), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G115), .A2(n869), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U976 ( .A(KEYINPUT47), .B(n872), .ZN(n873) );
  XNOR2_X1 U977 ( .A(KEYINPUT109), .B(n873), .ZN(n874) );
  NOR2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n914) );
  XNOR2_X1 U979 ( .A(G164), .B(n914), .ZN(n876) );
  XNOR2_X1 U980 ( .A(n877), .B(n876), .ZN(n885) );
  XOR2_X1 U981 ( .A(G162), .B(n878), .Z(n881) );
  XOR2_X1 U982 ( .A(G160), .B(n879), .Z(n880) );
  XNOR2_X1 U983 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U984 ( .A(n883), .B(n882), .Z(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U986 ( .A1(G37), .A2(n886), .ZN(G395) );
  XNOR2_X1 U987 ( .A(G286), .B(n887), .ZN(n889) );
  XNOR2_X1 U988 ( .A(G171), .B(n983), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U990 ( .A(n890), .B(n975), .Z(n891) );
  NOR2_X1 U991 ( .A1(G37), .A2(n891), .ZN(G397) );
  OR2_X1 U992 ( .A1(n892), .A2(G401), .ZN(n895) );
  NOR2_X1 U993 ( .A1(G229), .A2(G227), .ZN(n893) );
  XNOR2_X1 U994 ( .A(KEYINPUT49), .B(n893), .ZN(n894) );
  NOR2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n897) );
  NOR2_X1 U996 ( .A1(G395), .A2(G397), .ZN(n896) );
  NAND2_X1 U997 ( .A1(n897), .A2(n896), .ZN(G225) );
  INV_X1 U998 ( .A(G225), .ZN(G308) );
  INV_X1 U999 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U1000 ( .A(G160), .B(G2084), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(n899), .A2(n898), .ZN(n900) );
  NOR2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n908) );
  XOR2_X1 U1004 ( .A(G2090), .B(G162), .Z(n904) );
  NOR2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(KEYINPUT51), .B(n906), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(KEYINPUT111), .B(n913), .Z(n921) );
  XOR2_X1 U1011 ( .A(G2072), .B(n914), .Z(n915) );
  XNOR2_X1 U1012 ( .A(KEYINPUT112), .B(n915), .ZN(n918) );
  XOR2_X1 U1013 ( .A(G164), .B(G2078), .Z(n917) );
  NOR2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(KEYINPUT50), .B(n919), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(KEYINPUT52), .B(n922), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n923), .A2(G29), .ZN(n1010) );
  XOR2_X1 U1019 ( .A(G1966), .B(G21), .Z(n936) );
  XNOR2_X1 U1020 ( .A(KEYINPUT123), .B(G1341), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(n924), .B(G19), .ZN(n930) );
  XOR2_X1 U1022 ( .A(G4), .B(KEYINPUT124), .Z(n926) );
  XNOR2_X1 U1023 ( .A(G1348), .B(KEYINPUT59), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n926), .B(n925), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(G1981), .B(G6), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1028 ( .A(G20), .B(n931), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(KEYINPUT60), .B(n934), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(KEYINPUT122), .B(G1961), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(G5), .B(n937), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(KEYINPUT125), .B(n940), .ZN(n948) );
  XOR2_X1 U1036 ( .A(G1986), .B(G24), .Z(n944) );
  XNOR2_X1 U1037 ( .A(G1976), .B(G23), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(G1971), .B(G22), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(KEYINPUT58), .B(n945), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT126), .B(n946), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(n949), .B(KEYINPUT61), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(G16), .B(KEYINPUT121), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(G11), .A2(n952), .ZN(n1008) );
  XNOR2_X1 U1048 ( .A(n953), .B(G25), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n954), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n955), .B(KEYINPUT113), .ZN(n965) );
  XOR2_X1 U1051 ( .A(n956), .B(G27), .Z(n961) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G2072), .B(G33), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(n959), .B(KEYINPUT114), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G32), .B(G1996), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n966), .B(KEYINPUT53), .ZN(n969) );
  XOR2_X1 U1061 ( .A(G2084), .B(G34), .Z(n967) );
  XNOR2_X1 U1062 ( .A(KEYINPUT54), .B(n967), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(G35), .B(G2090), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1066 ( .A(KEYINPUT115), .B(n972), .Z(n973) );
  NOR2_X1 U1067 ( .A1(G29), .A2(n973), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(KEYINPUT55), .B(n974), .ZN(n1006) );
  XNOR2_X1 U1069 ( .A(n975), .B(G1341), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(KEYINPUT119), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(KEYINPUT116), .B(KEYINPUT57), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(G168), .B(G1966), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(n980), .B(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n1001) );
  XNOR2_X1 U1076 ( .A(n983), .B(G1348), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(G171), .B(G1961), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n998) );
  XOR2_X1 U1079 ( .A(n986), .B(G1956), .Z(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n996) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n993) );
  INV_X1 U1082 ( .A(G1971), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(G166), .A2(n991), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1085 ( .A(KEYINPUT117), .B(n994), .Z(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT118), .B(n999), .Z(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(G16), .B(KEYINPUT56), .Z(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1092 ( .A(KEYINPUT120), .B(n1004), .Z(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(n1011), .B(KEYINPUT127), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(KEYINPUT62), .B(n1012), .ZN(G311) );
  INV_X1 U1098 ( .A(G311), .ZN(G150) );
endmodule

