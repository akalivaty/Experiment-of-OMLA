//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  NAND2_X1  g001(.A1(G234), .A2(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G952), .A3(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT21), .B(G898), .Z(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(G902), .A3(G953), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(G210), .B1(G237), .B2(G902), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G128), .Z(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT64), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n196), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n195), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(new_n200), .A3(new_n196), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n197), .A2(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n197), .A2(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n201), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n202), .A3(G128), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n216), .B1(new_n204), .B2(new_n205), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n214), .A2(new_n217), .B1(new_n209), .B2(new_n216), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT87), .B1(new_n218), .B2(new_n212), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n214), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n209), .A2(new_n216), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT87), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G125), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT88), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n225), .A2(new_n226), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n213), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G224), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G953), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n229), .B(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G104), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT3), .B1(new_n233), .B2(G107), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n235));
  INV_X1    g049(.A(G107), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G104), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(G107), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G101), .ZN(new_n240));
  INV_X1    g054(.A(G101), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n234), .A2(new_n237), .A3(new_n241), .A4(new_n238), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(KEYINPUT4), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT76), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT76), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n240), .A2(new_n245), .A3(KEYINPUT4), .A4(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(G116), .B(G119), .Z(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT2), .B(G113), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n239), .A2(new_n251), .A3(G101), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(KEYINPUT77), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT83), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n257));
  INV_X1    g071(.A(G119), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G116), .ZN(new_n259));
  OAI211_X1 g073(.A(G113), .B(new_n259), .C1(new_n248), .C2(new_n257), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n248), .B2(new_n249), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n236), .A2(G104), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n238), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G101), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT78), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT78), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n266), .A3(G101), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n242), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n247), .A2(KEYINPUT83), .A3(new_n250), .A4(new_n253), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n256), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g088(.A(G110), .B(G122), .Z(new_n275));
  XOR2_X1   g089(.A(new_n275), .B(KEYINPUT85), .Z(new_n276));
  NAND4_X1  g090(.A1(new_n256), .A2(KEYINPUT84), .A3(new_n270), .A4(new_n271), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n272), .A2(new_n275), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n274), .A2(new_n281), .A3(new_n276), .A4(new_n277), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT86), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n232), .B(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT89), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n282), .B(new_n283), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n289), .A2(KEYINPUT89), .A3(new_n232), .A4(new_n280), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n225), .A2(new_n213), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT7), .B1(new_n230), .B2(G953), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n295), .A2(KEYINPUT91), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(KEYINPUT91), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(new_n275), .B(KEYINPUT8), .Z(new_n299));
  AND2_X1   g113(.A1(new_n261), .A2(new_n268), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n269), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n301), .A2(KEYINPUT90), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(KEYINPUT90), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n298), .A2(new_n279), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n229), .A2(new_n294), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n292), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n194), .B1(new_n291), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n194), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n309), .B(new_n306), .C1(new_n288), .C2(new_n290), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n187), .B(new_n193), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G128), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(G119), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT66), .B(G128), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT23), .ZN(new_n317));
  OR3_X1    g131(.A1(new_n258), .A2(KEYINPUT23), .A3(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G110), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT16), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(G125), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n212), .A2(new_n323), .ZN(new_n325));
  NOR2_X1   g139(.A1(G125), .A2(G140), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n324), .B1(new_n327), .B2(new_n322), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(G146), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT24), .B(G110), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n195), .B2(new_n258), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(new_n332), .B2(new_n316), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n330), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n320), .A2(new_n319), .B1(new_n334), .B2(new_n331), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT72), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n198), .A2(new_n200), .ZN(new_n338));
  INV_X1    g152(.A(new_n327), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n336), .A2(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n328), .A2(new_n197), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n319), .A2(new_n320), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n334), .A2(new_n331), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n341), .B1(new_n344), .B2(KEYINPUT72), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n340), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n340), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n335), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G137), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n350), .B(new_n351), .Z(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n352), .B(new_n353), .Z(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n335), .B(new_n354), .C1(new_n347), .C2(new_n348), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n292), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT25), .A4(new_n292), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT70), .B(G217), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(G234), .B2(new_n292), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n365), .B2(new_n358), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n207), .A2(new_n210), .ZN(new_n368));
  INV_X1    g182(.A(G134), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G137), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n369), .A2(G137), .ZN(new_n372));
  OAI21_X1  g186(.A(G131), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT11), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n369), .B2(G137), .ZN(new_n375));
  INV_X1    g189(.A(G137), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT11), .A3(G134), .ZN(new_n377));
  INV_X1    g191(.A(G131), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n375), .A2(new_n377), .A3(new_n378), .A4(new_n370), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n368), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(new_n370), .A3(new_n377), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G131), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n379), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n218), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n250), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(KEYINPUT28), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT65), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n373), .B2(new_n379), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n373), .A2(new_n391), .A3(new_n379), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n386), .B1(new_n211), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n250), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n399));
  INV_X1    g213(.A(G237), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n189), .A3(G210), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n399), .B(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(G101), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT67), .ZN(new_n407));
  INV_X1    g221(.A(new_n394), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(new_n392), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n409), .A2(new_n368), .B1(new_n385), .B2(new_n218), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n407), .B1(new_n410), .B2(KEYINPUT30), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n396), .A2(KEYINPUT67), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n382), .A2(KEYINPUT30), .A3(new_n386), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n411), .A2(new_n413), .A3(new_n250), .A4(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n389), .A3(new_n404), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT31), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT31), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n415), .A2(new_n418), .A3(new_n389), .A4(new_n404), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n419), .A2(KEYINPUT69), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(KEYINPUT69), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n406), .B(new_n417), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(G472), .A2(G902), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT32), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT32), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n404), .B1(new_n398), .B2(KEYINPUT29), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n387), .A2(new_n388), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n390), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n292), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n415), .A2(new_n389), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n405), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT29), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G472), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n367), .B1(new_n428), .B2(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n265), .A2(new_n242), .A3(new_n267), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n368), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n313), .B1(new_n205), .B2(KEYINPUT1), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n209), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n268), .B1(new_n441), .B2(new_n210), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n385), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT12), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n444), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT81), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n449));
  OR2_X1    g263(.A1(new_n442), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n368), .A2(new_n438), .A3(KEYINPUT10), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n247), .A2(new_n218), .A3(new_n253), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n385), .B(KEYINPUT80), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G140), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n189), .A2(G227), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n455), .B(new_n456), .Z(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT81), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n445), .A2(new_n460), .A3(new_n446), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n448), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT82), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n459), .A2(new_n461), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT82), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n465), .A3(new_n448), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n457), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n469), .A2(new_n385), .ZN(new_n470));
  INV_X1    g284(.A(new_n454), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G469), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n292), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n292), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n447), .A2(new_n454), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n468), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n470), .A2(new_n458), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(G469), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n475), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT9), .B(G234), .Z(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G221), .B1(new_n484), .B2(G902), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(G113), .B(G122), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(new_n233), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n327), .A2(KEYINPUT93), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(KEYINPUT19), .Z(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT64), .B(G146), .ZN(new_n491));
  OR3_X1    g305(.A1(new_n490), .A2(KEYINPUT94), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT94), .B1(new_n490), .B2(new_n491), .ZN(new_n493));
  INV_X1    g307(.A(new_n341), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n400), .A2(new_n189), .A3(G214), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(G143), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(new_n378), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n496), .A2(new_n378), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT18), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n496), .B1(new_n501), .B2(new_n378), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n327), .A2(G146), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n491), .B2(new_n327), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n488), .B1(new_n498), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n499), .A2(KEYINPUT17), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n329), .B(new_n509), .C1(new_n497), .C2(KEYINPUT17), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n488), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G475), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n292), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n488), .B1(new_n507), .B2(new_n510), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n292), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G475), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n514), .A4(new_n292), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G478), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT13), .B1(new_n315), .B2(G143), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(new_n369), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n313), .A2(G143), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n315), .B2(G143), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n526), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G116), .B(G122), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(new_n236), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n236), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n533), .B(KEYINPUT95), .Z(new_n534));
  INV_X1    g348(.A(G116), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT14), .A3(G122), .ZN(new_n536));
  INV_X1    g350(.A(new_n530), .ZN(new_n537));
  OAI211_X1 g351(.A(G107), .B(new_n536), .C1(new_n537), .C2(KEYINPUT14), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n528), .A2(G134), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n528), .A2(G134), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n534), .A2(new_n538), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n484), .A2(G953), .A3(new_n364), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT96), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n532), .A2(new_n541), .A3(new_n543), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n542), .A2(KEYINPUT96), .A3(new_n544), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n292), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n524), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n524), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(new_n553), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n522), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n486), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n312), .A2(new_n437), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(G101), .ZN(G3));
  XNOR2_X1  g374(.A(new_n542), .B(KEYINPUT98), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n544), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(KEYINPUT99), .A3(new_n544), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n564), .A2(KEYINPUT33), .A3(new_n547), .A4(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT33), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n548), .A2(new_n567), .A3(new_n549), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n566), .A2(G478), .A3(new_n292), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n550), .A2(new_n523), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT100), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n367), .ZN(new_n576));
  INV_X1    g390(.A(G472), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n422), .B2(new_n292), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n423), .B2(new_n422), .ZN(new_n579));
  AND4_X1   g393(.A1(new_n576), .A2(new_n482), .A3(new_n485), .A4(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n312), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT34), .B(G104), .Z(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(G6));
  NOR2_X1   g397(.A1(new_n573), .A2(new_n556), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n312), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G107), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT101), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n585), .B(new_n587), .ZN(G9));
  INV_X1    g402(.A(new_n579), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n349), .A2(KEYINPUT36), .A3(new_n354), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n356), .A2(new_n357), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n354), .A2(KEYINPUT36), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n365), .A2(G902), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n362), .A2(new_n365), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OR3_X1    g409(.A1(new_n589), .A2(KEYINPUT102), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT102), .B1(new_n589), .B2(new_n595), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n312), .A2(new_n596), .A3(new_n558), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT37), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n320), .ZN(G12));
  INV_X1    g414(.A(new_n556), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n190), .B1(new_n192), .B2(G900), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n601), .A2(new_n522), .A3(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n187), .B(new_n603), .C1(new_n308), .C2(new_n310), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n428), .A2(new_n436), .ZN(new_n606));
  INV_X1    g420(.A(new_n595), .ZN(new_n607));
  AND4_X1   g421(.A1(new_n606), .A2(new_n485), .A3(new_n482), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT103), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n313), .ZN(G30));
  NAND2_X1  g425(.A1(new_n291), .A2(new_n307), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n309), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n291), .A2(new_n194), .A3(new_n307), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT38), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n602), .B(KEYINPUT39), .Z(new_n617));
  OR2_X1    g431(.A1(new_n486), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT40), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n595), .A3(new_n619), .ZN(new_n620));
  OR3_X1    g434(.A1(new_n486), .A2(KEYINPUT40), .A3(new_n617), .ZN(new_n621));
  INV_X1    g435(.A(new_n428), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n433), .A2(new_n405), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n430), .A2(new_n405), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n625), .B2(new_n389), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n577), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n601), .A2(new_n573), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n621), .A2(new_n187), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n620), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n196), .ZN(G45));
  INV_X1    g448(.A(new_n486), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n606), .A3(new_n607), .ZN(new_n636));
  INV_X1    g450(.A(new_n187), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n613), .B2(new_n614), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n572), .A2(new_n573), .A3(new_n602), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n187), .B(new_n640), .C1(new_n308), .C2(new_n310), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n636), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n197), .ZN(G48));
  NAND2_X1  g459(.A1(new_n606), .A2(new_n576), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n470), .A2(new_n471), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n463), .A2(new_n466), .B1(new_n647), .B2(new_n468), .ZN(new_n648));
  OAI21_X1  g462(.A(G469), .B1(new_n648), .B2(G902), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n475), .A2(new_n649), .A3(new_n485), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n312), .A2(new_n652), .A3(new_n575), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT41), .B(G113), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G15));
  NAND3_X1  g469(.A1(new_n312), .A2(new_n652), .A3(new_n584), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G116), .ZN(G18));
  OAI211_X1 g471(.A(new_n650), .B(new_n187), .C1(new_n308), .C2(new_n310), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n193), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n557), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n659), .A2(new_n606), .A3(new_n607), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G119), .ZN(G21));
  NAND2_X1  g477(.A1(new_n431), .A2(new_n405), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n664), .B(new_n417), .C1(new_n420), .C2(new_n421), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n423), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT105), .ZN(new_n667));
  INV_X1    g481(.A(new_n578), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n576), .A2(new_n667), .A3(new_n193), .A4(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n659), .A2(new_n631), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G122), .ZN(G24));
  NAND3_X1  g486(.A1(new_n667), .A2(new_n668), .A3(new_n607), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n638), .A2(new_n674), .A3(new_n640), .A4(new_n650), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G125), .ZN(G27));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n308), .A2(new_n310), .A3(new_n637), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(new_n437), .A3(new_n635), .ZN(new_n679));
  INV_X1    g493(.A(new_n640), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n677), .B(KEYINPUT42), .C1(new_n679), .C2(new_n680), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n378), .ZN(G33));
  NAND3_X1  g500(.A1(new_n613), .A2(new_n187), .A3(new_n614), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n646), .A3(new_n486), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n584), .A2(new_n602), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n690), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n688), .A2(KEYINPUT108), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n678), .A2(new_n693), .A3(new_n437), .A4(new_n635), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n695), .B1(new_n696), .B2(new_n691), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G134), .ZN(G36));
  NAND2_X1  g513(.A1(new_n522), .A2(new_n572), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n589), .A3(new_n607), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n687), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n479), .A2(new_n480), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n479), .A2(KEYINPUT45), .A3(new_n480), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(G469), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(KEYINPUT46), .A3(new_n477), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n475), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n475), .A2(new_n711), .A3(KEYINPUT109), .ZN(new_n715));
  INV_X1    g529(.A(new_n710), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n476), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n714), .B(new_n715), .C1(KEYINPUT46), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n485), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n617), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n705), .B(new_n720), .C1(new_n704), .C2(new_n703), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT110), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G137), .ZN(G39));
  NAND3_X1  g537(.A1(new_n428), .A2(new_n367), .A3(new_n436), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n687), .A2(new_n680), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT111), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n719), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n718), .A2(KEYINPUT47), .A3(new_n485), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n323), .ZN(G42));
  NAND3_X1  g546(.A1(new_n576), .A2(new_n667), .A3(new_n668), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n190), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n702), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT117), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n650), .A2(new_n637), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n616), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n739), .B(new_n740), .C1(new_n737), .C2(new_n738), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n735), .A2(new_n678), .A3(new_n702), .A4(new_n650), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT118), .ZN(new_n747));
  OR3_X1    g561(.A1(new_n747), .A2(KEYINPUT119), .A3(new_n673), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT119), .B1(new_n747), .B2(new_n673), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n475), .A2(new_n649), .ZN(new_n751));
  INV_X1    g565(.A(new_n485), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n730), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n736), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n678), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n678), .A2(new_n628), .A3(new_n650), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n757), .A2(new_n367), .A3(new_n190), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n522), .A3(new_n571), .A4(new_n569), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n745), .A2(new_n750), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n747), .A2(new_n646), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT48), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(G952), .B(new_n189), .C1(new_n736), .C2(new_n658), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n758), .B2(new_n575), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT120), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(KEYINPUT120), .A3(new_n769), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n763), .B(new_n764), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n608), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n642), .A2(new_n651), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n777), .A2(new_n674), .B1(new_n605), .B2(new_n608), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n595), .A2(new_n779), .A3(new_n602), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(new_n595), .B2(new_n602), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n486), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n638), .A3(new_n629), .A4(new_n631), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(new_n778), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n776), .A2(new_n778), .A3(KEYINPUT52), .A4(new_n783), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n674), .A2(new_n635), .A3(new_n575), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n636), .B2(new_n557), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n602), .A3(new_n678), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n698), .A2(new_n683), .A3(new_n684), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n609), .A2(new_n675), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n644), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(KEYINPUT115), .A3(KEYINPUT52), .A4(new_n783), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n638), .A2(KEYINPUT113), .A3(new_n193), .A4(new_n584), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n799));
  INV_X1    g613(.A(new_n584), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n799), .B1(new_n311), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(new_n801), .A3(new_n580), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n559), .A3(new_n581), .A4(new_n598), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n662), .A2(new_n671), .A3(new_n653), .A4(new_n656), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n789), .A2(new_n794), .A3(new_n797), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n805), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n598), .A2(new_n559), .A3(new_n581), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(KEYINPUT53), .A3(new_n802), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n793), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(KEYINPUT116), .A3(new_n797), .A4(new_n789), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n805), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n658), .A2(new_n630), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n311), .A2(new_n574), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n670), .A2(new_n817), .B1(new_n818), .B2(new_n652), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(KEYINPUT112), .A3(new_n656), .A4(new_n662), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n803), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n786), .A2(new_n788), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n794), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n804), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n809), .A2(new_n814), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n823), .A2(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n789), .A2(new_n797), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n821), .A2(new_n794), .A3(new_n804), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n827), .B(KEYINPUT54), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n773), .A2(new_n831), .B1(G952), .B2(G953), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n751), .B(KEYINPUT49), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n700), .A2(new_n367), .A3(new_n637), .A4(new_n752), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n740), .A2(new_n628), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n832), .A2(new_n835), .ZN(G75));
  NAND3_X1  g650(.A1(new_n809), .A2(new_n824), .A3(new_n814), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(G210), .A3(G902), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n289), .A2(new_n280), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(new_n232), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT55), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n838), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n838), .B2(new_n839), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n189), .A2(G952), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G51));
  NAND2_X1  g660(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n826), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n476), .B(KEYINPUT57), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n473), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n837), .A2(G902), .A3(new_n716), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n845), .B1(new_n851), .B2(new_n852), .ZN(G54));
  INV_X1    g667(.A(new_n845), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n837), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n855));
  INV_X1    g669(.A(new_n513), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT121), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n855), .A2(new_n860), .A3(new_n856), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n857), .B1(new_n859), .B2(new_n861), .ZN(G60));
  AND2_X1   g676(.A1(new_n566), .A2(new_n568), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n848), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(G478), .A2(G902), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT59), .Z(new_n866));
  NOR2_X1   g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n866), .B1(new_n826), .B2(new_n830), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n854), .B1(new_n868), .B2(new_n863), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n867), .A2(new_n869), .ZN(G63));
  NAND2_X1  g684(.A1(G217), .A2(G902), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT60), .Z(new_n872));
  NAND2_X1  g686(.A1(new_n837), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n591), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n837), .A2(new_n593), .A3(new_n872), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n854), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n874), .A2(KEYINPUT61), .A3(new_n854), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(G66));
  AOI21_X1  g694(.A(new_n189), .B1(new_n191), .B2(G224), .ZN(new_n881));
  INV_X1    g695(.A(new_n821), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n882), .B2(new_n189), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT122), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n840), .B1(G898), .B2(new_n189), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n884), .B(new_n885), .ZN(G69));
  NAND3_X1  g700(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(new_n490), .Z(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(G900), .B2(G953), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n721), .A2(new_n796), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT125), .Z(new_n891));
  INV_X1    g705(.A(new_n731), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n685), .B1(new_n697), .B2(new_n694), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n720), .A2(new_n437), .A3(new_n638), .A4(new_n631), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(new_n895), .B2(G953), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT62), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n776), .A2(new_n778), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n633), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(KEYINPUT62), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n796), .B1(new_n632), .B2(new_n620), .ZN(new_n903));
  INV_X1    g717(.A(new_n898), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n731), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n618), .B1(new_n574), .B2(new_n800), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n437), .A3(new_n678), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n902), .A2(new_n905), .A3(new_n721), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n189), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n888), .B(KEYINPUT123), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n896), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n912), .B(new_n915), .Z(G72));
  NAND2_X1  g730(.A1(G472), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT63), .Z(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n895), .B2(new_n882), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n433), .A3(new_n405), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n624), .A2(new_n434), .A3(new_n918), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n827), .B(new_n921), .C1(new_n828), .C2(new_n829), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n854), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n918), .B1(new_n908), .B2(new_n882), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT127), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n623), .B2(new_n925), .ZN(G57));
endmodule


