//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT23), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G169gat), .Z(new_n220));
  AND2_X1   g019(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT25), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT23), .ZN(new_n225));
  OR2_X1    g024(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n227));
  AOI21_X1  g026(.A(G190gat), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n217), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n210), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT25), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n214), .A2(KEYINPUT27), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT27), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(G183gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n233), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(G183gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n214), .A2(KEYINPUT27), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT68), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n232), .B1(new_n241), .B2(new_n215), .ZN(new_n242));
  AND2_X1   g041(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT27), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(KEYINPUT67), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(new_n235), .A3(G183gat), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n245), .A2(new_n246), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n209), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n224), .A2(KEYINPUT26), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(new_n254), .A3(new_n211), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n223), .B(new_n231), .C1(new_n242), .C2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n257));
  INV_X1    g056(.A(G120gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(G113gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260));
  INV_X1    g059(.A(G113gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(G120gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n258), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n259), .A2(new_n262), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n266));
  XNOR2_X1  g065(.A(G127gat), .B(G134gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n267), .ZN(new_n269));
  XNOR2_X1  g068(.A(G113gat), .B(G120gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n269), .B1(KEYINPUT1), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n205), .B1(new_n256), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n274), .B(KEYINPUT64), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n252), .A2(new_n253), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n247), .A2(new_n249), .ZN(new_n278));
  INV_X1    g077(.A(new_n246), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT66), .B(G183gat), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(KEYINPUT27), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(G190gat), .B1(new_n237), .B2(new_n240), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n282), .B(new_n211), .C1(new_n232), .C2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n272), .ZN(new_n285));
  AOI22_X1  g084(.A1(KEYINPUT25), .A2(new_n230), .B1(new_n219), .B2(new_n222), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n284), .A2(KEYINPUT71), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n256), .A2(new_n272), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n273), .A2(new_n276), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n289), .B(KEYINPUT34), .Z(new_n290));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n288), .A3(new_n287), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n275), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT33), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(KEYINPUT32), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(G71gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(G99gat), .ZN(new_n296));
  XOR2_X1   g095(.A(G15gat), .B(G43gat), .Z(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(KEYINPUT33), .ZN(new_n300));
  AND4_X1   g099(.A1(KEYINPUT73), .A2(new_n292), .A3(KEYINPUT32), .A4(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(new_n291), .B2(new_n275), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT73), .B1(new_n303), .B2(new_n300), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n290), .B(new_n299), .C1(new_n301), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n292), .A2(KEYINPUT32), .A3(new_n300), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n303), .A2(KEYINPUT73), .A3(new_n300), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n290), .B1(new_n311), .B2(new_n299), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n203), .B(new_n204), .C1(new_n306), .C2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n299), .B1(new_n301), .B2(new_n304), .ZN(new_n314));
  INV_X1    g113(.A(new_n290), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n316), .A2(KEYINPUT74), .A3(new_n202), .A4(new_n305), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT77), .ZN(new_n320));
  INV_X1    g119(.A(G141gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(G148gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(G148gat), .ZN(new_n323));
  INV_X1    g122(.A(G148gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  INV_X1    g126(.A(G155gat), .ZN(new_n328));
  INV_X1    g127(.A(G162gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n327), .B1(new_n330), .B2(KEYINPUT2), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n327), .ZN(new_n333));
  NOR2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G141gat), .B(G148gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(KEYINPUT2), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n332), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n272), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n272), .B2(new_n338), .ZN(new_n344));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346));
  INV_X1    g145(.A(new_n323), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n321), .A2(G148gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n349), .A2(new_n335), .B1(new_n326), .B2(new_n331), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n350), .A2(KEYINPUT4), .A3(new_n271), .A4(new_n268), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n342), .A2(new_n344), .A3(new_n345), .A4(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT5), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n353), .A2(KEYINPUT78), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n272), .A2(new_n338), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n350), .A2(new_n271), .A3(new_n268), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n345), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(new_n353), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n352), .B(new_n354), .C1(new_n353), .C2(new_n358), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT0), .B(G57gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(G85gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G1gat), .B(G29gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n360), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n360), .B2(new_n361), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n368));
  NOR3_X1   g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n360), .A2(new_n361), .A3(new_n365), .ZN(new_n370));
  INV_X1    g169(.A(new_n368), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n319), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n367), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(new_n370), .A3(new_n371), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT80), .ZN(new_n376));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n256), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n377), .B1(new_n284), .B2(new_n286), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT75), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G197gat), .B(G204gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT22), .ZN(new_n384));
  INV_X1    g183(.A(G211gat), .ZN(new_n385));
  INV_X1    g184(.A(G218gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(G211gat), .B(G218gat), .Z(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT75), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n284), .B2(new_n286), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(new_n378), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n382), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n390), .B1(new_n380), .B2(new_n381), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT76), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G8gat), .ZN(new_n401));
  INV_X1    g200(.A(G36gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n397), .A2(new_n398), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n397), .A2(new_n404), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n395), .A2(new_n396), .A3(new_n403), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(KEYINPUT30), .A3(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n373), .A2(new_n376), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n379), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n350), .B1(new_n411), .B2(new_n340), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n390), .B1(new_n379), .B2(new_n341), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n340), .B1(new_n411), .B2(KEYINPUT81), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n390), .B2(new_n379), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n338), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n413), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n414), .B1(new_n420), .B2(new_n410), .ZN(new_n421));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT31), .B(G50gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(KEYINPUT82), .A3(G22gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(G22gat), .B2(new_n424), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n421), .B(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n369), .A2(new_n372), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n382), .A2(new_n390), .A3(new_n394), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(new_n391), .C1(new_n380), .C2(new_n381), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n391), .B1(new_n380), .B2(new_n381), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT84), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT37), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n397), .B2(new_n439), .ZN(new_n440));
  AOI211_X1 g239(.A(KEYINPUT85), .B(KEYINPUT37), .C1(new_n395), .C2(new_n396), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n403), .B(new_n437), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT38), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n406), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n397), .A2(new_n439), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(new_n443), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n446), .B(new_n403), .C1(new_n440), .C2(new_n441), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n430), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n342), .A2(new_n344), .A3(new_n351), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(G225gat), .A3(G233gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n356), .A2(new_n345), .A3(new_n357), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(KEYINPUT39), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n365), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT83), .B(KEYINPUT39), .Z(new_n454));
  OAI211_X1 g253(.A(new_n452), .B(new_n453), .C1(new_n450), .C2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT40), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n408), .A2(new_n370), .A3(new_n405), .A4(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n455), .A2(new_n456), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n428), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI221_X1 g259(.A(new_n318), .B1(new_n409), .B2(new_n428), .C1(new_n448), .C2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT35), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n408), .A2(new_n405), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n463), .A2(new_n316), .A3(new_n428), .A4(new_n305), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n464), .B2(new_n429), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n316), .A2(new_n428), .A3(new_n305), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(KEYINPUT35), .A3(new_n409), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT93), .B(G211gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(G231gat), .A2(G233gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT89), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT16), .ZN(new_n477));
  AOI21_X1  g276(.A(G1gat), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G8gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n478), .A2(new_n479), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n478), .A2(new_n479), .ZN(new_n484));
  INV_X1    g283(.A(new_n476), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n480), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G71gat), .A2(G78gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT9), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(G57gat), .A2(G64gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(G57gat), .A2(G64gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT92), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(G71gat), .B2(G78gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G71gat), .B(G78gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n493), .A2(new_n497), .A3(new_n495), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT21), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(G183gat), .ZN(new_n504));
  XOR2_X1   g303(.A(G127gat), .B(G155gat), .Z(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n503), .B(new_n214), .ZN(new_n507));
  INV_X1    g306(.A(new_n505), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n474), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(new_n509), .A3(new_n474), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n501), .A2(KEYINPUT21), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n513), .B(new_n514), .Z(new_n515));
  NAND3_X1  g314(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n515), .ZN(new_n517));
  INV_X1    g316(.A(new_n512), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n510), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G99gat), .B(G106gat), .Z(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G85gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT95), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT95), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G85gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G92gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n527), .A2(new_n528), .B1(KEYINPUT8), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n522), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(KEYINPUT8), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT95), .B(G85gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(G92gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT7), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n531), .B(new_n537), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n536), .A2(new_n521), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G29gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(new_n402), .ZN(new_n542));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(KEYINPUT15), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n402), .A3(KEYINPUT14), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT14), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT87), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT87), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT15), .ZN(new_n552));
  INV_X1    g351(.A(G43gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(G50gat), .ZN(new_n554));
  INV_X1    g353(.A(G50gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(G43gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n552), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n544), .A2(new_n549), .A3(new_n551), .A4(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(KEYINPUT15), .B(new_n543), .C1(new_n548), .C2(new_n542), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n561), .A2(KEYINPUT88), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(KEYINPUT88), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n558), .A2(KEYINPUT88), .A3(new_n561), .A4(new_n559), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n540), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G190gat), .B(G218gat), .Z(new_n568));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n540), .A2(new_n560), .B1(KEYINPUT41), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n568), .ZN(new_n573));
  INV_X1    g372(.A(new_n571), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n566), .ZN(new_n575));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT94), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n572), .A2(KEYINPUT96), .A3(new_n575), .A4(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n575), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(KEYINPUT96), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n567), .A2(new_n568), .A3(new_n571), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT97), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n581), .A2(new_n582), .A3(new_n587), .A4(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n520), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n470), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n564), .A2(new_n565), .B1(new_n486), .B2(new_n483), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n483), .A2(new_n486), .A3(new_n560), .ZN(new_n593));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT90), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT18), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n599));
  INV_X1    g398(.A(new_n565), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n487), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n593), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n602), .A3(new_n594), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT18), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(KEYINPUT90), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n560), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n487), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n594), .B(KEYINPUT91), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n598), .A2(new_n605), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G169gat), .B(G197gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n598), .A2(new_n605), .A3(new_n611), .A4(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n493), .A2(new_n497), .A3(new_n495), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n497), .B1(new_n493), .B2(new_n495), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n539), .B2(new_n533), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n530), .A2(new_n522), .A3(new_n532), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n521), .B1(new_n536), .B2(new_n538), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n501), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n540), .A2(KEYINPUT10), .A3(new_n501), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n627), .A2(new_n630), .ZN(new_n637));
  INV_X1    g436(.A(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(new_n207), .ZN(new_n642));
  INV_X1    g441(.A(G204gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n639), .A2(KEYINPUT98), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n644), .B1(new_n639), .B2(KEYINPUT98), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n647), .A2(new_n636), .A3(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n623), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n591), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n373), .A2(new_n376), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT99), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n373), .A2(new_n655), .A3(new_n376), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660));
  INV_X1    g459(.A(new_n463), .ZN(new_n661));
  NOR2_X1   g460(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n591), .A2(new_n651), .A3(new_n661), .A4(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n477), .A2(new_n479), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n664), .A2(new_n660), .A3(new_n665), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n479), .B1(new_n652), .B2(new_n661), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(G1325gat));
  NOR2_X1   g472(.A1(new_n306), .A2(new_n312), .ZN(new_n674));
  AOI21_X1  g473(.A(G15gat), .B1(new_n652), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n313), .A2(new_n317), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n652), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(G15gat), .B2(new_n677), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n652), .A2(new_n427), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(new_n589), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n651), .A2(new_n520), .ZN(new_n683));
  AOI211_X1 g482(.A(new_n682), .B(new_n683), .C1(new_n461), .C2(new_n469), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n541), .A3(new_n657), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT45), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n468), .A2(KEYINPUT102), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n465), .A2(new_n467), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n444), .A2(new_n447), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n429), .ZN(new_n692));
  INV_X1    g491(.A(new_n460), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n676), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n409), .B2(new_n428), .ZN(new_n696));
  INV_X1    g495(.A(new_n376), .ZN(new_n697));
  INV_X1    g496(.A(new_n372), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT80), .B1(new_n375), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n463), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(KEYINPUT101), .A3(new_n427), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n688), .A2(new_n690), .B1(new_n694), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n687), .B1(new_n703), .B2(new_n682), .ZN(new_n704));
  INV_X1    g503(.A(new_n683), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n470), .A2(KEYINPUT44), .A3(new_n589), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n657), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n686), .A2(new_n709), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n684), .A2(new_n402), .A3(new_n661), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT46), .Z(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n707), .B2(new_n463), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1329gat));
  OAI21_X1  g513(.A(G43gat), .B1(new_n707), .B2(new_n318), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n684), .A2(new_n553), .A3(new_n674), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT103), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n717), .A2(KEYINPUT103), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT104), .Z(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n719), .B(new_n722), .ZN(G1330gat));
  OAI21_X1  g522(.A(G50gat), .B1(new_n707), .B2(new_n428), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n684), .A2(new_n555), .A3(new_n427), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT48), .B1(new_n725), .B2(KEYINPUT105), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1331gat));
  AND3_X1   g527(.A1(new_n465), .A2(new_n467), .A3(new_n689), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n689), .B1(new_n465), .B2(new_n467), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n317), .B(new_n313), .C1(new_n448), .C2(new_n460), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n696), .A2(new_n701), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n729), .A2(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n520), .A2(new_n622), .A3(new_n589), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n650), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n708), .A2(KEYINPUT106), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n657), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g540(.A1(new_n735), .A2(new_n463), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  INV_X1    g545(.A(new_n735), .ZN(new_n747));
  INV_X1    g546(.A(G71gat), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n674), .B(KEYINPUT107), .Z(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G71gat), .B1(new_n735), .B2(new_n318), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g552(.A1(new_n735), .A2(new_n428), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT108), .B(G78gat), .Z(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1335gat));
  INV_X1    g555(.A(new_n520), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n622), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n733), .A2(new_n589), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n589), .A4(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n657), .A3(new_n650), .ZN(new_n764));
  AOI211_X1 g563(.A(new_n687), .B(new_n682), .C1(new_n461), .C2(new_n469), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT44), .B1(new_n733), .B2(new_n589), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n758), .A2(new_n650), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n708), .A2(new_n527), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n764), .A2(new_n527), .B1(new_n768), .B2(new_n769), .ZN(G1336gat));
  NOR2_X1   g569(.A1(new_n463), .A2(G92gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n688), .A2(new_n690), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n694), .A2(new_n702), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n682), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT51), .B1(new_n774), .B2(new_n758), .ZN(new_n775));
  INV_X1    g574(.A(new_n762), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n650), .B(new_n771), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n767), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n704), .A2(new_n661), .A3(new_n706), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n777), .A2(new_n780), .A3(KEYINPUT110), .A4(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n777), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n763), .A2(KEYINPUT109), .A3(new_n650), .A4(new_n771), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n780), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n786), .A2(new_n791), .ZN(G1337gat));
  NAND2_X1  g591(.A1(new_n676), .A2(G99gat), .ZN(new_n793));
  NOR4_X1   g592(.A1(new_n765), .A2(new_n766), .A3(new_n767), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n763), .A2(new_n650), .A3(new_n674), .ZN(new_n795));
  INV_X1    g594(.A(G99gat), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1338gat));
  NAND4_X1  g598(.A1(new_n704), .A2(new_n427), .A3(new_n706), .A4(new_n778), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  INV_X1    g600(.A(new_n650), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n802), .A2(new_n428), .A3(G106gat), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT112), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n761), .B2(new_n762), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT53), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n800), .A2(KEYINPUT113), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n800), .A2(KEYINPUT113), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n807), .A2(G106gat), .A3(new_n808), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n805), .A2(KEYINPUT53), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(G1339gat));
  NAND3_X1  g610(.A1(new_n632), .A2(new_n633), .A3(new_n638), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n636), .A2(KEYINPUT54), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n634), .A2(new_n635), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n644), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT55), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n813), .A2(new_n818), .A3(new_n644), .A4(new_n815), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n649), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n622), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n608), .A2(new_n610), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n594), .B1(new_n601), .B2(new_n602), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n617), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n621), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n650), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n589), .B1(new_n821), .B2(new_n826), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n589), .A2(new_n820), .A3(new_n825), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT115), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n589), .A2(new_n820), .A3(new_n825), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n622), .A2(new_n820), .B1(new_n825), .B2(new_n650), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(new_n589), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n829), .A2(new_n520), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n734), .A2(new_n802), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n834), .B2(new_n836), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n736), .A2(new_n463), .A3(new_n738), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n466), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n261), .A3(new_n622), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n837), .A2(new_n838), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(new_n657), .A3(new_n463), .A4(new_n466), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n623), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n847), .B(new_n848), .ZN(G1340gat));
  NAND3_X1  g648(.A1(new_n842), .A2(new_n258), .A3(new_n650), .ZN(new_n850));
  OAI21_X1  g649(.A(G120gat), .B1(new_n845), .B2(new_n802), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(G1341gat));
  INV_X1    g651(.A(G127gat), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n845), .A2(new_n853), .A3(new_n520), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n842), .A2(new_n757), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n853), .ZN(G1342gat));
  OR2_X1    g655(.A1(new_n682), .A2(G134gat), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT56), .B1(new_n841), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n841), .A2(KEYINPUT56), .A3(new_n857), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n845), .B2(new_n682), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n859), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(G1343gat));
  NAND2_X1  g663(.A1(new_n834), .A2(new_n836), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT116), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n427), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n657), .A2(new_n463), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT119), .B1(new_n870), .B2(new_n676), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n318), .A2(new_n872), .A3(new_n657), .A4(new_n463), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n520), .B1(new_n827), .B2(new_n828), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n836), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n427), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n874), .B1(KEYINPUT57), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n869), .A2(new_n622), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G141gat), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n676), .A2(new_n428), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n840), .A2(new_n321), .A3(new_n622), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT58), .ZN(new_n884));
  XNOR2_X1  g683(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n879), .B2(G141gat), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  INV_X1    g686(.A(new_n839), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n866), .A2(new_n868), .A3(new_n888), .A4(new_n881), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(G141gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n887), .B1(new_n890), .B2(new_n622), .ZN(new_n891));
  NOR4_X1   g690(.A1(new_n889), .A2(KEYINPUT120), .A3(G141gat), .A4(new_n623), .ZN(new_n892));
  OAI211_X1 g691(.A(KEYINPUT122), .B(new_n886), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n882), .A2(KEYINPUT120), .ZN(new_n895));
  INV_X1    g694(.A(new_n889), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n896), .A2(new_n887), .A3(new_n321), .A4(new_n622), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT122), .B1(new_n898), .B2(new_n886), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n884), .B1(new_n894), .B2(new_n899), .ZN(G1344gat));
  NAND3_X1  g699(.A1(new_n869), .A2(new_n650), .A3(new_n878), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n902), .A3(G148gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n324), .B1(new_n889), .B2(new_n802), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n866), .A2(KEYINPUT57), .A3(new_n868), .A4(new_n427), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n877), .A2(new_n867), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n324), .B(new_n802), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n874), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g709(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n911));
  OAI211_X1 g710(.A(KEYINPUT124), .B(new_n903), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n906), .A2(new_n907), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n914), .A2(G148gat), .A3(new_n650), .A4(new_n909), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n911), .B1(new_n915), .B2(new_n904), .ZN(new_n916));
  INV_X1    g715(.A(new_n903), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n912), .A2(new_n918), .ZN(G1345gat));
  OAI21_X1  g718(.A(new_n328), .B1(new_n889), .B2(new_n520), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n869), .A2(G155gat), .A3(new_n878), .A4(new_n757), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(G1346gat));
  OAI21_X1  g721(.A(new_n329), .B1(new_n889), .B2(new_n682), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n869), .A2(G162gat), .A3(new_n878), .A4(new_n589), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(G1347gat));
  NAND3_X1  g724(.A1(new_n844), .A2(new_n428), .A3(new_n749), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n739), .A2(new_n661), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n623), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n466), .A2(new_n661), .ZN(new_n930));
  NOR4_X1   g729(.A1(new_n837), .A2(new_n838), .A3(new_n657), .A4(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n622), .A3(new_n220), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n929), .A2(new_n932), .ZN(G1348gat));
  AOI21_X1  g732(.A(G176gat), .B1(new_n931), .B2(new_n650), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n928), .A2(new_n802), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(G176gat), .ZN(G1349gat));
  NAND3_X1  g735(.A1(new_n931), .A2(new_n757), .A3(new_n241), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n926), .A2(new_n520), .A3(new_n927), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n280), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n928), .B2(new_n682), .ZN(new_n941));
  XOR2_X1   g740(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n931), .A2(new_n215), .A3(new_n589), .ZN(new_n945));
  OAI211_X1 g744(.A(G190gat), .B(new_n942), .C1(new_n928), .C2(new_n682), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G1351gat));
  NAND3_X1  g746(.A1(new_n739), .A2(new_n661), .A3(new_n318), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n914), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n623), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n837), .A2(new_n838), .A3(new_n657), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n661), .A3(new_n881), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(G197gat), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n952), .B1(new_n955), .B2(new_n622), .ZN(new_n956));
  NOR4_X1   g755(.A1(new_n954), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n623), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(G1352gat));
  INV_X1    g757(.A(new_n954), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n643), .A4(new_n650), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n914), .A2(new_n650), .A3(new_n949), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G204gat), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n953), .A2(new_n643), .A3(new_n661), .A4(new_n881), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT62), .B1(new_n964), .B2(new_n802), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n961), .A2(new_n963), .A3(new_n968), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n959), .A2(new_n385), .A3(new_n757), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n914), .A2(new_n757), .A3(new_n949), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  OAI21_X1  g774(.A(G218gat), .B1(new_n950), .B2(new_n682), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n386), .A3(new_n589), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1355gat));
endmodule


