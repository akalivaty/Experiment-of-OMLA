//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n582, new_n583, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n642, new_n643, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  XOR2_X1   g034(.A(G325), .B(KEYINPUT67), .Z(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  INV_X1    g037(.A(G113), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT69), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n471), .B(G125), .C1(new_n466), .C2(new_n467), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n465), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT70), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n471), .B1(new_n476), .B2(G125), .ZN(new_n477));
  INV_X1    g052(.A(new_n472), .ZN(new_n478));
  OAI22_X1  g053(.A1(new_n477), .A2(new_n478), .B1(new_n463), .B2(new_n464), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  OR2_X1    g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G137), .ZN(new_n486));
  INV_X1    g061(.A(G101), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n474), .A2(G2104), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G160));
  AND2_X1   g067(.A1(new_n476), .A2(KEYINPUT71), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n476), .A2(KEYINPUT71), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(new_n474), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G124), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n474), .B1(new_n493), .B2(new_n494), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G136), .ZN(new_n500));
  INV_X1    g075(.A(G100), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n501), .A2(new_n474), .A3(KEYINPUT72), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT72), .B1(new_n501), .B2(new_n474), .ZN(new_n503));
  OAI221_X1 g078(.A(G2104), .B1(G112), .B2(new_n474), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n497), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G162));
  AOI21_X1  g081(.A(KEYINPUT4), .B1(new_n485), .B2(G138), .ZN(new_n507));
  NAND2_X1  g082(.A1(G126), .A2(G2105), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT4), .A2(G138), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(G2105), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n476), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G114), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G2105), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n507), .A2(new_n517), .ZN(G164));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  OR2_X1    g099(.A1(KEYINPUT73), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT73), .A2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT74), .B1(new_n530), .B2(KEYINPUT6), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT6), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(new_n533), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n525), .A2(KEYINPUT6), .A3(new_n526), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n535), .A2(new_n536), .A3(G50), .A4(G543), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT75), .B(G88), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n535), .A2(new_n536), .A3(new_n523), .A4(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n540), .B1(new_n537), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n529), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT77), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g120(.A(KEYINPUT77), .B(new_n529), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G166));
  NAND4_X1  g122(.A1(new_n535), .A2(new_n536), .A3(G51), .A4(G543), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n535), .A2(new_n536), .A3(G89), .A4(new_n523), .ZN(new_n549));
  AND2_X1   g124(.A1(G63), .A2(G651), .ZN(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT7), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n553), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n523), .A2(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n548), .A2(new_n549), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT78), .A4(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(G168));
  NAND3_X1  g135(.A1(new_n535), .A2(new_n536), .A3(G543), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G52), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n528), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n535), .A2(new_n536), .A3(new_n523), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G90), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(G301));
  INV_X1    g143(.A(G301), .ZN(G171));
  AOI22_X1  g144(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(new_n528), .ZN(new_n571));
  XOR2_X1   g146(.A(KEYINPUT79), .B(G43), .Z(new_n572));
  NAND2_X1  g147(.A1(new_n562), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n566), .A2(G81), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n574), .B1(new_n573), .B2(new_n575), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n571), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G860), .ZN(G153));
  NAND4_X1  g155(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g156(.A1(G1), .A2(G3), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT8), .ZN(new_n583));
  NAND4_X1  g158(.A1(G319), .A2(G483), .A3(G661), .A4(new_n583), .ZN(G188));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n523), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n521), .A2(KEYINPUT82), .A3(new_n522), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(G78), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT81), .B(KEYINPUT9), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n562), .A2(G53), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n566), .A2(G91), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT9), .ZN(new_n595));
  INV_X1    g170(.A(G53), .ZN(new_n596));
  OAI211_X1 g171(.A(KEYINPUT81), .B(new_n595), .C1(new_n561), .C2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n591), .A2(new_n593), .A3(new_n594), .A4(new_n597), .ZN(G299));
  INV_X1    g173(.A(G168), .ZN(G286));
  INV_X1    g174(.A(G166), .ZN(G303));
  NAND2_X1  g175(.A1(new_n562), .A2(G49), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n566), .A2(G87), .ZN(new_n602));
  OAI21_X1  g177(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(G288));
  INV_X1    g179(.A(G86), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n521), .B2(new_n522), .ZN(new_n606));
  AND2_X1   g181(.A1(G48), .A2(G543), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n536), .B(new_n535), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G61), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n521), .B2(new_n522), .ZN(new_n610));
  AND2_X1   g185(.A1(G73), .A2(G543), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n527), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(G305));
  NAND2_X1  g188(.A1(new_n562), .A2(G47), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(new_n528), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n566), .A2(G85), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(G290));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(G301), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n566), .A2(G92), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT10), .Z(new_n622));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  AND2_X1   g199(.A1(new_n587), .A2(new_n588), .ZN(new_n625));
  INV_X1    g200(.A(G66), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n626), .B1(new_n587), .B2(new_n588), .ZN(new_n628));
  INV_X1    g203(.A(new_n624), .ZN(new_n629));
  OAI21_X1  g204(.A(KEYINPUT83), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n627), .A2(G651), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n562), .A2(G54), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n631), .A2(KEYINPUT84), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(KEYINPUT84), .B1(new_n631), .B2(new_n632), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n622), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT85), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT85), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n637), .B(new_n622), .C1(new_n633), .C2(new_n634), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n620), .B1(new_n639), .B2(new_n619), .ZN(G284));
  AOI21_X1  g215(.A(new_n620), .B1(new_n639), .B2(new_n619), .ZN(G321));
  NOR2_X1   g216(.A1(G286), .A2(new_n619), .ZN(new_n642));
  XNOR2_X1  g217(.A(G299), .B(KEYINPUT86), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(new_n619), .ZN(G297));
  AOI21_X1  g219(.A(new_n642), .B1(new_n643), .B2(new_n619), .ZN(G280));
  INV_X1    g220(.A(G559), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n639), .B1(new_n646), .B2(G860), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT87), .ZN(G148));
  OAI21_X1  g223(.A(KEYINPUT88), .B1(new_n579), .B2(G868), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n639), .A2(new_n646), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G868), .ZN(new_n651));
  MUX2_X1   g226(.A(KEYINPUT88), .B(new_n649), .S(new_n651), .Z(G323));
  XNOR2_X1  g227(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g228(.A1(new_n468), .A2(new_n488), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT13), .ZN(new_n657));
  AOI22_X1  g232(.A1(new_n656), .A2(new_n657), .B1(KEYINPUT89), .B2(G2100), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n656), .ZN(new_n659));
  OR3_X1    g234(.A1(new_n659), .A2(KEYINPUT89), .A3(G2100), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n496), .A2(G123), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n499), .A2(G135), .ZN(new_n662));
  OR2_X1    g237(.A1(G99), .A2(G2105), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n663), .B(G2104), .C1(G111), .C2(new_n474), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(G2096), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n659), .B1(KEYINPUT89), .B2(G2100), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(G2096), .ZN(new_n668));
  NAND4_X1  g243(.A1(new_n660), .A2(new_n666), .A3(new_n667), .A4(new_n668), .ZN(G156));
  XNOR2_X1  g244(.A(G2427), .B(G2438), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2430), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT15), .B(G2435), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(KEYINPUT14), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2451), .B(G2454), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT16), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2443), .B(G2446), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1341), .B(G1348), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT90), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n685), .A2(G14), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n684), .A2(new_n686), .ZN(G401));
  XNOR2_X1  g262(.A(G2072), .B(G2078), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT17), .Z(new_n689));
  XOR2_X1   g264(.A(G2084), .B(G2090), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT91), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2067), .B(G2678), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n689), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT92), .Z(new_n695));
  NAND3_X1  g270(.A1(new_n691), .A2(new_n688), .A3(new_n692), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT18), .Z(new_n697));
  NOR2_X1   g272(.A1(new_n689), .A2(new_n693), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n688), .A2(new_n692), .ZN(new_n699));
  OR3_X1    g274(.A1(new_n698), .A2(new_n691), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n695), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G2096), .B(G2100), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(G227));
  XNOR2_X1  g278(.A(G1956), .B(G2474), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1961), .B(G1966), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1971), .B(G1976), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT19), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n705), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n706), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n708), .A2(new_n709), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT20), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(G1991), .B(G1996), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(G1981), .B(G1986), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(G229));
  NAND3_X1  g298(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT25), .Z(new_n725));
  AOI22_X1  g300(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n726));
  INV_X1    g301(.A(G139), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n725), .B1(new_n474), .B2(new_n726), .C1(new_n498), .C2(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G33), .B(new_n728), .S(G29), .Z(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G2072), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT98), .Z(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G26), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT28), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n496), .A2(G128), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n499), .A2(G140), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n474), .A2(G116), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n739), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2067), .ZN(new_n741));
  NOR2_X1   g316(.A1(G27), .A2(G29), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G164), .B2(G29), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2078), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT31), .B(G11), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT101), .ZN(new_n746));
  INV_X1    g321(.A(G28), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n747), .B2(KEYINPUT30), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n665), .B2(new_n732), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n744), .B(new_n751), .C1(G2072), .C2(new_n729), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n731), .A2(new_n741), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n732), .A2(G32), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT26), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G105), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n488), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n496), .B2(G129), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n499), .A2(G141), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n754), .B1(new_n765), .B2(new_n732), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G16), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n732), .A2(G35), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G162), .B2(new_n732), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT29), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n768), .B(new_n773), .C1(new_n776), .C2(G2090), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G21), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G168), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1966), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT95), .B(G16), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G19), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n579), .B2(new_n782), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1341), .ZN(new_n785));
  OR4_X1    g360(.A1(new_n753), .A2(new_n777), .A3(new_n780), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n769), .A2(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n639), .B2(new_n769), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(G1348), .ZN(new_n789));
  INV_X1    g364(.A(G2084), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G34), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(new_n732), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n491), .B2(new_n732), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n776), .A2(G2090), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n790), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT100), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n781), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT23), .ZN(new_n799));
  INV_X1    g374(.A(G299), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n769), .ZN(new_n801));
  INV_X1    g376(.A(G1956), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n795), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n786), .A2(new_n789), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n788), .A2(G1348), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n808));
  MUX2_X1   g383(.A(G6), .B(G305), .S(G16), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT32), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1981), .ZN(new_n811));
  NOR2_X1   g386(.A1(G16), .A2(G23), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT96), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G288), .B2(new_n769), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT33), .B(G1976), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(G1971), .ZN(new_n818));
  NAND2_X1  g393(.A1(G303), .A2(new_n782), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n781), .A2(G22), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n819), .A2(new_n818), .A3(new_n820), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n817), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  NOR2_X1   g400(.A1(G25), .A2(G29), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n827));
  INV_X1    g402(.A(G107), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(G2105), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n496), .B2(G119), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n499), .A2(new_n831), .A3(G131), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n499), .B2(G131), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n826), .B1(new_n835), .B2(G29), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT35), .B(G1991), .Z(new_n837));
  XOR2_X1   g412(.A(new_n836), .B(new_n837), .Z(new_n838));
  NOR2_X1   g413(.A1(new_n782), .A2(G24), .ZN(new_n839));
  INV_X1    g414(.A(G290), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(new_n782), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1986), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(KEYINPUT97), .B1(new_n825), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n843), .B(new_n846), .C1(KEYINPUT34), .C2(new_n824), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n808), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n808), .A3(new_n849), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n807), .B1(new_n851), .B2(new_n852), .ZN(G311));
  INV_X1    g428(.A(new_n852), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n806), .B(new_n805), .C1(new_n854), .C2(new_n850), .ZN(G150));
  AOI22_X1  g430(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n528), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT102), .ZN(new_n858));
  AOI22_X1  g433(.A1(G55), .A2(new_n562), .B1(new_n566), .B2(G93), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT103), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n862), .A3(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n639), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT38), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n578), .A3(new_n863), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n579), .A2(new_n860), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n868), .B(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  INV_X1    g448(.A(G860), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n872), .B2(KEYINPUT39), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n866), .B1(new_n873), .B2(new_n875), .ZN(G145));
  XNOR2_X1  g451(.A(new_n491), .B(KEYINPUT104), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n665), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n834), .B(new_n656), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n764), .B(new_n728), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G164), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n739), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n496), .A2(G130), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n499), .A2(G142), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n474), .A2(G118), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n885), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n883), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n880), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n883), .B(new_n891), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n879), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g473(.A1(new_n864), .A2(new_n619), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n900));
  INV_X1    g475(.A(new_n871), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n650), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n639), .A2(new_n646), .A3(new_n871), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n635), .B(G299), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n635), .B(new_n800), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n903), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n871), .B1(new_n639), .B2(new_n646), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n904), .A2(KEYINPUT105), .A3(new_n908), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(G303), .A2(G290), .ZN(new_n919));
  NOR2_X1   g494(.A1(G166), .A2(new_n840), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(G288), .B(KEYINPUT106), .Z(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(G305), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n923), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n619), .B1(new_n918), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n927), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n926), .B(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n931), .A2(new_n911), .A3(new_n916), .A4(new_n917), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n900), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  OAI22_X1  g509(.A1(new_n914), .A2(new_n915), .B1(new_n904), .B2(new_n910), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT105), .B1(new_n904), .B2(new_n908), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n928), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND4_X1   g512(.A1(new_n934), .A2(new_n937), .A3(new_n932), .A4(G868), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n933), .A2(new_n938), .ZN(G295));
  NOR2_X1   g514(.A1(new_n933), .A2(new_n938), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  NOR2_X1   g516(.A1(G286), .A2(KEYINPUT109), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G171), .B1(G286), .B2(KEYINPUT109), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n869), .A2(new_n870), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n869), .B2(new_n870), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n948), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n942), .A3(new_n946), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n908), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n907), .A2(new_n909), .A3(new_n951), .A4(new_n949), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n955), .B2(new_n926), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n953), .A2(new_n954), .A3(new_n925), .A4(new_n924), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n941), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n958), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(KEYINPUT44), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n961), .A2(new_n965), .ZN(G397));
  INV_X1    g541(.A(G2067), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n739), .B(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n765), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n764), .A2(G1996), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(KEYINPUT110), .B(G40), .Z(new_n973));
  NOR2_X1   g548(.A1(new_n489), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n475), .A2(new_n481), .A3(new_n974), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n476), .A2(new_n510), .B1(new_n513), .B2(new_n515), .ZN(new_n976));
  OAI211_X1 g551(.A(G138), .B(new_n474), .C1(new_n466), .C2(new_n467), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT4), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n975), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n972), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n972), .A2(KEYINPUT111), .A3(new_n981), .ZN(new_n985));
  INV_X1    g560(.A(new_n981), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n834), .B(new_n837), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n984), .B(new_n985), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(G290), .B(G1986), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n981), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n980), .B(KEYINPUT45), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n975), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n443), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n475), .A2(new_n481), .A3(new_n974), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n507), .B2(new_n517), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n980), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n993), .A2(new_n994), .B1(new_n772), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n994), .A2(G2078), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n992), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G171), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n997), .B(KEYINPUT45), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1966), .B1(new_n995), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n998), .A2(new_n1000), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n975), .A2(new_n1010), .A3(G2084), .ZN(new_n1011));
  OAI21_X1  g586(.A(G8), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n558), .A2(G8), .A3(new_n559), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT122), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1013), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT51), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n995), .A2(new_n1001), .A3(new_n790), .ZN(new_n1021));
  INV_X1    g596(.A(G1966), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n975), .B2(new_n991), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1016), .B1(new_n1024), .B2(G8), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1018), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT62), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1007), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n545), .A2(G8), .A3(new_n546), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(KEYINPUT113), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n545), .A2(G8), .A3(new_n546), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT112), .B(G1971), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n995), .B2(new_n1008), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n975), .A2(new_n1010), .A3(G2090), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G2090), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n995), .A2(new_n1001), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1036), .B1(new_n975), .B2(new_n991), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1032), .A2(new_n1045), .A3(G8), .A4(new_n1034), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n475), .A2(new_n481), .A3(new_n980), .A4(new_n974), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  INV_X1    g626(.A(G1981), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n608), .B2(new_n612), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n608), .A2(new_n1052), .A3(new_n612), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n1055), .B(new_n1052), .C1(new_n608), .C2(new_n612), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT115), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1051), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1061), .B2(new_n1051), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1057), .A2(new_n1059), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1050), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n601), .A2(new_n602), .A3(G1976), .A4(new_n603), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1049), .A2(G8), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT52), .ZN(new_n1070));
  INV_X1    g645(.A(G1976), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(G288), .B2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1072), .A2(new_n1049), .A3(G8), .A4(new_n1068), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1048), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1056), .A2(new_n1055), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n1053), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(new_n1058), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT116), .B1(new_n1079), .B2(KEYINPUT115), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1065), .B1(new_n1080), .B2(new_n1051), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT117), .B(new_n1076), .C1(new_n1081), .C2(new_n1050), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1047), .B1(new_n1075), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1018), .B(KEYINPUT62), .C1(new_n1020), .C2(new_n1025), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(KEYINPUT51), .A3(new_n1019), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(KEYINPUT124), .A3(KEYINPUT62), .A4(new_n1018), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1028), .A2(new_n1083), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1046), .A2(new_n1067), .A3(new_n1074), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1050), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1081), .ZN(new_n1093));
  OR2_X1    g668(.A1(G288), .A2(G1976), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1056), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1091), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1012), .A2(G286), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT63), .B1(new_n1083), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(KEYINPUT63), .ZN(new_n1099));
  NOR4_X1   g674(.A1(new_n1047), .A2(new_n1099), .A3(new_n1067), .A4(new_n1074), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1090), .B(new_n1096), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1026), .ZN(new_n1102));
  XNOR2_X1  g677(.A(G301), .B(KEYINPUT54), .ZN(new_n1103));
  AND4_X1   g678(.A1(G40), .A2(new_n1008), .A3(new_n490), .A4(new_n1004), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n474), .B1(new_n479), .B2(KEYINPUT123), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(KEYINPUT123), .B2(new_n479), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1103), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1006), .A2(new_n1103), .B1(new_n1003), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1083), .A2(new_n1102), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1002), .ZN(new_n1110));
  OAI22_X1  g685(.A1(new_n1110), .A2(G1348), .B1(G2067), .B2(new_n1049), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n639), .A2(KEYINPUT60), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n636), .B(new_n638), .C1(new_n1111), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(new_n442), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n802), .A2(new_n1002), .B1(new_n992), .B2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1122));
  NAND2_X1  g697(.A1(G299), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n800), .A2(KEYINPUT57), .ZN(new_n1126));
  NAND3_X1  g701(.A1(G299), .A2(KEYINPUT119), .A3(new_n1122), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1121), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1121), .A2(new_n1128), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1118), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  NAND3_X1  g708(.A1(new_n1049), .A2(KEYINPUT121), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n995), .A2(new_n1008), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1135), .B2(G1996), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT121), .B1(new_n1049), .B2(new_n1133), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n579), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT59), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1131), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n1129), .A3(KEYINPUT61), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1117), .A2(new_n1132), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n639), .A2(new_n1111), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1129), .B1(new_n1143), .B2(new_n1131), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1109), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n990), .B1(new_n1101), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n835), .A2(new_n837), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n984), .A2(new_n985), .A3(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n739), .A2(G2067), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1147), .B1(new_n1152), .B2(new_n981), .ZN(new_n1153));
  AOI211_X1 g728(.A(KEYINPUT125), .B(new_n986), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n968), .A2(new_n765), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT46), .B1(new_n986), .B2(G1996), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT46), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n981), .A2(new_n1157), .A3(new_n969), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1155), .A2(new_n981), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT47), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n986), .A2(G1986), .A3(G290), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT48), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1161), .B1(new_n988), .B2(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1153), .A2(new_n1154), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1146), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1146), .A2(new_n1165), .A3(KEYINPUT126), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g745(.A(new_n461), .ZN(new_n1172));
  OR2_X1    g746(.A1(G227), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g747(.A(new_n1173), .B1(new_n684), .B2(new_n686), .ZN(new_n1174));
  OR2_X1    g748(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1175));
  AOI21_X1  g749(.A(G229), .B1(new_n1174), .B2(KEYINPUT127), .ZN(new_n1176));
  NAND3_X1  g750(.A1(new_n897), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g751(.A(new_n1177), .B1(new_n963), .B2(new_n964), .ZN(G308));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1179), .B1(new_n960), .B2(new_n959), .ZN(G225));
endmodule


