//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G110), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(new_n192), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT24), .B(G110), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT71), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(new_n201), .A3(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT72), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT72), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n210), .A2(new_n207), .A3(new_n201), .A4(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT71), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n202), .A2(new_n204), .A3(new_n213), .A4(KEYINPUT16), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n206), .A2(new_n212), .A3(G146), .A4(new_n214), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n200), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G137), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(KEYINPUT74), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n224), .B(KEYINPUT75), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n222), .B(new_n225), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT73), .B(G110), .Z(new_n227));
  OR2_X1    g041(.A1(new_n195), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n198), .A2(new_n199), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n202), .A2(new_n204), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n228), .A2(new_n229), .B1(new_n216), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n218), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n220), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n225), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n222), .B(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n232), .A2(new_n218), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(new_n219), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n188), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G217), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(new_n187), .B2(G234), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n239), .B2(new_n240), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n234), .A2(new_n238), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT76), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n234), .A2(new_n238), .A3(KEYINPUT76), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n244), .A2(G902), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n242), .A2(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  NOR2_X1   g069(.A1(G237), .A2(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G210), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n255), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n258), .B(new_n259), .Z(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n216), .A2(G143), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n193), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n263), .A2(KEYINPUT1), .A3(G146), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT11), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(G137), .ZN(new_n274));
  INV_X1    g088(.A(G137), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT11), .A3(G134), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(G137), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n274), .A2(new_n276), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n273), .A2(G137), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n275), .A2(G134), .ZN(new_n281));
  OAI21_X1  g095(.A(G131), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n279), .A2(new_n282), .A3(KEYINPUT67), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT67), .B1(new_n279), .B2(new_n282), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n271), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n190), .B2(G116), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT66), .A3(G119), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n190), .A2(G116), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(KEYINPUT2), .A2(G113), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT65), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT2), .A3(G113), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT2), .ZN(new_n298));
  INV_X1    g112(.A(G113), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n287), .A2(new_n289), .B1(G116), .B2(new_n190), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n300), .A3(new_n297), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n274), .A2(new_n276), .A3(new_n278), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G131), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n279), .ZN(new_n308));
  NOR2_X1   g122(.A1(KEYINPUT0), .A2(G128), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT0), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(new_n193), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n265), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n262), .B(new_n264), .C1(new_n310), .C2(new_n193), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n285), .A2(new_n305), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT64), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n279), .A2(new_n282), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n279), .B2(new_n282), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n271), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n305), .B1(new_n321), .B2(new_n315), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT28), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n261), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n302), .A2(new_n304), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT30), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n321), .A2(new_n328), .A3(new_n315), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n285), .B2(new_n315), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n261), .A3(new_n316), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT31), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n331), .A2(KEYINPUT31), .A3(new_n261), .A4(new_n316), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n326), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(G472), .A2(G902), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT32), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n326), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n268), .A2(new_n262), .A3(new_n264), .ZN(new_n341));
  AOI21_X1  g155(.A(G128), .B1(new_n262), .B2(new_n264), .ZN(new_n342));
  INV_X1    g156(.A(new_n270), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n279), .A2(new_n282), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n279), .A2(new_n282), .A3(KEYINPUT67), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n308), .A2(new_n314), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT30), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n321), .A2(new_n328), .A3(new_n315), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n317), .B1(new_n353), .B2(new_n327), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT31), .B1(new_n354), .B2(new_n261), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n305), .B1(new_n351), .B2(new_n352), .ZN(new_n356));
  NOR4_X1   g170(.A1(new_n356), .A2(new_n333), .A3(new_n317), .A4(new_n260), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n340), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT32), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n337), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n339), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n260), .B1(new_n356), .B2(new_n317), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n323), .A2(new_n325), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n260), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n305), .B1(new_n285), .B2(new_n315), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n316), .B1(new_n366), .B2(KEYINPUT69), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT69), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n285), .A2(new_n368), .A3(new_n305), .A4(new_n315), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n325), .B1(new_n370), .B2(new_n324), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n261), .A2(KEYINPUT29), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n365), .B(new_n187), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G472), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n254), .B1(new_n361), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n230), .A2(KEYINPUT88), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT88), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n202), .A2(new_n204), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(G146), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT89), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n231), .A2(new_n216), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n376), .A2(KEYINPUT89), .A3(G146), .A4(new_n378), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT90), .ZN(new_n385));
  INV_X1    g199(.A(G237), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n223), .A3(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n263), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n256), .A2(G143), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT18), .A2(G131), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n385), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AND4_X1   g207(.A1(G143), .A2(new_n386), .A3(new_n223), .A4(G214), .ZN(new_n394));
  AOI21_X1  g208(.A(G143), .B1(new_n256), .B2(G214), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT90), .A3(new_n391), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n391), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT86), .B1(new_n394), .B2(new_n395), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n388), .A2(new_n400), .A3(new_n389), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n402), .A2(new_n404), .A3(new_n399), .A4(new_n392), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n384), .B(new_n398), .C1(new_n403), .C2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G113), .B(G122), .ZN(new_n408));
  INV_X1    g222(.A(G104), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n396), .A2(new_n277), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n390), .A2(G131), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n390), .A2(KEYINPUT17), .A3(G131), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n414), .A2(new_n217), .A3(new_n218), .A4(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n410), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT92), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n376), .A2(KEYINPUT19), .A3(new_n378), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n420));
  OR3_X1    g234(.A1(new_n230), .A2(new_n420), .A3(KEYINPUT19), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n420), .B1(new_n230), .B2(KEYINPUT19), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n419), .A2(new_n421), .A3(new_n216), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n411), .A2(new_n412), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n218), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n402), .A2(new_n404), .A3(new_n392), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT87), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n427), .A2(new_n405), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n379), .A2(new_n380), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n383), .A2(new_n382), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n398), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n418), .B(new_n425), .C1(new_n428), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n410), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n418), .B1(new_n407), .B2(new_n425), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n417), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n437));
  NOR2_X1   g251(.A1(G475), .A2(G902), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT93), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT93), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n436), .A2(new_n441), .A3(new_n437), .A4(new_n438), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n407), .A2(new_n410), .A3(new_n416), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n383), .A2(new_n382), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n444), .A2(new_n381), .B1(new_n393), .B2(new_n397), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n427), .A2(new_n405), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n424), .A2(new_n218), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n445), .A2(new_n446), .B1(new_n447), .B2(new_n423), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n410), .B1(new_n448), .B2(new_n418), .ZN(new_n449));
  INV_X1    g263(.A(new_n435), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n443), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n438), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT20), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n440), .A2(new_n442), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G902), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n410), .B1(new_n407), .B2(new_n416), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n455), .B1(new_n443), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT94), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n459), .B(new_n455), .C1(new_n443), .C2(new_n456), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(G475), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT97), .ZN(new_n462));
  INV_X1    g276(.A(G107), .ZN(new_n463));
  INV_X1    g277(.A(G122), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G116), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n463), .B1(new_n465), .B2(KEYINPUT14), .ZN(new_n466));
  XNOR2_X1  g280(.A(G116), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n263), .A2(G128), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n193), .A2(G143), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT96), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT96), .ZN(new_n473));
  AOI21_X1  g287(.A(G134), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n475), .A2(new_n273), .A3(new_n471), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n468), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n288), .A2(G122), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n465), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(new_n463), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n467), .A2(G107), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT95), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n273), .B1(new_n475), .B2(new_n471), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT13), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n193), .B2(G143), .ZN(new_n485));
  INV_X1    g299(.A(new_n469), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n469), .A2(new_n484), .ZN(new_n488));
  OAI21_X1  g302(.A(G134), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n479), .A2(new_n463), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n467), .A2(G107), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n482), .A2(new_n483), .A3(new_n489), .A4(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT9), .B(G234), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n495), .A2(new_n243), .A3(G953), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n477), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n477), .B2(new_n494), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n462), .B(new_n187), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G478), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(KEYINPUT15), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n477), .A2(new_n494), .ZN(new_n503));
  INV_X1    g317(.A(new_n496), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n477), .A2(new_n494), .A3(new_n496), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n462), .B1(new_n507), .B2(new_n187), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  AOI211_X1 g323(.A(new_n462), .B(new_n501), .C1(new_n507), .C2(new_n187), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n223), .A2(G952), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(G234), .B2(G237), .ZN(new_n513));
  AOI211_X1 g327(.A(new_n223), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT21), .B(G898), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n454), .A2(new_n461), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G214), .B1(G237), .B2(G902), .ZN(new_n519));
  XNOR2_X1  g333(.A(G110), .B(G122), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(KEYINPUT78), .A2(G101), .ZN(new_n522));
  NOR2_X1   g336(.A1(KEYINPUT78), .A2(G101), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n409), .A2(G107), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n463), .A2(KEYINPUT3), .A3(G104), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT3), .B1(new_n463), .B2(G104), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n524), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G101), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT3), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n409), .B2(G107), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n463), .A2(KEYINPUT3), .A3(G104), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n531), .A2(new_n532), .B1(new_n409), .B2(G107), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n528), .B(KEYINPUT4), .C1(new_n529), .C2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT82), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(G101), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n327), .A2(new_n534), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n409), .A2(KEYINPUT80), .A3(G107), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT80), .B1(new_n409), .B2(G107), .ZN(new_n541));
  OAI22_X1  g355(.A1(new_n540), .A2(new_n541), .B1(new_n409), .B2(G107), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n542), .A2(G101), .B1(new_n533), .B2(new_n524), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n303), .A2(KEYINPUT5), .ZN(new_n544));
  OAI21_X1  g358(.A(G113), .B1(new_n291), .B2(KEYINPUT5), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n543), .B(new_n304), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n539), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n533), .A2(new_n529), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n302), .A2(new_n304), .B1(new_n548), .B2(new_n537), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n535), .B1(new_n549), .B2(new_n534), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n521), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n327), .A2(new_n534), .A3(new_n538), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT82), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n553), .A2(new_n539), .A3(new_n546), .A4(new_n520), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(KEYINPUT6), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT6), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n556), .B(new_n521), .C1(new_n547), .C2(new_n550), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n311), .A2(new_n309), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n313), .B(G125), .C1(new_n558), .C2(new_n267), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT83), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n312), .A2(KEYINPUT83), .A3(G125), .A4(new_n313), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n342), .A2(new_n343), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n203), .A3(new_n269), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G224), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G953), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n565), .B(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n555), .A2(new_n557), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT84), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n561), .A2(new_n570), .A3(new_n562), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT7), .B1(new_n566), .B2(G953), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n565), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n565), .B1(new_n572), .B2(new_n571), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n520), .B(KEYINPUT8), .Z(new_n575));
  INV_X1    g389(.A(new_n524), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n409), .A2(G107), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT80), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n463), .B2(G104), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n409), .A2(KEYINPUT80), .A3(G107), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI22_X1  g395(.A1(new_n536), .A2(new_n576), .B1(new_n581), .B2(new_n529), .ZN(new_n582));
  INV_X1    g396(.A(new_n304), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n545), .B1(new_n303), .B2(KEYINPUT5), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n575), .B1(new_n546), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n573), .A2(new_n574), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n587), .B2(new_n554), .ZN(new_n588));
  OAI21_X1  g402(.A(G210), .B1(G237), .B2(G902), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT85), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n569), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n569), .B2(new_n588), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n519), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G221), .B1(new_n495), .B2(G902), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT77), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G469), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n538), .A2(new_n314), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT10), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n563), .B2(new_n269), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n599), .A2(new_n534), .B1(new_n543), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n269), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n268), .A2(new_n262), .A3(new_n264), .A4(KEYINPUT81), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n563), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT10), .B1(new_n606), .B2(new_n543), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n308), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n602), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n542), .A2(G101), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n271), .A2(new_n611), .A3(KEYINPUT10), .A4(new_n528), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT4), .B1(new_n533), .B2(new_n529), .ZN(new_n613));
  INV_X1    g427(.A(new_n528), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n538), .A2(new_n314), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n308), .B1(new_n617), .B2(new_n607), .ZN(new_n618));
  XNOR2_X1  g432(.A(G110), .B(G140), .ZN(new_n619));
  INV_X1    g433(.A(G227), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(G953), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n619), .B(new_n621), .Z(new_n622));
  NAND3_X1  g436(.A1(new_n610), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n266), .A2(new_n270), .A3(new_n605), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT81), .B1(new_n267), .B2(new_n268), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n528), .B(new_n611), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n582), .A2(new_n344), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n308), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT12), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n628), .A2(KEYINPUT12), .A3(new_n308), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n617), .A2(new_n607), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n631), .A2(new_n632), .B1(new_n633), .B2(new_n609), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n623), .B1(new_n634), .B2(new_n622), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n598), .B1(new_n635), .B2(new_n455), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n610), .A2(new_n618), .ZN(new_n637));
  INV_X1    g451(.A(new_n622), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n632), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT12), .B1(new_n628), .B2(new_n308), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n610), .B(new_n622), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  AOI211_X1 g456(.A(G469), .B(new_n188), .C1(new_n639), .C2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n597), .B1(new_n636), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n594), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n375), .A2(new_n518), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n576), .ZN(G3));
  INV_X1    g461(.A(new_n516), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n648), .B(new_n519), .C1(new_n592), .C2(new_n593), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n454), .A2(new_n461), .ZN(new_n650));
  AOI21_X1  g464(.A(G478), .B1(new_n507), .B2(new_n187), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT98), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n505), .A2(new_n506), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n652), .A2(KEYINPUT98), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n188), .A2(new_n500), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n651), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n658), .B1(new_n454), .B2(new_n461), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n649), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n253), .B(new_n597), .C1(new_n636), .C2(new_n643), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n336), .B2(new_n188), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n358), .A2(new_n337), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT100), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(new_n649), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n437), .B1(new_n436), .B2(new_n438), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n461), .B(new_n511), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n675), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT101), .B1(new_n649), .B2(new_n678), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n670), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT102), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT35), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G107), .ZN(G9));
  INV_X1    g501(.A(KEYINPUT36), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n220), .A2(new_n236), .A3(new_n688), .A4(new_n233), .ZN(new_n689));
  OAI22_X1  g503(.A1(new_n237), .A2(new_n219), .B1(new_n226), .B2(KEYINPUT36), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n252), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT103), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n689), .A2(new_n690), .A3(new_n693), .A4(new_n252), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n246), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n695), .B1(new_n696), .B2(new_n241), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n669), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n518), .A2(new_n699), .A3(new_n645), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT37), .B(G110), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G12));
  AOI21_X1  g516(.A(new_n698), .B1(new_n361), .B2(new_n374), .ZN(new_n703));
  INV_X1    g517(.A(G900), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n513), .B1(new_n514), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n678), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n645), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  XOR2_X1   g522(.A(new_n705), .B(KEYINPUT39), .Z(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  OR3_X1    g524(.A1(new_n644), .A2(KEYINPUT40), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT40), .B1(new_n644), .B2(new_n710), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n519), .A2(new_n711), .A3(new_n698), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n569), .A2(new_n588), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n590), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n569), .A2(new_n588), .A3(new_n591), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT38), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n332), .B1(new_n370), .B2(new_n261), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n455), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G472), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n361), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n511), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n454), .B2(new_n461), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n713), .A2(new_n718), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT104), .B(G143), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G45));
  INV_X1    g541(.A(new_n705), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n703), .A2(new_n645), .A3(new_n663), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  AOI22_X1  g544(.A1(new_n339), .A2(new_n360), .B1(G472), .B2(new_n373), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n639), .A2(new_n642), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n187), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G469), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n598), .A3(new_n187), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n597), .A3(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n731), .A2(new_n254), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n664), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n675), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND2_X1  g556(.A1(new_n683), .A2(new_n737), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT105), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n683), .A2(new_n745), .A3(new_n737), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR2_X1   g562(.A1(new_n594), .A2(new_n736), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n703), .A2(new_n518), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n703), .A2(new_n518), .A3(KEYINPUT106), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G119), .ZN(G21));
  AOI21_X1  g569(.A(new_n324), .B1(new_n367), .B2(new_n369), .ZN(new_n756));
  INV_X1    g570(.A(new_n325), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n260), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n355), .B2(new_n357), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n337), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n667), .A2(new_n253), .A3(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n761), .A2(new_n516), .A3(new_n736), .ZN(new_n762));
  INV_X1    g576(.A(new_n594), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n724), .A2(KEYINPUT107), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT107), .B1(new_n724), .B2(new_n763), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT108), .B(G122), .Z(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G24));
  NAND3_X1  g583(.A1(new_n667), .A2(new_n697), .A3(new_n760), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n667), .A2(new_n760), .A3(new_n697), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n705), .B(new_n658), .C1(new_n454), .C2(new_n461), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(new_n749), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G125), .ZN(G27));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n336), .A2(KEYINPUT32), .A3(new_n338), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n359), .B1(new_n358), .B2(new_n337), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n374), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n715), .A2(new_n519), .A3(new_n716), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n644), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n783), .A3(new_n253), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n650), .A2(new_n659), .A3(new_n728), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n778), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n775), .A2(KEYINPUT42), .A3(new_n375), .A4(new_n783), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G131), .ZN(G33));
  NAND3_X1  g603(.A1(new_n375), .A2(new_n706), .A3(new_n783), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  OR3_X1    g605(.A1(new_n650), .A2(KEYINPUT43), .A3(new_n658), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT43), .B1(new_n650), .B2(new_n658), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n669), .A3(new_n697), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n635), .B(KEYINPUT45), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(G469), .ZN(new_n798));
  NAND2_X1  g612(.A1(G469), .A2(G902), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n801), .B(G469), .C1(new_n797), .C2(G902), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n735), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n597), .A3(new_n709), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n796), .A2(new_n782), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n794), .A2(new_n795), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G137), .ZN(G39));
  NOR4_X1   g622(.A1(new_n785), .A2(new_n253), .A3(new_n781), .A4(new_n782), .ZN(new_n809));
  NAND2_X1  g623(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n803), .A2(new_n597), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI211_X1 g627(.A(KEYINPUT110), .B(KEYINPUT47), .C1(new_n803), .C2(new_n597), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n809), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(KEYINPUT111), .B(new_n809), .C1(new_n813), .C2(new_n814), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  AND2_X1   g634(.A1(new_n734), .A2(new_n735), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT49), .Z(new_n822));
  NAND3_X1  g636(.A1(new_n253), .A2(new_n519), .A3(new_n597), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n822), .A2(new_n718), .A3(new_n823), .ZN(new_n824));
  OR4_X1    g638(.A1(new_n650), .A2(new_n824), .A3(new_n658), .A4(new_n722), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n645), .B(new_n703), .C1(new_n775), .C2(new_n706), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n776), .ZN(new_n829));
  INV_X1    g643(.A(new_n644), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n697), .A2(new_n705), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n722), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n650), .A2(new_n511), .A3(new_n763), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT107), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n832), .B1(new_n835), .B2(new_n764), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n827), .B1(new_n829), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n832), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(new_n765), .B2(new_n766), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(KEYINPUT52), .A3(new_n776), .A4(new_n828), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n782), .A2(new_n644), .A3(new_n705), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n660), .B1(new_n773), .B2(new_n771), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n461), .B1(new_n676), .B2(new_n677), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n731), .A2(new_n511), .A3(new_n844), .A4(new_n698), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n842), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n788), .A3(new_n790), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n841), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n518), .B(new_n645), .C1(new_n375), .C2(new_n699), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n454), .A2(new_n461), .A3(new_n511), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n670), .B(new_n675), .C1(new_n851), .C2(new_n663), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n850), .A2(new_n852), .A3(KEYINPUT112), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n665), .A2(new_n737), .B1(new_n752), .B2(new_n753), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n747), .A3(new_n767), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n826), .B1(new_n849), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n847), .B1(new_n837), .B2(new_n840), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n754), .A2(new_n767), .A3(new_n740), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n683), .A2(new_n745), .A3(new_n737), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n745), .B1(new_n683), .B2(new_n737), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT114), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n858), .A2(new_n747), .A3(new_n868), .A4(new_n767), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n826), .B1(new_n855), .B2(new_n856), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n862), .A2(new_n867), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n860), .A2(new_n861), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n860), .A2(KEYINPUT113), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT113), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n874), .B(new_n826), .C1(new_n849), .C2(new_n859), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n850), .A2(new_n852), .A3(KEYINPUT112), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT112), .B1(new_n850), .B2(new_n852), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n878), .A2(new_n863), .A3(new_n866), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(KEYINPUT53), .A3(new_n862), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n873), .A2(new_n875), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n872), .B1(new_n881), .B2(KEYINPUT54), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n792), .A2(new_n513), .A3(new_n793), .ZN(new_n883));
  INV_X1    g697(.A(new_n761), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(new_n782), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT115), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n813), .A2(new_n814), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n821), .A2(new_n596), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n782), .A2(new_n736), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n771), .A2(new_n773), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n253), .A3(new_n513), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n722), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n454), .A2(new_n461), .A3(new_n658), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n892), .A2(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT50), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n718), .A2(new_n519), .A3(new_n736), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n885), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n899), .B1(new_n885), .B2(new_n901), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n898), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n890), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT51), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n890), .A2(KEYINPUT51), .A3(new_n905), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n883), .A2(new_n749), .A3(new_n884), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n895), .B1(new_n739), .B2(new_n738), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n910), .A2(G952), .A3(new_n223), .A4(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n375), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n892), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n914), .B(new_n915), .Z(new_n916));
  NAND2_X1  g730(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND4_X1   g732(.A1(new_n882), .A2(new_n908), .A3(new_n909), .A4(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(G952), .A2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n825), .B1(new_n919), .B2(new_n920), .ZN(G75));
  NOR2_X1   g735(.A1(new_n223), .A2(G952), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n187), .B1(new_n860), .B2(new_n871), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT56), .B1(new_n924), .B2(new_n590), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n555), .A2(new_n557), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n568), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n923), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(KEYINPUT117), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n925), .A2(KEYINPUT118), .A3(new_n930), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(G51));
  XOR2_X1   g749(.A(new_n799), .B(KEYINPUT57), .Z(new_n936));
  AOI21_X1  g750(.A(new_n861), .B1(new_n860), .B2(new_n871), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n872), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n732), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n798), .B(KEYINPUT119), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n924), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n922), .B1(new_n939), .B2(new_n941), .ZN(G54));
  NAND2_X1  g756(.A1(new_n860), .A2(new_n871), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n188), .ZN(new_n944));
  NAND2_X1  g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n451), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .A4(new_n436), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n923), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G60));
  INV_X1    g764(.A(new_n656), .ZN(new_n951));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT59), .Z(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AND4_X1   g769(.A1(new_n862), .A2(new_n867), .A3(new_n869), .A4(new_n870), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT53), .B1(new_n879), .B2(new_n862), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT54), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n860), .A2(new_n861), .A3(new_n871), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT121), .B1(new_n960), .B2(new_n922), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n954), .B1(new_n872), .B2(new_n937), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT121), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n963), .A3(new_n923), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT122), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n875), .A2(new_n880), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n957), .A2(new_n874), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT54), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n953), .B1(new_n969), .B2(new_n959), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n966), .B1(new_n970), .B2(new_n656), .ZN(new_n971));
  OAI211_X1 g785(.A(KEYINPUT122), .B(new_n951), .C1(new_n882), .C2(new_n953), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n965), .B1(new_n971), .B2(new_n972), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT60), .Z(new_n975));
  NAND2_X1  g789(.A1(new_n943), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n251), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n922), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n689), .A2(new_n690), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n976), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G66));
  OAI21_X1  g796(.A(G953), .B1(new_n515), .B2(new_n566), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT123), .Z(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n859), .B2(new_n223), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n926), .B1(G898), .B2(new_n223), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n985), .B(new_n986), .Z(G69));
  XNOR2_X1  g801(.A(new_n353), .B(KEYINPUT124), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n988), .B(new_n989), .Z(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(new_n620), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n991), .A2(new_n704), .A3(new_n223), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n709), .B1(new_n851), .B2(new_n663), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n993), .A2(new_n784), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n805), .B2(new_n806), .ZN(new_n995));
  INV_X1    g809(.A(new_n829), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n725), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT62), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(new_n725), .A3(KEYINPUT62), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n995), .A2(new_n819), .A3(new_n1001), .A4(new_n990), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n829), .B1(new_n805), .B2(new_n806), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n804), .A2(new_n913), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n765), .A2(new_n766), .ZN(new_n1005));
  OR3_X1    g819(.A1(new_n1004), .A2(KEYINPUT125), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT125), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n788), .A2(new_n790), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1003), .A2(new_n1008), .A3(new_n819), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1002), .B1(new_n1012), .B2(new_n990), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n992), .B1(new_n1013), .B2(new_n223), .ZN(G72));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT63), .Z(new_n1016));
  NAND3_X1  g830(.A1(new_n995), .A2(new_n819), .A3(new_n1001), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1016), .B1(new_n1017), .B2(new_n859), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(KEYINPUT126), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1020), .B(new_n1016), .C1(new_n1017), .C2(new_n859), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n354), .A2(new_n260), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n362), .A2(new_n332), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n881), .A2(new_n1016), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1016), .B1(new_n1011), .B2(new_n859), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n356), .A2(new_n261), .A3(new_n317), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n922), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1023), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT127), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1023), .A2(KEYINPUT127), .A3(new_n1025), .A4(new_n1028), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(G57));
endmodule


