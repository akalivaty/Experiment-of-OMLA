//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935;
  XNOR2_X1  g000(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n202));
  XNOR2_X1  g001(.A(G155gat), .B(G183gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT87), .ZN(new_n206));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207));
  INV_X1    g006(.A(G1gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT16), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n207), .A2(G1gat), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n210), .A2(new_n211), .A3(G8gat), .ZN(new_n212));
  INV_X1    g011(.A(G8gat), .ZN(new_n213));
  XOR2_X1   g012(.A(G15gat), .B(G22gat), .Z(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n207), .A2(new_n209), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n206), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(G8gat), .B1(new_n210), .B2(new_n211), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n215), .A2(new_n213), .A3(new_n216), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT87), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G71gat), .A2(G78gat), .ZN(new_n223));
  OR2_X1    g022(.A1(G71gat), .A2(G78gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT9), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G57gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G64gat), .ZN(new_n228));
  INV_X1    g027(.A(G64gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G57gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G71gat), .B2(G78gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT91), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(G71gat), .B2(G78gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n223), .A2(KEYINPUT91), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n223), .A2(KEYINPUT91), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(G71gat), .A3(G78gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n238), .A2(new_n239), .A3(new_n224), .A4(new_n232), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT92), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(new_n228), .B2(new_n230), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n225), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n229), .A2(G57gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n227), .A2(G64gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(KEYINPUT92), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n241), .A2(new_n248), .A3(KEYINPUT93), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT93), .B1(new_n241), .B2(new_n248), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n231), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT21), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n222), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n251), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(KEYINPUT21), .ZN(new_n256));
  INV_X1    g055(.A(G127gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n256), .A2(new_n257), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n254), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n260), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(new_n258), .A3(new_n253), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n205), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G231gat), .A2(G233gat), .ZN(new_n266));
  INV_X1    g065(.A(G211gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n261), .A2(new_n263), .A3(new_n205), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n265), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n268), .B1(new_n265), .B2(new_n269), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT15), .ZN(new_n274));
  NOR2_X1   g073(.A1(G29gat), .A2(G36gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(G29gat), .A2(G36gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(KEYINPUT14), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G43gat), .B(G50gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT14), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n279), .A2(G29gat), .A3(G36gat), .ZN(new_n280));
  OR4_X1    g079(.A1(new_n274), .A2(new_n277), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n274), .B1(new_n277), .B2(new_n280), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(KEYINPUT14), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n279), .B1(G29gat), .B2(G36gat), .ZN(new_n284));
  OAI211_X1 g083(.A(KEYINPUT15), .B(new_n283), .C1(new_n284), .C2(new_n275), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n285), .A3(new_n278), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n281), .A2(KEYINPUT17), .A3(new_n286), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n287), .A2(KEYINPUT86), .A3(new_n288), .ZN(new_n293));
  NAND2_X1  g092(.A1(G85gat), .A2(G92gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT7), .ZN(new_n295));
  NAND2_X1  g094(.A1(G99gat), .A2(G106gat), .ZN(new_n296));
  INV_X1    g095(.A(G85gat), .ZN(new_n297));
  INV_X1    g096(.A(G92gat), .ZN(new_n298));
  AOI22_X1  g097(.A1(KEYINPUT8), .A2(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G99gat), .B(G106gat), .Z(new_n301));
  OR2_X1    g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(KEYINPUT95), .A3(new_n301), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT95), .B1(new_n300), .B2(new_n301), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n287), .B(new_n302), .C1(new_n305), .C2(new_n304), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G190gat), .B(G218gat), .Z(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n307), .A2(new_n311), .A3(new_n308), .A4(new_n309), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT94), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(G134gat), .ZN(new_n318));
  INV_X1    g117(.A(G162gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n321), .A2(KEYINPUT96), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT96), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT97), .B1(new_n310), .B2(new_n312), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n324), .B1(new_n315), .B2(KEYINPUT97), .ZN(new_n325));
  INV_X1    g124(.A(new_n320), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n322), .B1(new_n327), .B2(new_n321), .ZN(new_n328));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(new_n229), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(new_n298), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n332));
  INV_X1    g131(.A(G169gat), .ZN(new_n333));
  INV_X1    g132(.A(G176gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT23), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT65), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n334), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n336), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n337), .A2(new_n338), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT66), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G183gat), .ZN(new_n346));
  INV_X1    g145(.A(G190gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT24), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(KEYINPUT24), .B2(new_n349), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n332), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT25), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n341), .A2(new_n335), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n351), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n357), .B(KEYINPUT68), .Z(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT27), .B(G183gat), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(new_n347), .ZN(new_n362));
  INV_X1    g161(.A(new_n349), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n339), .B(KEYINPUT26), .Z(new_n364));
  AOI211_X1 g163(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n338), .ZN(new_n365));
  OR3_X1    g164(.A1(new_n346), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT27), .B1(new_n346), .B2(KEYINPUT69), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n347), .A3(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n368), .A2(KEYINPUT70), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(KEYINPUT70), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n360), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n359), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(G226gat), .A3(G233gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n352), .A2(new_n358), .B1(new_n371), .B2(new_n365), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(KEYINPUT29), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT22), .ZN(new_n378));
  INV_X1    g177(.A(G218gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n378), .B1(new_n267), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT74), .ZN(new_n381));
  XNOR2_X1  g180(.A(G197gat), .B(G204gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n383), .B(new_n378), .C1(new_n267), .C2(new_n379), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G211gat), .B(G218gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  NAND3_X1  g186(.A1(new_n374), .A2(new_n377), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n374), .B2(new_n377), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n331), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n377), .ZN(new_n392));
  INV_X1    g191(.A(new_n387), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n331), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT75), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n396), .A2(new_n399), .A3(new_n397), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n396), .B2(new_n397), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n391), .B(new_n398), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(G127gat), .B(G134gat), .Z(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G120gat), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT72), .B1(new_n405), .B2(G113gat), .ZN(new_n406));
  INV_X1    g205(.A(G113gat), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT71), .B1(new_n407), .B2(G120gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT72), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n407), .A3(G120gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT71), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(new_n405), .A3(G113gat), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n406), .A2(new_n408), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT1), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n404), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G113gat), .B(G120gat), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n403), .B1(new_n416), .B2(KEYINPUT1), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT79), .ZN(new_n419));
  NAND2_X1  g218(.A1(G155gat), .A2(G162gat), .ZN(new_n420));
  INV_X1    g219(.A(G155gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n319), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n420), .B1(new_n422), .B2(KEYINPUT2), .ZN(new_n423));
  INV_X1    g222(.A(G141gat), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT77), .B1(new_n424), .B2(G148gat), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT76), .ZN(new_n426));
  INV_X1    g225(.A(G148gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(G141gat), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT77), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(new_n427), .A3(G141gat), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n424), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n425), .A2(new_n428), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT2), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n424), .A2(G148gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n427), .A2(G141gat), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n422), .A2(new_n420), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n423), .A2(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n438), .B(KEYINPUT78), .Z(new_n441));
  OAI211_X1 g240(.A(new_n419), .B(new_n440), .C1(new_n441), .C2(new_n439), .ZN(new_n442));
  INV_X1    g241(.A(new_n418), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n438), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n442), .B(new_n446), .C1(new_n444), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n441), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n419), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n444), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n451), .B(KEYINPUT39), .C1(new_n450), .C2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G1gat), .B(G29gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT0), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(G57gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(new_n297), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n455), .B(new_n459), .C1(KEYINPUT39), .C2(new_n451), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT40), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n454), .A2(new_n450), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n450), .B1(new_n444), .B2(new_n447), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n442), .B(new_n463), .C1(new_n445), .C2(new_n444), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(KEYINPUT5), .A3(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n450), .A2(KEYINPUT5), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(new_n448), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n459), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n402), .A2(new_n461), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G228gat), .A2(G233gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT82), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT29), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT3), .B1(new_n387), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(new_n438), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n387), .B1(new_n475), .B2(new_n440), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n478), .A2(new_n473), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n441), .B2(new_n476), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G22gat), .B(G78gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT31), .B(G50gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G106gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n485), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n481), .A2(new_n489), .A3(new_n483), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n486), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n402), .A2(new_n461), .A3(KEYINPUT84), .A4(new_n469), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n394), .A2(KEYINPUT37), .A3(new_n388), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT37), .B1(new_n394), .B2(new_n388), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n331), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n498), .A2(KEYINPUT38), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n467), .B2(new_n468), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(new_n469), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(KEYINPUT38), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n499), .A2(new_n502), .A3(new_n396), .A4(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n472), .A2(new_n494), .A3(new_n495), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n373), .A2(new_n443), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n376), .A2(new_n418), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G227gat), .A2(G233gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT64), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT34), .B1(new_n511), .B2(KEYINPUT73), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OR3_X1    g312(.A1(new_n508), .A2(KEYINPUT73), .A3(new_n510), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G43gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G71gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G99gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n506), .A2(new_n510), .A3(new_n507), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT33), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(KEYINPUT32), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n518), .B(KEYINPUT32), .C1(new_n519), .C2(new_n517), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n514), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n514), .B1(new_n523), .B2(new_n522), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n513), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n523), .ZN(new_n528));
  INV_X1    g327(.A(new_n514), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(new_n512), .A3(new_n524), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n527), .A2(KEYINPUT36), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT36), .B1(new_n527), .B2(new_n531), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n493), .B1(new_n402), .B2(new_n502), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n505), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n527), .A2(new_n531), .ZN(new_n537));
  INV_X1    g336(.A(new_n502), .ZN(new_n538));
  INV_X1    g337(.A(new_n402), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n537), .A2(new_n494), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT35), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n493), .B1(new_n527), .B2(new_n531), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n542), .A2(new_n543), .A3(new_n538), .A4(new_n539), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  AOI211_X1 g344(.A(new_n273), .B(new_n328), .C1(new_n536), .C2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G120gat), .B(G148gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(new_n334), .ZN(new_n548));
  INV_X1    g347(.A(G204gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT99), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT100), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n241), .A2(new_n248), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n241), .A2(new_n248), .A3(KEYINPUT93), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n300), .A2(new_n301), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n558), .A2(new_n231), .A3(new_n302), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n251), .A2(new_n306), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT10), .ZN(new_n564));
  INV_X1    g363(.A(new_n305), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(new_n565), .B2(new_n303), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n255), .A2(new_n302), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G230gat), .A2(G233gat), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n553), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n569), .ZN(new_n571));
  AOI211_X1 g370(.A(KEYINPUT100), .B(new_n571), .C1(new_n563), .C2(new_n567), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n560), .A2(new_n561), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n571), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n552), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n571), .B1(new_n563), .B2(new_n567), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n550), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n579), .A3(new_n575), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n212), .A2(new_n217), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n291), .A2(new_n292), .A3(new_n584), .A4(new_n293), .ZN(new_n585));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n218), .A2(new_n221), .A3(new_n287), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT18), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT88), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n222), .A2(new_n281), .A3(new_n286), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n587), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n586), .B(KEYINPUT13), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n218), .A2(new_n287), .A3(KEYINPUT89), .A4(new_n221), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n589), .A2(KEYINPUT88), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G197gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT11), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G169gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n583), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n546), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(new_n538), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n208), .ZN(G1324gat));
  OAI21_X1  g417(.A(G8gat), .B1(new_n616), .B2(new_n539), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT42), .ZN(new_n620));
  INV_X1    g419(.A(new_n616), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT101), .B(G8gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT16), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n402), .A3(new_n623), .ZN(new_n624));
  MUX2_X1   g423(.A(KEYINPUT42), .B(new_n620), .S(new_n624), .Z(G1325gat));
  INV_X1    g424(.A(new_n534), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n621), .A2(G15gat), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(G15gat), .B1(new_n621), .B2(new_n537), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(G1326gat));
  NOR2_X1   g428(.A1(new_n616), .A2(new_n494), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT43), .B(G22gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(G1327gat));
  NAND2_X1  g431(.A1(new_n315), .A2(KEYINPUT97), .ZN(new_n633));
  INV_X1    g432(.A(new_n324), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n326), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(KEYINPUT96), .A3(new_n321), .ZN(new_n636));
  INV_X1    g435(.A(new_n322), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n536), .B2(new_n545), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI211_X1 g440(.A(KEYINPUT44), .B(new_n638), .C1(new_n536), .C2(new_n545), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n272), .A2(new_n614), .A3(new_n583), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT102), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n502), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(G29gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n639), .A2(new_n644), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n649), .A2(G29gat), .A3(new_n538), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT45), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(G1328gat));
  NAND2_X1  g451(.A1(new_n646), .A2(new_n402), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(G36gat), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n649), .A2(G36gat), .A3(new_n539), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT46), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(G1329gat));
  INV_X1    g456(.A(new_n537), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n649), .A2(G43gat), .A3(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n626), .B(new_n645), .C1(new_n641), .C2(new_n642), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n660), .B2(G43gat), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(KEYINPUT103), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g462(.A(G50gat), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n639), .A2(new_n664), .A3(new_n493), .A4(new_n644), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n493), .B(new_n645), .C1(new_n641), .C2(new_n642), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT104), .ZN(new_n667));
  OAI211_X1 g466(.A(KEYINPUT48), .B(new_n665), .C1(new_n667), .C2(new_n664), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(G50gat), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n669), .A2(new_n665), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(KEYINPUT48), .B2(new_n670), .ZN(G1331gat));
  NAND3_X1  g470(.A1(new_n272), .A2(new_n638), .A3(new_n614), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n536), .B2(new_n545), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n538), .A2(new_n582), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n583), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n402), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT105), .ZN(new_n681));
  NOR2_X1   g480(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1333gat));
  OAI21_X1  g482(.A(G71gat), .B1(new_n677), .B2(new_n534), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n658), .A2(G71gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n677), .B2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g486(.A1(new_n678), .A2(new_n493), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g488(.A1(new_n273), .A2(new_n614), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT106), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n643), .A2(new_n674), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G85gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n639), .A2(new_n691), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT51), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n639), .A2(KEYINPUT51), .A3(new_n691), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT107), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n694), .B2(new_n695), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n674), .A2(new_n297), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n693), .B1(new_n701), .B2(new_n702), .ZN(G1336gat));
  NAND3_X1  g502(.A1(new_n402), .A2(new_n298), .A3(new_n583), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT108), .Z(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(new_n698), .B2(new_n700), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT52), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n583), .B(new_n691), .C1(new_n641), .C2(new_n642), .ZN(new_n708));
  OAI21_X1  g507(.A(G92gat), .B1(new_n708), .B2(new_n539), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n696), .ZN(new_n711));
  INV_X1    g510(.A(new_n697), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n705), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n707), .B1(new_n709), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT109), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n709), .A2(new_n713), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n707), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n719), .ZN(G1337gat));
  OAI21_X1  g519(.A(G99gat), .B1(new_n708), .B2(new_n534), .ZN(new_n721));
  OR3_X1    g520(.A1(new_n701), .A2(G99gat), .A3(new_n582), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(new_n658), .ZN(G1338gat));
  OR3_X1    g522(.A1(new_n708), .A2(KEYINPUT111), .A3(new_n494), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT111), .B1(new_n708), .B2(new_n494), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(G106gat), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT53), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n494), .A2(G106gat), .A3(new_n582), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n698), .B2(new_n700), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n711), .B2(new_n712), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G106gat), .B1(new_n708), .B2(new_n494), .ZN(new_n734));
  OAI211_X1 g533(.A(KEYINPUT110), .B(new_n728), .C1(new_n711), .C2(new_n712), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n730), .B1(new_n727), .B2(new_n736), .ZN(G1339gat));
  INV_X1    g536(.A(KEYINPUT118), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n539), .A2(new_n502), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n658), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT116), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n563), .A2(new_n742), .A3(new_n571), .A4(new_n567), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(KEYINPUT54), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n563), .A2(new_n571), .A3(new_n567), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n577), .B2(KEYINPUT113), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT54), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n570), .B2(new_n572), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n749), .A3(new_n550), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n747), .A2(new_n749), .A3(KEYINPUT55), .A4(new_n550), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n752), .A2(new_n613), .A3(new_n580), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n597), .A2(new_n600), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n598), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n585), .A2(new_n587), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(G229gat), .A3(G233gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n608), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n594), .A2(new_n603), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n611), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n576), .B2(new_n581), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n638), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n752), .A2(new_n761), .A3(new_n580), .A4(new_n753), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n766), .A2(new_n638), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n328), .B1(new_n754), .B2(new_n762), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n766), .A2(new_n638), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT114), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(new_n273), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n272), .A2(new_n638), .A3(new_n582), .A4(new_n614), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT112), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n772), .A2(KEYINPUT115), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT115), .B1(new_n772), .B2(new_n774), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n741), .B1(new_n777), .B2(new_n494), .ZN(new_n778));
  NOR4_X1   g577(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT116), .A4(new_n493), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n740), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT117), .B(new_n740), .C1(new_n778), .C2(new_n779), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n613), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G113gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n772), .A2(new_n774), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n774), .A3(KEYINPUT115), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n538), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n542), .A2(new_n539), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n793), .A2(G113gat), .A3(new_n614), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n738), .B1(new_n785), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g595(.A(KEYINPUT118), .B(new_n794), .C1(new_n784), .C2(G113gat), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(G1340gat));
  INV_X1    g597(.A(new_n793), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n405), .A3(new_n583), .ZN(new_n800));
  INV_X1    g599(.A(new_n782), .ZN(new_n801));
  INV_X1    g600(.A(new_n783), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n801), .A2(new_n802), .A3(new_n582), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n803), .B2(new_n405), .ZN(G1341gat));
  AOI21_X1  g603(.A(G127gat), .B1(new_n799), .B2(new_n272), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n801), .A2(new_n802), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n273), .A2(new_n257), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(G1342gat));
  NOR3_X1   g607(.A1(new_n793), .A2(G134gat), .A3(new_n638), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT56), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n801), .A2(new_n802), .A3(new_n638), .ZN(new_n811));
  INV_X1    g610(.A(G134gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(G1343gat));
  NOR2_X1   g612(.A1(new_n626), .A2(new_n494), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n790), .A2(new_n538), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT120), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n614), .A2(G141gat), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n818), .A2(new_n402), .A3(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n752), .A2(KEYINPUT119), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n753), .A2(new_n580), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n822), .A2(new_n614), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(KEYINPUT119), .B2(new_n752), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n762), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n638), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n272), .B1(new_n827), .B2(new_n767), .ZN(new_n828));
  INV_X1    g627(.A(new_n774), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n493), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI211_X1 g629(.A(new_n626), .B(new_n739), .C1(new_n830), .C2(KEYINPUT57), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n777), .A2(new_n832), .A3(new_n493), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n613), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G141gat), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n816), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n402), .A3(new_n820), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n834), .B2(G141gat), .ZN(new_n840));
  OAI22_X1  g639(.A1(new_n821), .A2(new_n837), .B1(new_n836), .B2(new_n840), .ZN(G1344gat));
  NOR2_X1   g640(.A1(new_n818), .A2(new_n402), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n427), .A3(new_n583), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT57), .B1(new_n790), .B2(new_n494), .ZN(new_n845));
  INV_X1    g644(.A(new_n773), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n832), .B(new_n493), .C1(new_n828), .C2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n583), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n626), .A2(new_n739), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n844), .B1(new_n851), .B2(G148gat), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n831), .A2(new_n833), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n844), .B1(new_n853), .B2(new_n582), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n427), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n843), .B1(new_n852), .B2(new_n855), .ZN(G1345gat));
  NAND4_X1  g655(.A1(new_n817), .A2(new_n421), .A3(new_n272), .A4(new_n539), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n853), .A2(new_n273), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n421), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT121), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n857), .B(new_n861), .C1(new_n421), .C2(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1346gat));
  NAND3_X1  g662(.A1(new_n842), .A2(new_n319), .A3(new_n328), .ZN(new_n864));
  OAI21_X1  g663(.A(G162gat), .B1(new_n853), .B2(new_n638), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1347gat));
  OAI21_X1  g665(.A(KEYINPUT122), .B1(new_n790), .B2(new_n502), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n777), .A2(new_n868), .A3(new_n538), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(new_n542), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n402), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n333), .A3(new_n613), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n538), .A2(new_n402), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n658), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT123), .Z(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n778), .B2(new_n779), .ZN(new_n878));
  OAI21_X1  g677(.A(G169gat), .B1(new_n878), .B2(new_n614), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n873), .A2(new_n879), .ZN(G1348gat));
  NOR3_X1   g679(.A1(new_n878), .A2(new_n334), .A3(new_n582), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n872), .A2(new_n583), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n334), .ZN(G1349gat));
  NAND4_X1  g682(.A1(new_n871), .A2(new_n272), .A3(new_n361), .A4(new_n402), .ZN(new_n884));
  OAI21_X1  g683(.A(G183gat), .B1(new_n878), .B2(new_n273), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT60), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n884), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(G1350gat));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n347), .A3(new_n328), .ZN(new_n891));
  INV_X1    g690(.A(new_n878), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n347), .B1(new_n892), .B2(new_n328), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(G1351gat));
  NAND3_X1  g696(.A1(new_n870), .A2(new_n402), .A3(new_n814), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT124), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n815), .B1(new_n867), .B2(new_n869), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n402), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n614), .A2(G197gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n626), .A2(new_n874), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n848), .A2(new_n613), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G197gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n904), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(new_n899), .B2(new_n902), .ZN(new_n912));
  INV_X1    g711(.A(new_n909), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT125), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n910), .A2(new_n914), .ZN(G1352gat));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n549), .A3(new_n583), .A4(new_n402), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n849), .A2(new_n907), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G204gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n917), .A2(KEYINPUT126), .A3(new_n918), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n916), .B2(KEYINPUT62), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n919), .B(new_n921), .C1(new_n922), .C2(new_n924), .ZN(G1353gat));
  NAND3_X1  g724(.A1(new_n848), .A2(new_n272), .A3(new_n907), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n926), .A2(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n903), .A2(new_n267), .A3(new_n272), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n926), .A2(new_n930), .A3(new_n931), .A4(G211gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n929), .A3(new_n932), .ZN(G1354gat));
  AND4_X1   g732(.A1(G218gat), .A2(new_n848), .A3(new_n328), .A4(new_n907), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n903), .A2(new_n328), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(new_n379), .ZN(G1355gat));
endmodule


