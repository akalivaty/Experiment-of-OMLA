//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(G134), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n192), .A3(G131), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(G128), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n200), .B(new_n202), .C1(KEYINPUT1), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT67), .B1(new_n205), .B2(new_n207), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n198), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G143), .B(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT0), .A3(G128), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT0), .B(G128), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT65), .A2(G131), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n193), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n189), .A2(new_n191), .A3(new_n192), .A4(new_n218), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n220), .A2(KEYINPUT66), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT66), .B1(new_n220), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n217), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n212), .A2(new_n224), .A3(KEYINPUT30), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n205), .A2(new_n207), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n198), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n221), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n227), .B1(new_n216), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G116), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G119), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT2), .B(G113), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n238), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n225), .A2(new_n232), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(G237), .A2(G953), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G210), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT27), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G101), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n241), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n212), .A2(new_n224), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n242), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n242), .A2(KEYINPUT68), .A3(new_n247), .A4(new_n249), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(KEYINPUT31), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT69), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n252), .A2(new_n256), .A3(KEYINPUT31), .A4(new_n253), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT31), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n242), .A2(new_n258), .A3(new_n247), .A4(new_n249), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n212), .A2(new_n224), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n248), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n249), .A2(KEYINPUT28), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n262), .A2(new_n263), .B1(new_n241), .B2(new_n230), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n259), .B1(new_n264), .B2(new_n247), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n255), .A2(new_n257), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT32), .ZN(new_n268));
  NOR2_X1   g082(.A1(G472), .A2(G902), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n247), .B1(new_n242), .B2(new_n249), .ZN(new_n273));
  AOI211_X1 g087(.A(KEYINPUT29), .B(new_n273), .C1(new_n264), .C2(new_n247), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n260), .A2(new_n248), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n263), .B2(new_n262), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT29), .A3(new_n247), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G472), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G469), .ZN(new_n282));
  XNOR2_X1  g096(.A(G110), .B(G140), .ZN(new_n283));
  INV_X1    g097(.A(G953), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n284), .A2(G227), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n283), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G104), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT71), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G104), .ZN(new_n290));
  AOI21_X1  g104(.A(G107), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G107), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(G104), .ZN(new_n293));
  OAI21_X1  g107(.A(G101), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n287), .A2(KEYINPUT3), .A3(G107), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n288), .A2(new_n290), .A3(G107), .ZN(new_n299));
  INV_X1    g113(.A(G101), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n294), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n208), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT71), .B(G104), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT3), .B1(new_n304), .B2(G107), .ZN(new_n305));
  AOI21_X1  g119(.A(G101), .B1(new_n304), .B2(G107), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n296), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n226), .A2(new_n307), .A3(new_n294), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n303), .A2(KEYINPUT74), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n302), .A2(new_n310), .A3(new_n208), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n309), .A2(KEYINPUT12), .A3(new_n228), .A4(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n222), .A2(new_n223), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n309), .A2(new_n315), .A3(new_n311), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT12), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT75), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(new_n320), .A3(new_n317), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n313), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n305), .A2(new_n299), .A3(new_n296), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT73), .B(KEYINPUT4), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(G101), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n217), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n288), .A2(new_n290), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n292), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n295), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n300), .B1(new_n330), .B2(new_n299), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT4), .B1(new_n298), .B2(new_n301), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n330), .B2(new_n306), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n323), .A2(G101), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(KEYINPUT72), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n326), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n302), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n339), .B(KEYINPUT10), .C1(new_n210), .C2(new_n211), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n308), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n338), .A2(new_n343), .A3(new_n315), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n286), .B1(new_n322), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n286), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n315), .B1(new_n338), .B2(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n282), .B1(new_n349), .B2(new_n278), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n352));
  INV_X1    g166(.A(new_n338), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n340), .A2(new_n342), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n314), .ZN(new_n355));
  INV_X1    g169(.A(new_n286), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n352), .B1(new_n322), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n316), .A2(new_n320), .A3(new_n317), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n320), .B1(new_n316), .B2(new_n317), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n312), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n346), .A3(KEYINPUT76), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n356), .B1(new_n355), .B2(new_n347), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(G902), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT77), .B1(new_n366), .B2(new_n282), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n358), .B2(new_n362), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n369));
  NOR4_X1   g183(.A1(new_n368), .A2(new_n369), .A3(G469), .A4(G902), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n351), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT9), .B(G234), .ZN(new_n372));
  OAI21_X1  g186(.A(G221), .B1(new_n372), .B2(G902), .ZN(new_n373));
  OAI21_X1  g187(.A(G214), .B1(G237), .B2(G902), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G110), .B(G122), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT79), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n234), .A2(new_n236), .A3(KEYINPUT5), .ZN(new_n378));
  OAI21_X1  g192(.A(G113), .B1(new_n234), .B2(KEYINPUT5), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n239), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n302), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n325), .A2(new_n241), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n331), .A2(new_n332), .A3(new_n327), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT72), .B1(new_n335), .B2(new_n336), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n382), .B1(new_n387), .B2(KEYINPUT78), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n383), .B1(new_n333), .B2(new_n337), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT78), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n377), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n381), .B1(new_n389), .B2(new_n390), .ZN(new_n393));
  INV_X1    g207(.A(new_n377), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n387), .A2(KEYINPUT78), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(KEYINPUT6), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT81), .B1(new_n216), .B2(G125), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n216), .A2(G125), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(G125), .B2(new_n226), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n400), .B2(KEYINPUT81), .ZN(new_n401));
  INV_X1    g215(.A(G224), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G953), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT82), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n401), .B(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n393), .A2(new_n395), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n407));
  AND4_X1   g221(.A1(KEYINPUT80), .A2(new_n406), .A3(new_n407), .A4(new_n377), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n394), .B1(new_n393), .B2(new_n395), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT80), .B1(new_n409), .B2(new_n407), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n397), .B(new_n405), .C1(new_n408), .C2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n401), .A2(KEYINPUT7), .A3(new_n404), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n404), .A2(KEYINPUT7), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n400), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n381), .A2(KEYINPUT83), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n302), .A2(new_n380), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n416), .B(new_n417), .Z(new_n418));
  XOR2_X1   g232(.A(new_n377), .B(KEYINPUT8), .Z(new_n419));
  AOI21_X1  g233(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n420), .B2(new_n396), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n411), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n411), .A2(new_n421), .A3(new_n423), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n375), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n281), .A2(new_n371), .A3(new_n373), .A4(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT90), .ZN(new_n429));
  AND2_X1   g243(.A1(KEYINPUT86), .A2(G122), .ZN(new_n430));
  NOR2_X1   g244(.A1(KEYINPUT86), .A2(G122), .ZN(new_n431));
  OAI21_X1  g245(.A(G116), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n432), .B(KEYINPUT87), .Z(new_n433));
  NAND2_X1  g247(.A1(new_n235), .A2(G122), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n292), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n432), .B(KEYINPUT87), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n434), .B(KEYINPUT14), .ZN(new_n437));
  OAI21_X1  g251(.A(G107), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G128), .B(G143), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n188), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G217), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n372), .A2(new_n442), .A3(G953), .ZN(new_n443));
  INV_X1    g257(.A(new_n434), .ZN(new_n444));
  OAI21_X1  g258(.A(G107), .B1(new_n436), .B2(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n435), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT13), .B1(new_n206), .B2(G143), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(new_n188), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n448), .B(new_n439), .Z(new_n449));
  OAI211_X1 g263(.A(new_n441), .B(new_n443), .C1(new_n446), .C2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n443), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n435), .A2(new_n438), .A3(new_n440), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n449), .B1(new_n435), .B2(new_n445), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT89), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n452), .A2(new_n453), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(KEYINPUT88), .A3(new_n443), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n456), .A2(new_n457), .A3(new_n278), .A4(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G478), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT15), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n460), .A2(new_n462), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n429), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n465), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(KEYINPUT90), .A3(new_n463), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n243), .A2(G214), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(new_n201), .ZN(new_n471));
  AOI21_X1  g285(.A(G143), .B1(new_n243), .B2(G214), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(new_n194), .ZN(new_n474));
  XNOR2_X1  g288(.A(G125), .B(G140), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT16), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT16), .ZN(new_n477));
  INV_X1    g291(.A(G140), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(G125), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(G146), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(KEYINPUT84), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT19), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n474), .B(new_n480), .C1(G146), .C2(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n471), .A2(new_n472), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(KEYINPUT18), .A3(G131), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT18), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n473), .B1(new_n486), .B2(new_n194), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n475), .B(new_n199), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G113), .B(G122), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(new_n287), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n480), .ZN(new_n495));
  AOI21_X1  g309(.A(G146), .B1(new_n476), .B2(new_n479), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n484), .A2(KEYINPUT17), .A3(G131), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n497), .B(new_n498), .C1(new_n474), .C2(KEYINPUT17), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n492), .A3(new_n489), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(G475), .A2(G902), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT85), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(KEYINPUT20), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n501), .B2(new_n502), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n509));
  INV_X1    g323(.A(new_n500), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n492), .B1(new_n499), .B2(new_n489), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n278), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n508), .A2(new_n509), .B1(new_n512), .B2(G475), .ZN(new_n513));
  NAND2_X1  g327(.A1(G234), .A2(G237), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(G952), .A3(new_n284), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT21), .B(G898), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(G902), .A3(G953), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n507), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n469), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n442), .B1(G234), .B2(new_n278), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT23), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n233), .B2(G128), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n526), .B(new_n527), .C1(G119), .C2(new_n206), .ZN(new_n528));
  XNOR2_X1  g342(.A(G119), .B(G128), .ZN(new_n529));
  XOR2_X1   g343(.A(KEYINPUT24), .B(G110), .Z(new_n530));
  AOI22_X1  g344(.A1(new_n528), .A2(G110), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n495), .B2(new_n496), .ZN(new_n532));
  OAI22_X1  g346(.A1(new_n528), .A2(G110), .B1(new_n529), .B2(new_n530), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n475), .A2(new_n199), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n480), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n284), .A2(G221), .A3(G234), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT70), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT22), .B(G137), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n540), .B1(new_n532), .B2(new_n535), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n524), .B1(new_n544), .B2(G902), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT25), .B(new_n278), .C1(new_n542), .C2(new_n543), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n523), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n542), .A2(new_n543), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n522), .A2(G902), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n521), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n428), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT91), .B(G101), .Z(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(G3));
  NOR3_X1   g368(.A1(new_n322), .A2(new_n352), .A3(new_n357), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT76), .B1(new_n361), .B2(new_n346), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n365), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(new_n282), .A3(new_n278), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n369), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n366), .A2(KEYINPUT77), .A3(new_n282), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n350), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n373), .ZN(new_n562));
  INV_X1    g376(.A(new_n550), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n411), .A2(new_n421), .A3(new_n423), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n423), .B1(new_n411), .B2(new_n421), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n374), .B(new_n519), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G472), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n267), .B2(new_n278), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT92), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n267), .A2(new_n278), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G472), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n267), .A2(new_n269), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n571), .B1(new_n575), .B2(KEYINPUT92), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n564), .A2(new_n568), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n461), .A2(G902), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n450), .A2(KEYINPUT93), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n454), .ZN(new_n581));
  OAI211_X1 g395(.A(KEYINPUT93), .B(new_n451), .C1(new_n452), .C2(new_n453), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT33), .B1(new_n456), .B2(new_n459), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n578), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n456), .A2(new_n459), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n461), .B1(new_n586), .B2(G902), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n507), .A2(new_n513), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n588), .A2(KEYINPUT94), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT94), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n577), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT34), .B(G104), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  AND2_X1   g409(.A1(new_n507), .A2(new_n513), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n469), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n567), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n564), .A2(new_n576), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT35), .B(G107), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G9));
  NOR2_X1   g415(.A1(new_n561), .A2(new_n562), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT95), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT96), .B1(new_n540), .B2(KEYINPUT36), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT36), .ZN(new_n606));
  INV_X1    g420(.A(new_n538), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n607), .A2(new_n539), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n539), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n605), .B(new_n606), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n603), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n536), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n604), .A2(new_n610), .A3(new_n603), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n604), .A2(new_n610), .A3(new_n603), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n536), .B1(new_n616), .B2(new_n611), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n549), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n545), .A2(new_n546), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n522), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n621), .A3(KEYINPUT97), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n623));
  INV_X1    g437(.A(new_n549), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n615), .B2(new_n617), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n623), .B1(new_n625), .B2(new_n547), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n520), .B(new_n627), .C1(new_n466), .C2(new_n468), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n570), .A2(KEYINPUT92), .ZN(new_n629));
  INV_X1    g443(.A(new_n574), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT92), .B1(new_n630), .B2(new_n570), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n602), .A2(new_n632), .A3(new_n427), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT98), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n633), .B(new_n635), .ZN(G12));
  XNOR2_X1  g450(.A(new_n515), .B(KEYINPUT99), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(G900), .B2(new_n518), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT100), .Z(new_n639));
  NOR2_X1   g453(.A1(new_n589), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n627), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n469), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n428), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT101), .B(G128), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G30));
  NOR2_X1   g461(.A1(new_n565), .A2(new_n566), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n648), .A2(KEYINPUT38), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(KEYINPUT38), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n252), .A2(new_n253), .ZN(new_n652));
  INV_X1    g466(.A(new_n249), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n275), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n247), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n278), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(G472), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n270), .B2(new_n271), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n466), .A2(new_n468), .A3(new_n589), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n625), .A2(new_n547), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n374), .A3(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n651), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n639), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n602), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n664), .B1(KEYINPUT40), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n201), .ZN(G45));
  INV_X1    g485(.A(new_n588), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n596), .ZN(new_n673));
  INV_X1    g487(.A(new_n639), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n428), .A2(new_n627), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n199), .ZN(G48));
  OAI21_X1  g491(.A(G469), .B1(new_n368), .B2(G902), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n373), .B(new_n678), .C1(new_n367), .C2(new_n370), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT103), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n563), .B1(new_n272), .B2(new_n280), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n559), .A2(new_n560), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n373), .A4(new_n678), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n592), .A2(new_n567), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n680), .A2(new_n681), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NAND4_X1  g502(.A1(new_n680), .A2(new_n681), .A3(new_n684), .A4(new_n598), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  NAND3_X1  g504(.A1(new_n680), .A2(new_n427), .A3(new_n684), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT104), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n680), .A2(new_n693), .A3(new_n684), .A4(new_n427), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n281), .A2(new_n628), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  XOR2_X1   g513(.A(new_n269), .B(KEYINPUT105), .Z(new_n700));
  AND3_X1   g514(.A1(new_n252), .A2(KEYINPUT31), .A3(new_n253), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n259), .B1(new_n276), .B2(new_n247), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(KEYINPUT106), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n573), .A2(new_n707), .A3(new_n550), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n567), .A2(new_n708), .A3(new_n660), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n680), .A2(new_n709), .A3(new_n684), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND2_X1  g525(.A1(new_n573), .A2(new_n707), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n675), .A2(new_n662), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n695), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n345), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g531(.A(KEYINPUT107), .B(new_n286), .C1(new_n322), .C2(new_n344), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n348), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n282), .B1(new_n719), .B2(new_n278), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n559), .B2(new_n560), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT108), .B1(new_n721), .B2(new_n562), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n565), .A2(new_n566), .A3(new_n375), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n719), .A2(new_n278), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n367), .B2(new_n370), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n373), .ZN(new_n728));
  AND4_X1   g542(.A1(new_n681), .A2(new_n722), .A3(new_n723), .A4(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n675), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(KEYINPUT42), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n722), .A2(new_n728), .A3(new_n681), .A4(new_n723), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n732), .B1(new_n733), .B2(new_n675), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  NAND2_X1  g550(.A1(new_n469), .A2(new_n640), .ZN(new_n737));
  XOR2_X1   g551(.A(new_n737), .B(KEYINPUT109), .Z(new_n738));
  NOR2_X1   g552(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n188), .ZN(G36));
  NAND2_X1  g554(.A1(new_n648), .A2(new_n374), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT110), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n741), .A2(KEYINPUT110), .ZN(new_n743));
  INV_X1    g557(.A(new_n576), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n596), .A2(new_n588), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(KEYINPUT43), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(KEYINPUT43), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n747), .A2(new_n748), .A3(new_n662), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n744), .A2(new_n745), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n745), .B1(new_n744), .B2(new_n749), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n742), .B(new_n743), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n282), .A2(new_n278), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n719), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n349), .ZN(new_n757));
  OAI21_X1  g571(.A(G469), .B1(new_n757), .B2(KEYINPUT45), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n754), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n682), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n373), .A3(new_n666), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n752), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n190), .ZN(G39));
  NOR4_X1   g580(.A1(new_n281), .A2(new_n741), .A3(new_n675), .A4(new_n550), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n373), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT47), .B1(new_n763), .B2(new_n373), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n770), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n768), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(KEYINPUT111), .A3(new_n767), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n374), .B1(new_n649), .B2(new_n650), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n747), .A2(new_n708), .A3(new_n748), .A4(new_n637), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n680), .A3(new_n781), .A4(new_n684), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(KEYINPUT50), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n782), .B(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n680), .A2(new_n684), .A3(new_n723), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n563), .A2(new_n515), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n786), .A2(new_n659), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n596), .A3(new_n672), .ZN(new_n789));
  INV_X1    g603(.A(new_n637), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n747), .A2(new_n748), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n786), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n712), .A2(new_n662), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n785), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n781), .A2(new_n743), .A3(new_n742), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT115), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n769), .A2(new_n770), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n682), .A2(new_n678), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n682), .A2(KEYINPUT116), .A3(new_n678), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n562), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n797), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n779), .B1(new_n795), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(G952), .ZN(new_n806));
  INV_X1    g620(.A(new_n592), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n806), .B(G953), .C1(new_n788), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT48), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n792), .A2(new_n809), .A3(new_n681), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n786), .A2(new_n790), .A3(new_n791), .ZN(new_n811));
  INV_X1    g625(.A(new_n681), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT48), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n695), .A2(new_n781), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n808), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n805), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n795), .ZN(new_n818));
  INV_X1    g632(.A(new_n797), .ZN(new_n819));
  INV_X1    g633(.A(new_n803), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n819), .B1(new_n775), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n818), .A2(KEYINPUT51), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT118), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n818), .A2(new_n824), .A3(KEYINPUT51), .A4(new_n821), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n817), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n427), .A2(new_n661), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n562), .B1(new_n682), .B2(new_n725), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n625), .A2(new_n547), .A3(new_n639), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n658), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n828), .A2(new_n829), .A3(new_n831), .A4(KEYINPUT114), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n726), .A2(new_n373), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n427), .A2(new_n658), .A3(new_n661), .A4(new_n830), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n371), .A2(new_n373), .A3(new_n427), .ZN(new_n838));
  INV_X1    g652(.A(new_n644), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n675), .A2(new_n627), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n838), .B(new_n281), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n714), .A2(new_n842), .A3(KEYINPUT52), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  INV_X1    g658(.A(new_n713), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n692), .B2(new_n694), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n837), .A2(new_n841), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n722), .A2(new_n728), .A3(new_n713), .A4(new_n723), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT113), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n741), .B1(new_n829), .B2(new_n727), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n853), .A3(new_n713), .A4(new_n722), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n642), .A2(new_n465), .A3(new_n464), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n281), .A2(new_n602), .A3(new_n723), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n738), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n857), .B1(new_n729), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT42), .B1(new_n729), .B2(new_n730), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n733), .A2(new_n732), .A3(new_n675), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n855), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n589), .B1(new_n467), .B2(new_n463), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n564), .A2(new_n568), .A3(new_n576), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n689), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n686), .A2(new_n710), .A3(new_n633), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n673), .A2(new_n564), .A3(new_n568), .A4(new_n576), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT112), .B1(new_n869), .B2(new_n552), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT112), .ZN(new_n871));
  INV_X1    g685(.A(new_n673), .ZN(new_n872));
  OAI221_X1 g686(.A(new_n871), .B1(new_n428), .B2(new_n551), .C1(new_n577), .C2(new_n872), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n698), .A2(new_n868), .A3(new_n870), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n849), .A2(new_n863), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n698), .A2(new_n868), .A3(new_n870), .A4(new_n873), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n862), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(KEYINPUT53), .A3(new_n849), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n877), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  AND4_X1   g696(.A1(KEYINPUT53), .A2(new_n849), .A3(new_n863), .A4(new_n874), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n880), .B2(new_n849), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT54), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n826), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n826), .A2(new_n885), .A3(KEYINPUT119), .A4(new_n882), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n806), .A2(new_n284), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n799), .B(KEYINPUT49), .Z(new_n892));
  NOR4_X1   g706(.A1(new_n746), .A2(new_n562), .A3(new_n375), .A4(new_n563), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n651), .A3(new_n659), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n891), .A2(new_n894), .ZN(G75));
  AOI21_X1  g709(.A(new_n278), .B1(new_n877), .B2(new_n881), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(G210), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n397), .B1(new_n408), .B2(new_n410), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n405), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT55), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n897), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n897), .B2(new_n898), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n284), .A2(G952), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G51));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n885), .A2(new_n906), .A3(new_n882), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n877), .A2(new_n881), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n753), .B(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n557), .ZN(new_n912));
  INV_X1    g726(.A(new_n896), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n913), .A2(new_n756), .A3(new_n758), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n904), .B1(new_n912), .B2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n500), .A3(new_n494), .ZN(new_n917));
  INV_X1    g731(.A(new_n904), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .A4(new_n501), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(G60));
  INV_X1    g734(.A(new_n583), .ZN(new_n921));
  INV_X1    g735(.A(new_n584), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AND4_X1   g740(.A1(new_n923), .A2(new_n907), .A3(new_n909), .A4(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(new_n885), .B2(new_n882), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n918), .B1(new_n928), .B2(new_n923), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(G63));
  XNOR2_X1  g744(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n442), .A2(new_n278), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n908), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n544), .B(KEYINPUT122), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n908), .A2(new_n618), .A3(new_n933), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n918), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n936), .A2(KEYINPUT61), .A3(new_n918), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G66));
  OAI21_X1  g756(.A(G953), .B1(new_n516), .B2(new_n402), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n874), .B2(G953), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n899), .B1(G898), .B2(new_n284), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT123), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n944), .B(new_n946), .ZN(G69));
  NAND2_X1  g761(.A1(new_n225), .A2(new_n232), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n482), .B(KEYINPUT124), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(G900), .A2(G953), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n846), .A2(new_n645), .A3(new_n676), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n764), .A2(new_n812), .A3(new_n827), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n765), .A2(new_n953), .A3(new_n739), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n777), .A2(new_n735), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n950), .B(new_n951), .C1(new_n955), .C2(G953), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n714), .B(new_n841), .C1(new_n669), .C2(new_n668), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n681), .B(new_n723), .C1(new_n673), .C2(new_n864), .ZN(new_n959));
  OAI22_X1  g773(.A1(new_n752), .A2(new_n764), .B1(new_n667), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n773), .B2(new_n776), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n958), .A2(new_n961), .A3(new_n965), .A4(new_n962), .ZN(new_n966));
  AOI21_X1  g780(.A(G953), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n956), .B1(new_n967), .B2(new_n950), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n284), .B1(G227), .B2(G900), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n969), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n971), .B(new_n956), .C1(new_n967), .C2(new_n950), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(G72));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n652), .B2(new_n273), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT127), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n908), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n975), .B1(new_n955), .B2(new_n879), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n242), .A2(new_n249), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n247), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n978), .A2(new_n982), .A3(new_n918), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n964), .A2(new_n874), .A3(new_n966), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT126), .B1(new_n984), .B2(new_n975), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n980), .A2(new_n247), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n984), .A2(KEYINPUT126), .A3(new_n975), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(G57));
endmodule


