//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n461), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n464), .A2(new_n468), .ZN(G160));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n460), .A2(new_n462), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G124), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT64), .ZN(new_n473));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n476), .B1(new_n461), .B2(G136), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n470), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n473), .A2(new_n470), .A3(new_n477), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n462), .C1(new_n458), .C2(new_n459), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n485), .A2(new_n486), .A3(G138), .A4(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n462), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT66), .B1(new_n495), .B2(new_n489), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n485), .A2(G126), .A3(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n488), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n505), .B2(KEYINPUT67), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n509), .A2(new_n511), .B1(new_n501), .B2(new_n502), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  OAI221_X1 g091(.A(new_n506), .B1(new_n507), .B2(new_n513), .C1(new_n514), .C2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND2_X1  g093(.A1(new_n515), .A2(G89), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(new_n522), .B1(new_n503), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n525), .B1(new_n509), .B2(new_n511), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n519), .A2(new_n524), .A3(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  NAND2_X1  g104(.A1(new_n515), .A2(G90), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(G52), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n530), .B(new_n531), .C1(new_n505), .C2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(new_n502), .ZN(new_n539));
  NOR2_X1   g114(.A1(KEYINPUT5), .A2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n526), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n515), .A2(G81), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  AOI22_X1  g128(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n505), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT69), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OR3_X1    g132(.A1(new_n513), .A2(KEYINPUT9), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n513), .B2(new_n557), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n558), .A2(new_n559), .B1(G91), .B2(new_n515), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  NAND2_X1  g137(.A1(new_n515), .A2(G87), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n526), .A2(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  NAND3_X1  g141(.A1(new_n512), .A2(G86), .A3(new_n503), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(KEYINPUT71), .B1(new_n515), .B2(G86), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(G61), .B1(new_n539), .B2(new_n540), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n505), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(KEYINPUT70), .B1(G48), .B2(new_n526), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n574), .A2(KEYINPUT70), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n571), .A2(new_n575), .A3(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(new_n515), .A2(G85), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n526), .A2(G47), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n578), .B(new_n579), .C1(new_n505), .C2(new_n580), .ZN(G290));
  INV_X1    g156(.A(G868), .ZN(new_n582));
  NOR2_X1   g157(.A1(G171), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT72), .ZN(new_n584));
  NAND2_X1  g159(.A1(G79), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G66), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n541), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n513), .A2(KEYINPUT73), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n590));
  OAI21_X1  g165(.A(G54), .B1(new_n526), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n588), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n588), .B(KEYINPUT74), .C1(new_n589), .C2(new_n591), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n515), .A2(G92), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT10), .Z(new_n598));
  AND2_X1   g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n584), .B1(G868), .B2(new_n599), .ZN(G284));
  OAI21_X1  g175(.A(new_n584), .B1(G868), .B2(new_n599), .ZN(G321));
  NOR2_X1   g176(.A1(G286), .A2(new_n582), .ZN(new_n602));
  XOR2_X1   g177(.A(G299), .B(KEYINPUT75), .Z(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n582), .ZN(G297));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n582), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n547), .A2(new_n582), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n596), .A2(new_n598), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n610), .B2(new_n582), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n485), .A2(new_n463), .ZN(new_n613));
  XOR2_X1   g188(.A(KEYINPUT76), .B(KEYINPUT12), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n617), .A2(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n471), .A2(G123), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT77), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(KEYINPUT78), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n621), .A2(KEYINPUT78), .B1(new_n623), .B2(G2105), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n461), .A2(G135), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n617), .A2(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(G2096), .ZN(new_n629));
  NAND4_X1  g204(.A1(new_n618), .A2(new_n627), .A3(new_n628), .A4(new_n629), .ZN(G156));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n636), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  OAI21_X1  g217(.A(G14), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(G401));
  XNOR2_X1  g219(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT17), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT81), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n651), .A2(new_n647), .ZN(new_n654));
  OR3_X1    g229(.A1(new_n654), .A2(KEYINPUT80), .A3(new_n649), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n648), .A2(new_n651), .ZN(new_n656));
  OAI21_X1  g231(.A(KEYINPUT80), .B1(new_n654), .B2(new_n649), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n649), .A2(new_n651), .A3(new_n647), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT79), .B(KEYINPUT18), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n653), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n646), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n645), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT86), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT84), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT19), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n677), .A2(KEYINPUT85), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(KEYINPUT85), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n684), .A2(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(KEYINPUT20), .ZN(new_n686));
  OAI221_X1 g261(.A(new_n681), .B1(new_n680), .B2(new_n676), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n689), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n672), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n687), .A2(new_n689), .ZN(new_n693));
  INV_X1    g268(.A(new_n672), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n687), .A2(new_n689), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n692), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n692), .B2(new_n696), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(G229));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NOR2_X1   g276(.A1(G162), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n701), .B2(G35), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n704));
  INV_X1    g279(.A(G2090), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G5), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G171), .B2(new_n707), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n703), .A2(new_n706), .B1(G1961), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT98), .ZN(new_n711));
  NOR2_X1   g286(.A1(G29), .A2(G33), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT93), .Z(new_n713));
  NAND3_X1  g288(.A1(new_n485), .A2(G139), .A3(new_n462), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT94), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT25), .ZN(new_n717));
  NAND2_X1  g292(.A1(G115), .A2(G2104), .ZN(new_n718));
  INV_X1    g293(.A(G127), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n460), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n717), .B1(G2105), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n715), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n713), .B1(new_n722), .B2(new_n701), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G2072), .Z(new_n724));
  NOR2_X1   g299(.A1(G29), .A2(G32), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n485), .A2(G129), .A3(G2105), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT96), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT26), .Z(new_n729));
  NAND3_X1  g304(.A1(new_n485), .A2(G141), .A3(new_n462), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n463), .A2(G105), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(KEYINPUT97), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT97), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n727), .B2(new_n732), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n725), .B1(new_n737), .B2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(KEYINPUT24), .A2(G34), .ZN(new_n742));
  NOR2_X1   g317(.A1(KEYINPUT24), .A2(G34), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n701), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT95), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G160), .B2(G29), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n724), .B(new_n741), .C1(G2084), .C2(new_n746), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n710), .B1(new_n703), .B2(new_n706), .C1(new_n711), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n711), .ZN(new_n749));
  NOR2_X1   g324(.A1(G4), .A2(G16), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n599), .B2(G16), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(G1348), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(G1348), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n749), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G16), .A2(G21), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G168), .B2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT99), .ZN(new_n757));
  INV_X1    g332(.A(G1966), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n738), .A2(new_n740), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n759), .B(new_n760), .C1(G1961), .C2(new_n709), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n707), .A2(G20), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT23), .Z(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G299), .B2(G16), .ZN(new_n764));
  INV_X1    g339(.A(G1956), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G164), .A2(new_n701), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G27), .B2(new_n701), .ZN(new_n768));
  INV_X1    g343(.A(G2078), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n548), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G16), .B2(G19), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT91), .B(G1341), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n770), .A2(new_n771), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n701), .A2(G26), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT28), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n461), .A2(G140), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n471), .A2(G128), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(G104), .A2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n783), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT92), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(new_n701), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2067), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT31), .B(G11), .Z(new_n789));
  INV_X1    g364(.A(G28), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT30), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n790), .B2(KEYINPUT30), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n793), .B1(new_n626), .B2(new_n701), .C1(G2084), .C2(new_n746), .ZN(new_n794));
  OR4_X1    g369(.A1(new_n766), .A2(new_n777), .A3(new_n788), .A4(new_n794), .ZN(new_n795));
  NOR4_X1   g370(.A1(new_n748), .A2(new_n754), .A3(new_n761), .A4(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n701), .A2(G25), .ZN(new_n798));
  OR2_X1    g373(.A1(G95), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT87), .ZN(new_n801));
  AOI22_X1  g376(.A1(G119), .A2(new_n471), .B1(new_n461), .B2(G131), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n798), .B1(new_n804), .B2(new_n701), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT35), .B(G1991), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT88), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n805), .B(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n707), .A2(G24), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G290), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(G1986), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n808), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n707), .A2(G22), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G166), .B2(new_n707), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1971), .ZN(new_n817));
  MUX2_X1   g392(.A(G6), .B(G305), .S(G16), .Z(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT32), .B(G1981), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT89), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n707), .A2(G23), .ZN(new_n822));
  INV_X1    g397(.A(G288), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n707), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT33), .B(G1976), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n817), .A2(new_n821), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n818), .A2(new_n820), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT90), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n827), .A2(KEYINPUT90), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT34), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n814), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n831), .A2(KEYINPUT34), .A3(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT36), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(new_n839), .A3(new_n836), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n797), .B1(new_n838), .B2(new_n840), .ZN(G311));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n796), .ZN(G150));
  NOR2_X1   g418(.A1(new_n609), .A2(new_n606), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n515), .A2(G93), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n526), .A2(G55), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n846), .B(new_n847), .C1(new_n505), .C2(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n547), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n547), .A2(new_n849), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n845), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n854));
  AOI21_X1  g429(.A(G860), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT101), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n849), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  INV_X1    g435(.A(G160), .ZN(new_n861));
  INV_X1    g436(.A(new_n480), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(new_n478), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n479), .A2(G160), .A3(new_n480), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n863), .B2(new_n864), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n626), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(new_n864), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT102), .ZN(new_n870));
  INV_X1    g445(.A(new_n626), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n461), .A2(G142), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n471), .A2(G130), .ZN(new_n875));
  OR2_X1    g450(.A1(G106), .A2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(new_n615), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n804), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n722), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n734), .B2(new_n736), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n733), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n727), .A2(new_n732), .A3(KEYINPUT105), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n722), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n491), .B1(new_n490), .B2(new_n493), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n495), .A2(new_n489), .A3(KEYINPUT66), .ZN(new_n891));
  OAI211_X1 g466(.A(KEYINPUT103), .B(new_n498), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n488), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT103), .B1(new_n497), .B2(new_n498), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n889), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n498), .B1(new_n890), .B2(new_n891), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n898), .A2(KEYINPUT104), .A3(new_n488), .A4(new_n892), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n895), .A2(new_n786), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n786), .B1(new_n895), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n888), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n883), .B(new_n887), .C1(new_n900), .C2(new_n901), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n868), .A2(new_n873), .B1(new_n881), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n880), .A3(new_n904), .ZN(new_n907));
  AOI21_X1  g482(.A(G37), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n868), .A2(new_n873), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n903), .A2(new_n880), .A3(KEYINPUT106), .A4(new_n904), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n905), .A2(new_n881), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n909), .A2(new_n914), .A3(KEYINPUT107), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT107), .B1(new_n909), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n908), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g494(.A(KEYINPUT108), .B(new_n908), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n919), .A2(KEYINPUT40), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT40), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(G395));
  NAND2_X1  g498(.A1(new_n849), .A2(new_n582), .ZN(new_n924));
  XOR2_X1   g499(.A(G288), .B(KEYINPUT109), .Z(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(G305), .ZN(new_n926));
  XNOR2_X1  g501(.A(G303), .B(G290), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n926), .A2(new_n927), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(KEYINPUT110), .B2(KEYINPUT42), .ZN(new_n932));
  NAND2_X1  g507(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n609), .A2(G299), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n596), .A2(new_n556), .A3(new_n560), .A4(new_n598), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT41), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(KEYINPUT41), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n937), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n610), .B(new_n852), .ZN(new_n944));
  MUX2_X1   g519(.A(new_n942), .B(new_n943), .S(new_n944), .Z(new_n945));
  XNOR2_X1  g520(.A(new_n934), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n924), .B1(new_n946), .B2(new_n582), .ZN(G295));
  OAI21_X1  g522(.A(new_n924), .B1(new_n946), .B2(new_n582), .ZN(G331));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n852), .A2(G171), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n535), .B(new_n536), .C1(new_n850), .C2(new_n851), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(G168), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT112), .B1(new_n953), .B2(new_n941), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n952), .B(G286), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n955), .A2(new_n956), .A3(new_n939), .A4(new_n940), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n953), .A2(new_n943), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n929), .B2(new_n930), .ZN(new_n961));
  INV_X1    g536(.A(new_n930), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(KEYINPUT113), .A3(new_n928), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n959), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n954), .A2(new_n957), .A3(new_n931), .A4(new_n958), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n949), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n958), .B1(new_n941), .B2(new_n953), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n964), .ZN(new_n969));
  INV_X1    g544(.A(G37), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n949), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n975));
  INV_X1    g550(.A(new_n965), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT44), .B1(new_n976), .B2(new_n972), .ZN(new_n977));
  INV_X1    g552(.A(new_n971), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n949), .B1(new_n978), .B2(new_n966), .ZN(new_n979));
  OAI22_X1  g554(.A1(new_n974), .A2(new_n975), .B1(new_n977), .B2(new_n979), .ZN(G397));
  INV_X1    g555(.A(G2067), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n786), .B(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(G1996), .B2(new_n733), .ZN(new_n983));
  INV_X1    g558(.A(G1996), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n737), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n803), .B(new_n807), .Z(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(G290), .B(new_n811), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(KEYINPUT114), .B(G1384), .Z(new_n991));
  NAND3_X1  g566(.A1(new_n895), .A2(new_n899), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n464), .A2(G40), .A3(new_n468), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n990), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G303), .A2(G8), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n893), .B2(new_n894), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT116), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n1001), .C1(new_n893), .C2(new_n894), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(KEYINPUT50), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n499), .A2(new_n1001), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n995), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n705), .A3(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n895), .A2(new_n899), .A3(KEYINPUT45), .A4(new_n991), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n995), .B1(new_n1007), .B2(new_n993), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT115), .B(G1971), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT119), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1011), .A2(new_n1016), .A3(KEYINPUT119), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1000), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT50), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n995), .B1(new_n1007), .B2(KEYINPUT50), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1022), .A2(G2090), .A3(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1026));
  OAI211_X1 g601(.A(G8), .B(new_n1000), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n995), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G288), .A2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1028), .A2(new_n1018), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n503), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1033), .B(new_n567), .C1(new_n1034), .C2(new_n505), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1035), .A2(new_n1036), .A3(G1981), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n1035), .B2(G1981), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n571), .A2(new_n1040), .A3(new_n576), .A4(new_n575), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT49), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1035), .A2(new_n1036), .A3(G1981), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1035), .A2(G1981), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT118), .ZN(new_n1045));
  AND4_X1   g620(.A1(KEYINPUT49), .A2(new_n1041), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1048));
  INV_X1    g623(.A(new_n995), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1018), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1031), .A2(new_n1032), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1030), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(KEYINPUT117), .A3(KEYINPUT52), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1031), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1027), .A2(new_n1051), .A3(new_n1054), .A4(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1003), .A2(new_n993), .A3(new_n1005), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n484), .A2(new_n487), .ZN(new_n1060));
  OAI211_X1 g635(.A(KEYINPUT45), .B(new_n1001), .C1(new_n1060), .C2(new_n896), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n499), .A2(KEYINPUT120), .A3(KEYINPUT45), .A4(new_n1001), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n995), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n758), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1005), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n898), .A2(new_n488), .A3(new_n892), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1004), .B1(new_n1069), .B2(new_n1001), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1009), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G2084), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n1023), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1018), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G168), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1021), .A2(new_n1058), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1024), .B1(new_n1048), .B2(new_n1009), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1077), .A2(new_n1072), .B1(new_n1066), .B2(new_n758), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1078), .A2(new_n1018), .A3(G286), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n705), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1018), .B1(new_n1080), .B2(new_n1016), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1079), .B(KEYINPUT63), .C1(new_n1000), .C2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1076), .A2(KEYINPUT63), .B1(new_n1058), .B2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1051), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1027), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n1029), .A3(new_n823), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1041), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1084), .A2(new_n1085), .B1(new_n1050), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n556), .A2(new_n1091), .A3(new_n560), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1956), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1012), .A2(new_n1013), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1093), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1348), .B1(new_n1071), .B2(new_n1023), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1028), .A2(new_n981), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n599), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1094), .A2(new_n1097), .A3(new_n1093), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1098), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT121), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1105), .B(new_n1098), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G1348), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1028), .A2(new_n981), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1109), .A2(new_n609), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n609), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT60), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1093), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n765), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1117), .B2(new_n1096), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1114), .B1(new_n1118), .B2(new_n1102), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n609), .A2(KEYINPUT60), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1109), .A2(new_n1110), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1096), .A3(new_n1115), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(KEYINPUT61), .A3(new_n1098), .ZN(new_n1123));
  AND4_X1   g698(.A1(new_n1113), .A2(new_n1119), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT58), .B(G1341), .Z(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1028), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1012), .A2(new_n984), .A3(new_n1013), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1128), .B(KEYINPUT122), .C1(new_n1028), .C2(new_n1126), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n548), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT59), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1134), .B(new_n548), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1107), .B1(new_n1124), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G1961), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(G2078), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1059), .A2(new_n1065), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1012), .A2(new_n769), .A3(new_n1013), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1140), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n535), .A2(KEYINPUT54), .A3(new_n536), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n464), .A2(G40), .A3(new_n1141), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n467), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n462), .B1(new_n467), .B2(new_n1152), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1151), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n994), .A2(new_n1012), .A3(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1148), .A2(new_n1139), .A3(new_n1144), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1150), .A2(new_n1157), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1021), .A2(new_n1058), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(G286), .A2(G8), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT123), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(KEYINPUT124), .B(KEYINPUT51), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1162), .B(new_n1163), .C1(new_n1078), .C2(new_n1018), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1161), .B1(new_n1165), .B2(G8), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1022), .A2(G2084), .A3(new_n1024), .ZN(new_n1167));
  AOI21_X1  g742(.A(G1966), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1161), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OR2_X1    g744(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1164), .B1(new_n1166), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT125), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1170), .B(new_n1169), .C1(new_n1074), .C2(new_n1161), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1174), .A2(new_n1175), .A3(new_n1164), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1159), .A2(new_n1173), .A3(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1083), .B(new_n1089), .C1(new_n1137), .C2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1174), .A2(new_n1175), .A3(new_n1164), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1175), .B1(new_n1174), .B2(new_n1164), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1173), .A2(KEYINPUT62), .A3(new_n1176), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1145), .A2(G171), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1021), .A2(new_n1058), .A3(new_n1184), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n997), .B1(new_n1178), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n996), .B1(new_n733), .B2(new_n982), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n996), .A2(new_n984), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1189), .A2(KEYINPUT46), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(KEYINPUT46), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1188), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n1192), .B(KEYINPUT47), .Z(new_n1193));
  INV_X1    g768(.A(new_n996), .ZN(new_n1194));
  OR3_X1    g769(.A1(new_n1194), .A2(G1986), .A3(G290), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT48), .ZN(new_n1196));
  OAI22_X1  g771(.A1(new_n1195), .A2(new_n1196), .B1(new_n988), .B2(new_n1194), .ZN(new_n1197));
  AND2_X1   g772(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1198));
  AND4_X1   g773(.A1(new_n807), .A2(new_n983), .A3(new_n804), .A4(new_n985), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1199), .B1(new_n981), .B2(new_n786), .ZN(new_n1200));
  OAI22_X1  g775(.A1(new_n1197), .A2(new_n1198), .B1(new_n1194), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1193), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1187), .A2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g778(.A1(new_n666), .A2(new_n669), .A3(G319), .ZN(new_n1205));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g781(.A1(new_n666), .A2(new_n669), .A3(KEYINPUT127), .A4(G319), .ZN(new_n1208));
  AOI21_X1  g782(.A(G401), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g783(.A(new_n1209), .B1(new_n698), .B2(new_n699), .ZN(new_n1210));
  INV_X1    g784(.A(new_n1210), .ZN(new_n1211));
  OAI21_X1  g785(.A(new_n1211), .B1(new_n967), .B2(new_n973), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1212), .B1(new_n919), .B2(new_n920), .ZN(G308));
  NAND2_X1  g787(.A1(new_n919), .A2(new_n920), .ZN(new_n1214));
  OAI211_X1 g788(.A(new_n1214), .B(new_n1211), .C1(new_n967), .C2(new_n973), .ZN(G225));
endmodule


