//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1300, new_n1301, new_n1303,
    new_n1304, new_n1305, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(G250), .B1(G257), .B2(G264), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n214));
  AND2_X1   g0014(.A1(KEYINPUT64), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(KEYINPUT64), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n203), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n213), .A2(KEYINPUT0), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n209), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n214), .A2(new_n222), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT65), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n240), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  OAI211_X1 g0052(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  OR2_X1    g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n260), .A2(G223), .B1(new_n263), .B2(G77), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1698), .B1(new_n258), .B2(new_n259), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G222), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n218), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n256), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G226), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT67), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n268), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT69), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n277), .A2(new_n281), .A3(new_n278), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n272), .B1(new_n273), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G150), .ZN(new_n290));
  INV_X1    g0090(.A(new_n216), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT64), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G33), .A3(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT8), .B(G58), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n288), .B(new_n290), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n218), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n299), .A2(new_n207), .A3(G1), .ZN(new_n300));
  INV_X1    g0100(.A(G50), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT70), .B1(new_n207), .B2(G1), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT70), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(new_n206), .A3(G20), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n297), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n299), .A2(G1), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G20), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n298), .B(new_n302), .C1(new_n301), .C2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n287), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT71), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n285), .A2(G179), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n313), .B1(new_n312), .B2(new_n314), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n285), .A2(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n311), .A2(KEYINPUT9), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n311), .A2(KEYINPUT9), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n285), .A2(G200), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT76), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT10), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n325), .A2(KEYINPUT10), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n320), .A2(new_n321), .B1(new_n285), .B2(G200), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n329), .A2(new_n325), .A3(KEYINPUT10), .A4(new_n319), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n300), .A2(new_n224), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n310), .B2(new_n224), .ZN(new_n333));
  INV_X1    g0133(.A(new_n294), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT64), .B(G20), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(new_n289), .B1(new_n335), .B2(G77), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT15), .B(G87), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n338), .A2(KEYINPUT74), .A3(G33), .A4(new_n217), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT74), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n293), .B2(new_n337), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n333), .B1(new_n342), .B2(new_n297), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT72), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n265), .A2(new_n345), .A3(G232), .ZN(new_n346));
  OAI211_X1 g0146(.A(G232), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT72), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(G238), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT3), .B(G33), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT73), .B(G107), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n270), .B1(new_n349), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n225), .B1(new_n280), .B2(new_n282), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n355), .A2(new_n356), .A3(new_n256), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n344), .B1(new_n357), .B2(G190), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n277), .A2(new_n281), .A3(new_n278), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n281), .B1(new_n277), .B2(new_n278), .ZN(new_n360));
  OAI21_X1  g0160(.A(G244), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n353), .B1(new_n346), .B2(new_n348), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n255), .C1(new_n362), .C2(new_n270), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G200), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n317), .A2(new_n331), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT17), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n201), .A2(new_n202), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G58), .A2(G68), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n289), .A2(G159), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT7), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n217), .A2(new_n263), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n258), .A2(new_n207), .A3(new_n259), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n202), .B1(new_n375), .B2(KEYINPUT7), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n372), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n307), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n373), .B1(new_n217), .B2(new_n263), .ZN(new_n380));
  NOR4_X1   g0180(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT7), .A4(G20), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n380), .A2(new_n381), .A3(new_n202), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n379), .B1(new_n382), .B2(new_n372), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n310), .A2(new_n334), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n309), .A2(new_n294), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n277), .A2(G232), .A3(new_n278), .ZN(new_n389));
  INV_X1    g0189(.A(G33), .ZN(new_n390));
  INV_X1    g0190(.A(G87), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G223), .A2(G1698), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n273), .B2(G1698), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n392), .B1(new_n394), .B2(new_n351), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n255), .B(new_n389), .C1(new_n395), .C2(new_n270), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G200), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n318), .B2(new_n396), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n367), .B1(new_n388), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n398), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n378), .A2(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT17), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n273), .A2(G1698), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n405), .B1(G223), .B2(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n271), .B1(new_n407), .B2(new_n392), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n408), .A2(G179), .A3(new_n255), .A4(new_n389), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n396), .A2(G169), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n404), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT83), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT83), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n404), .C1(new_n401), .C2(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n411), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n388), .A3(KEYINPUT18), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n403), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G179), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n357), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n343), .B1(new_n363), .B2(new_n286), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(KEYINPUT75), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT75), .ZN(new_n424));
  AOI211_X1 g0224(.A(new_n424), .B(new_n343), .C1(new_n363), .C2(new_n286), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n366), .A2(new_n419), .A3(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n293), .B2(new_n224), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n297), .ZN(new_n431));
  XOR2_X1   g0231(.A(new_n431), .B(KEYINPUT11), .Z(new_n432));
  INV_X1    g0232(.A(KEYINPUT79), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n300), .A2(new_n202), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(KEYINPUT80), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT12), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT79), .B1(new_n300), .B2(new_n202), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n437), .A2(KEYINPUT12), .ZN(new_n438));
  OAI221_X1 g0238(.A(new_n436), .B1(new_n202), .B2(new_n310), .C1(new_n438), .C2(new_n435), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n283), .A2(G238), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n255), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT77), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n351), .A2(G1698), .ZN(new_n444));
  INV_X1    g0244(.A(G232), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n260), .A2(KEYINPUT77), .A3(G232), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT78), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(G33), .A3(G97), .ZN(new_n450));
  INV_X1    g0250(.A(G97), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT78), .B1(new_n390), .B2(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n265), .A2(G226), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n270), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT13), .B1(new_n442), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n448), .A2(new_n453), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n271), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT13), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n256), .B1(new_n283), .B2(G238), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n440), .B1(new_n461), .B2(new_n318), .ZN(new_n462));
  INV_X1    g0262(.A(G200), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n455), .B2(new_n460), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n455), .A2(G179), .A3(new_n460), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT14), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT81), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n442), .A2(KEYINPUT13), .A3(new_n454), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n458), .B1(new_n457), .B2(new_n459), .ZN(new_n471));
  OAI21_X1  g0271(.A(G169), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n467), .A2(KEYINPUT81), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n461), .A2(G169), .A3(new_n473), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n469), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OR3_X1    g0277(.A1(new_n432), .A2(new_n439), .A3(KEYINPUT82), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT82), .B1(new_n432), .B2(new_n439), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n465), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n428), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(KEYINPUT23), .A2(G107), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n215), .B2(new_n216), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT91), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT91), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n335), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n391), .A2(KEYINPUT90), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n217), .A2(new_n351), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n488), .B1(new_n491), .B2(KEYINPUT22), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT23), .ZN(new_n493));
  OAI21_X1  g0293(.A(G20), .B1(new_n352), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G116), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n390), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n217), .A2(new_n351), .A3(KEYINPUT22), .A4(new_n489), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n492), .A2(new_n499), .A3(KEYINPUT24), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT24), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n491), .A2(KEYINPUT22), .B1(new_n494), .B2(new_n496), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT22), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n485), .A2(new_n487), .B1(new_n490), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n501), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n297), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n307), .B(new_n309), .C1(G1), .C2(new_n390), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n300), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT25), .B1(new_n300), .B2(new_n226), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n507), .A2(new_n226), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(G250), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n513));
  OAI211_X1 g0313(.A(G257), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n514));
  INV_X1    g0314(.A(G294), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n514), .C1(new_n390), .C2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n218), .B1(new_n274), .B2(new_n269), .ZN(new_n517));
  XNOR2_X1  g0317(.A(KEYINPUT5), .B(G41), .ZN(new_n518));
  INV_X1    g0318(.A(G45), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G1), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n276), .A2(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n516), .A2(new_n271), .B1(new_n521), .B2(G264), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n277), .A2(G274), .A3(new_n520), .A4(new_n518), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(G190), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n516), .A2(new_n271), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n521), .A2(G264), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G200), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n506), .A2(new_n512), .A3(new_n524), .A4(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(G169), .B1(new_n522), .B2(new_n523), .ZN(new_n530));
  AND4_X1   g0330(.A1(new_n420), .A2(new_n525), .A3(new_n523), .A4(new_n526), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT24), .B1(new_n492), .B2(new_n499), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n502), .A2(new_n504), .A3(new_n501), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n307), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n532), .B1(new_n535), .B2(new_n511), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G87), .A2(G97), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n352), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n352), .A2(KEYINPUT87), .A3(new_n537), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n452), .A2(new_n450), .A3(KEYINPUT19), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n540), .A2(new_n541), .B1(new_n217), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n263), .A2(new_n335), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G68), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n217), .A2(G33), .A3(G97), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n297), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n337), .A2(new_n300), .ZN(new_n551));
  INV_X1    g0351(.A(new_n507), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n338), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n351), .A2(G238), .A3(new_n257), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT86), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n265), .A2(KEYINPUT86), .A3(G238), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n260), .A2(G244), .B1(G33), .B2(G116), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n270), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n277), .B(G250), .C1(G1), .C2(new_n519), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n520), .A2(G274), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n286), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n564), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n444), .A2(new_n225), .B1(new_n390), .B2(new_n495), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n557), .B2(new_n558), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n420), .B(new_n566), .C1(new_n568), .C2(new_n270), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n554), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(G200), .B1(new_n561), .B2(new_n564), .ZN(new_n571));
  OAI211_X1 g0371(.A(G190), .B(new_n566), .C1(new_n568), .C2(new_n270), .ZN(new_n572));
  AOI22_X1  g0372(.A1(G68), .A2(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n542), .A2(new_n217), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n352), .A2(KEYINPUT87), .A3(new_n537), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT87), .B1(new_n352), .B2(new_n537), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n297), .B1(new_n300), .B2(new_n337), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n552), .A2(G87), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n571), .A2(new_n572), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n529), .A2(new_n536), .A3(new_n570), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n300), .A2(new_n495), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n507), .B2(new_n495), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT89), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G283), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n390), .A2(G97), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n217), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n587), .B1(new_n451), .B2(G33), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT89), .B1(new_n335), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n297), .B1(new_n207), .B2(G116), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT20), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT20), .ZN(new_n596));
  AOI211_X1 g0396(.A(new_n596), .B(new_n593), .C1(new_n589), .C2(new_n591), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n585), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n518), .A2(new_n520), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(G270), .A3(new_n277), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n600), .A2(new_n523), .ZN(new_n601));
  OAI211_X1 g0401(.A(G257), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n258), .A2(G303), .A3(new_n259), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(G264), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT88), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n605), .A2(new_n602), .A3(KEYINPUT88), .A4(new_n603), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n271), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n601), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n598), .A2(G169), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n598), .A2(KEYINPUT21), .A3(G169), .A4(new_n609), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n609), .A2(new_n420), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n598), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n609), .A2(G200), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n592), .A2(new_n594), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n596), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n594), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n584), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n601), .B(G190), .C1(new_n606), .C2(new_n608), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n616), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n612), .A2(new_n613), .A3(new_n615), .A4(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(G244), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT4), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n351), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n351), .A2(G250), .A3(G1698), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n587), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n271), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n599), .A2(G257), .A3(new_n277), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n523), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n286), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n632), .B1(new_n271), .B2(new_n629), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n420), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n380), .A2(new_n381), .A3(new_n352), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n289), .A2(KEYINPUT84), .A3(G77), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT84), .B1(new_n289), .B2(G77), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g0441(.A(G97), .B(G107), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT6), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(new_n451), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n642), .A2(new_n643), .B1(new_n226), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n641), .B1(new_n645), .B2(new_n217), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n297), .B1(new_n638), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n300), .A2(new_n451), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n507), .B2(new_n451), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n635), .A2(new_n637), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(G97), .A2(G107), .ZN(new_n653));
  NOR2_X1   g0453(.A1(G97), .A2(G107), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n643), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n226), .A2(KEYINPUT6), .A3(G97), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n217), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n289), .A2(G77), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT84), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n289), .A2(KEYINPUT84), .A3(G77), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT7), .B1(new_n335), .B2(new_n351), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n263), .A2(new_n373), .A3(new_n207), .ZN(new_n665));
  INV_X1    g0465(.A(new_n352), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n649), .B1(new_n668), .B2(new_n297), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n630), .A2(new_n633), .A3(G190), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n669), .B(new_n670), .C1(new_n463), .C2(new_n636), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n652), .A2(new_n671), .A3(KEYINPUT85), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT85), .B1(new_n652), .B2(new_n671), .ZN(new_n673));
  NOR4_X1   g0473(.A1(new_n582), .A2(new_n623), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n482), .A2(new_n674), .ZN(G372));
  NAND2_X1  g0475(.A1(new_n418), .A2(new_n412), .ZN(new_n676));
  INV_X1    g0476(.A(new_n477), .ZN(new_n677));
  INV_X1    g0477(.A(new_n480), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n677), .A2(new_n678), .B1(new_n465), .B2(new_n426), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n676), .B1(new_n679), .B2(new_n403), .ZN(new_n680));
  INV_X1    g0480(.A(new_n331), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n317), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n482), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n581), .A2(new_n570), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n528), .A2(new_n524), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n535), .A2(new_n686), .A3(new_n511), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n652), .A2(new_n671), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n615), .A2(new_n613), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n612), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n527), .A2(new_n286), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n522), .A2(new_n420), .A3(new_n523), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n506), .B2(new_n512), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n685), .B(new_n689), .C1(new_n691), .C2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT26), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n684), .B2(new_n652), .ZN(new_n698));
  INV_X1    g0498(.A(new_n652), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n581), .A3(new_n570), .A4(KEYINPUT26), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n570), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n682), .B1(new_n683), .B2(new_n703), .ZN(G369));
  NAND2_X1  g0504(.A1(new_n217), .A2(new_n308), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G213), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n620), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n691), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n623), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n536), .A2(new_n710), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n535), .A2(new_n511), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n529), .B1(new_n717), .B2(new_n711), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n716), .B1(new_n718), .B2(new_n536), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n536), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n710), .B1(new_n690), .B2(new_n612), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n716), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(new_n725), .ZN(G399));
  NOR2_X1   g0526(.A1(new_n211), .A2(G41), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n540), .A2(new_n495), .A3(new_n541), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n727), .A2(new_n728), .A3(new_n206), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n221), .B2(new_n727), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  NAND2_X1  g0531(.A1(new_n702), .A2(new_n711), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT93), .B1(new_n733), .B2(KEYINPUT29), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n698), .A2(KEYINPUT94), .A3(new_n700), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n700), .A2(KEYINPUT94), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n696), .A2(new_n735), .A3(new_n570), .A4(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n737), .A2(new_n711), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT29), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT93), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT29), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n732), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n734), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n674), .B2(new_n711), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n566), .B1(new_n568), .B2(new_n270), .ZN(new_n746));
  INV_X1    g0546(.A(new_n522), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n746), .A2(new_n634), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n614), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(KEYINPUT30), .A3(new_n614), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n636), .A2(G179), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(new_n609), .A3(new_n746), .A4(new_n527), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n710), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n745), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n751), .A2(new_n754), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT92), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n751), .A2(KEYINPUT92), .A3(new_n754), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n761), .A2(new_n752), .A3(new_n762), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n764));
  OAI21_X1  g0564(.A(G330), .B1(new_n758), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n743), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n731), .B1(new_n767), .B2(G1), .ZN(G364));
  NOR2_X1   g0568(.A1(new_n335), .A2(new_n299), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G45), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G1), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n727), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n714), .B2(G330), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G330), .B2(new_n714), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n211), .A2(new_n263), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G355), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G116), .B2(new_n210), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n211), .A2(new_n351), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n519), .B2(new_n221), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n248), .A2(new_n519), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n218), .B1(G20), .B2(new_n286), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT95), .Z(new_n788));
  OAI21_X1  g0588(.A(new_n772), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n335), .A2(G179), .A3(G200), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n790), .A2(KEYINPUT97), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(KEYINPUT97), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n791), .A2(G190), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n791), .A2(new_n318), .A3(new_n792), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G326), .A2(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n217), .A2(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G179), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT98), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT98), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G329), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n463), .A2(G179), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n799), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n420), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n799), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n807), .A2(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n808), .A2(G20), .A3(G190), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT101), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n813), .B1(G303), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n217), .B1(G190), .B2(new_n800), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n263), .B1(new_n817), .B2(new_n515), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n335), .A2(G190), .A3(new_n810), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(KEYINPUT96), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n819), .A2(KEYINPUT96), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n818), .B1(new_n823), .B2(G322), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n798), .A2(new_n806), .A3(new_n816), .A4(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G159), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n804), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n814), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n263), .B1(new_n830), .B2(G87), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n831), .B1(new_n811), .B2(new_n224), .C1(new_n226), .C2(new_n809), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G58), .B2(new_n823), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n829), .B(new_n833), .C1(new_n301), .C2(new_n793), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n817), .A2(new_n451), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n796), .B2(G68), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT100), .Z(new_n837));
  OAI21_X1  g0637(.A(new_n825), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n789), .B1(new_n838), .B2(new_n786), .ZN(new_n839));
  INV_X1    g0639(.A(new_n785), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n714), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n774), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  INV_X1    g0643(.A(KEYINPUT103), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n423), .B2(new_n425), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n349), .A2(new_n354), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n256), .B1(new_n846), .B2(new_n271), .ZN(new_n847));
  AOI21_X1  g0647(.A(G169), .B1(new_n847), .B2(new_n361), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n424), .B1(new_n848), .B2(new_n343), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(new_n850), .A3(KEYINPUT103), .A4(new_n421), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n711), .A2(new_n343), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n358), .B2(new_n364), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n845), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT104), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n845), .A2(new_n851), .A3(KEYINPUT104), .A4(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n426), .A2(new_n852), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT105), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n854), .A2(new_n855), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT105), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n861), .A2(new_n862), .A3(new_n857), .A4(new_n858), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n732), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n733), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n772), .B1(new_n868), .B2(new_n765), .ZN(new_n869));
  INV_X1    g0669(.A(G330), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n687), .A2(new_n695), .ZN(new_n871));
  INV_X1    g0671(.A(new_n673), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n652), .A2(new_n671), .A3(KEYINPUT85), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n871), .A2(new_n872), .A3(new_n685), .A4(new_n873), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n874), .A2(new_n623), .A3(new_n710), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n756), .B1(new_n875), .B2(new_n744), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n870), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n866), .A2(new_n878), .A3(new_n867), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n869), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n786), .A2(new_n783), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n772), .B1(G77), .B2(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n805), .A2(G311), .B1(G303), .B2(new_n794), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n811), .A2(new_n495), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n809), .A2(new_n391), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n885), .B(new_n886), .C1(G107), .C2(new_n815), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n351), .B(new_n835), .C1(new_n823), .C2(G294), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n796), .A2(G283), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n884), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n811), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n823), .A2(G143), .B1(G159), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(G137), .ZN(new_n893));
  INV_X1    g0693(.A(G150), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n892), .B1(new_n893), .B2(new_n793), .C1(new_n894), .C2(new_n795), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT102), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT34), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n815), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n899), .A2(new_n301), .B1(new_n201), .B2(new_n817), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n809), .A2(new_n202), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n900), .A2(new_n263), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(G132), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n898), .B(new_n902), .C1(new_n903), .C2(new_n804), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n896), .A2(new_n897), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n890), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n883), .B1(new_n906), .B2(new_n786), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n864), .B2(new_n784), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT106), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n880), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(G384));
  INV_X1    g0711(.A(new_n645), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n912), .A2(KEYINPUT35), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(KEYINPUT35), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n913), .A2(new_n914), .A3(G116), .A4(new_n219), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT36), .Z(new_n916));
  OR3_X1    g0716(.A1(new_n220), .A2(new_n224), .A3(new_n368), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n301), .A2(G68), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n206), .B(G13), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n708), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n676), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n417), .A2(new_n388), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n388), .A2(new_n921), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n400), .A2(new_n401), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT37), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n923), .A2(new_n924), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n378), .B1(KEYINPUT16), .B2(new_n377), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n387), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n417), .B2(new_n921), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n930), .A2(new_n925), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n927), .B1(new_n931), .B2(new_n926), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(new_n921), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n932), .B1(new_n419), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT38), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n932), .B(KEYINPUT38), .C1(new_n419), .C2(new_n933), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n936), .A2(KEYINPUT39), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT108), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n403), .A2(new_n939), .B1(new_n418), .B2(new_n412), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n399), .A2(KEYINPUT108), .A3(new_n402), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n924), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT37), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n944), .A2(new_n927), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n935), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT39), .B1(new_n946), .B2(new_n937), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n938), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n677), .A2(new_n678), .A3(new_n711), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n922), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n845), .A2(new_n851), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n711), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n867), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n936), .A2(new_n937), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT107), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n465), .B(new_n956), .C1(new_n477), .C2(new_n480), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n478), .A2(new_n479), .A3(new_n710), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n465), .A2(new_n477), .A3(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n465), .B(KEYINPUT107), .C1(new_n477), .C2(new_n480), .ZN(new_n960));
  INV_X1    g0760(.A(new_n958), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n957), .A2(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n954), .A2(new_n955), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n951), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n734), .A2(new_n482), .A3(new_n739), .A4(new_n742), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n682), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n757), .A2(KEYINPUT31), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n745), .B2(new_n757), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n403), .A2(new_n939), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(new_n676), .A3(new_n941), .ZN(new_n972));
  INV_X1    g0772(.A(new_n924), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n972), .A2(new_n973), .B1(new_n927), .B2(new_n944), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n937), .B1(new_n974), .B2(KEYINPUT38), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n864), .A2(new_n970), .A3(new_n962), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT40), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT40), .B1(new_n936), .B2(new_n937), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n978), .A2(new_n864), .A3(new_n962), .A4(new_n970), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n482), .A2(new_n970), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n980), .A2(new_n981), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n983), .A2(new_n984), .A3(new_n870), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n968), .A2(new_n985), .B1(new_n206), .B2(new_n769), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n968), .A2(new_n985), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n920), .B1(new_n986), .B2(new_n987), .ZN(G367));
  AOI21_X1  g0788(.A(new_n711), .B1(new_n579), .B2(new_n580), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT109), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n685), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n570), .B2(new_n990), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT110), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT43), .B1(new_n992), .B2(new_n993), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(KEYINPUT43), .B2(new_n992), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n719), .A2(new_n724), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n699), .A2(new_n710), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n652), .B(new_n671), .C1(new_n669), .C2(new_n711), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT112), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(KEYINPUT112), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1003), .A2(KEYINPUT42), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n652), .B1(new_n1000), .B2(new_n536), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT111), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n711), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(KEYINPUT42), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n997), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1012), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1014), .A2(new_n996), .A3(new_n1005), .A4(new_n1010), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1001), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n722), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1013), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n727), .B(KEYINPUT41), .Z(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n719), .A2(new_n724), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n998), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(new_n715), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n743), .A2(new_n765), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT115), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n743), .A2(new_n1027), .A3(KEYINPUT115), .A4(new_n765), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n725), .A2(new_n1001), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT45), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT44), .ZN(new_n1035));
  OR3_X1    g0835(.A1(new_n725), .A2(new_n1035), .A3(new_n1001), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n725), .B2(new_n1001), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(KEYINPUT113), .B1(new_n722), .B2(KEYINPUT114), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(KEYINPUT114), .B1(new_n1039), .B2(KEYINPUT113), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n721), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1030), .A2(new_n1031), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1024), .B1(new_n1045), .B2(new_n766), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n771), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1022), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n992), .A2(new_n840), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n788), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n210), .B2(new_n337), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n244), .A2(new_n779), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n772), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G294), .A2(new_n796), .B1(new_n794), .B2(G311), .ZN(new_n1054));
  INV_X1    g0854(.A(G317), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n804), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n823), .A2(G303), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT46), .B1(new_n830), .B2(G116), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n351), .B(new_n1058), .C1(G283), .C2(new_n891), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n815), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n809), .A2(new_n451), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n817), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1061), .B1(new_n666), .B2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n794), .A2(G143), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n826), .B2(new_n795), .C1(new_n804), .C2(new_n893), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n351), .B1(new_n814), .B2(new_n201), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n809), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(G77), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n817), .A2(new_n202), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G50), .B2(new_n891), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n823), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1069), .B(new_n1071), .C1(new_n1072), .C2(new_n894), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1056), .A2(new_n1064), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT47), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1053), .B1(new_n1075), .B2(new_n786), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1049), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1048), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(G387));
  NOR2_X1   g0880(.A1(new_n814), .A2(new_n224), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1061), .A2(new_n263), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1062), .A2(new_n338), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(new_n202), .C2(new_n811), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G50), .B2(new_n823), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n805), .A2(G150), .B1(new_n334), .B2(new_n796), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n826), .C2(new_n793), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n805), .A2(G326), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n351), .B1(new_n1068), .B2(G116), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n823), .A2(G317), .B1(G303), .B2(new_n891), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n794), .A2(G322), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n812), .C2(new_n795), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT48), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1062), .A2(G283), .B1(new_n830), .B2(G294), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT49), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1088), .B(new_n1089), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1087), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n786), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n772), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n719), .A2(new_n840), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n779), .B1(new_n240), .B2(G45), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n728), .B2(new_n775), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n294), .A2(G50), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT50), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n519), .B1(new_n202), .B2(new_n224), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n728), .B(new_n1109), .C1(new_n1108), .C2(new_n1107), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1106), .A2(new_n1110), .B1(G107), .B2(new_n210), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1103), .B(new_n1104), .C1(new_n1050), .C2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1027), .A2(new_n771), .B1(new_n1102), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n767), .A2(new_n1027), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1028), .A2(new_n727), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(G393));
  OAI221_X1 g0916(.A(new_n263), .B1(new_n807), .B2(new_n814), .C1(new_n809), .C2(new_n226), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n805), .B2(G322), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1072), .A2(new_n812), .B1(new_n1055), .B2(new_n793), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT52), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n796), .A2(G303), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n891), .A2(G294), .B1(new_n1062), .B2(G116), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1072), .A2(new_n826), .B1(new_n894), .B2(new_n793), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT51), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n891), .A2(new_n334), .B1(new_n1062), .B2(G77), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n301), .B2(new_n795), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT116), .Z(new_n1129));
  OAI21_X1  g0929(.A(new_n351), .B1(new_n814), .B2(new_n202), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n886), .B(new_n1130), .C1(new_n805), .C2(G143), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1126), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1124), .B1(new_n1133), .B2(KEYINPUT117), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n786), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n788), .B1(G97), .B2(new_n211), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n778), .A2(new_n251), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1103), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1137), .B(new_n1140), .C1(new_n840), .C2(new_n1001), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1039), .B(new_n721), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n1047), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n727), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n1142), .B2(new_n1028), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1143), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(G390));
  AOI21_X1  g0950(.A(new_n732), .B1(new_n860), .B2(new_n863), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n953), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n962), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n949), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n948), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n878), .A2(new_n864), .A3(new_n962), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1152), .B1(new_n864), .B2(new_n738), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n962), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n949), .B(new_n975), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1156), .A2(new_n1157), .A3(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n864), .A2(new_n970), .A3(G330), .A4(new_n962), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n948), .B1(new_n1153), .B2(new_n949), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n975), .A2(new_n949), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n859), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n862), .B1(new_n1166), .B2(new_n861), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n863), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n738), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n953), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1165), .B1(new_n1170), .B2(new_n962), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1163), .B1(new_n1164), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1161), .A2(new_n1172), .A3(new_n771), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT119), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT119), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1161), .A2(new_n1172), .A3(new_n1175), .A4(new_n771), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n482), .A2(new_n970), .A3(G330), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n965), .A2(new_n682), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n864), .A2(new_n970), .A3(G330), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1159), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1159), .B1(new_n765), .B2(new_n865), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1186), .B2(new_n1162), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1180), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1162), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1157), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1164), .A2(new_n1171), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1188), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n962), .B1(new_n878), .B2(new_n864), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n954), .B1(new_n1163), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1179), .B1(new_n1194), .B2(new_n1183), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(new_n1161), .A3(new_n1172), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1192), .A2(new_n727), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n772), .B1(new_n334), .B2(new_n882), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n351), .B(new_n901), .C1(new_n823), .C2(G116), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n891), .A2(G97), .B1(new_n1062), .B2(G77), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n391), .C2(new_n899), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n805), .A2(G294), .B1(new_n666), .B2(new_n796), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n807), .B2(new_n793), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n805), .A2(G125), .B1(G128), .B2(new_n794), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n893), .B2(new_n795), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n823), .A2(G132), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(KEYINPUT54), .B(G143), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT120), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n891), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n830), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT53), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n814), .B2(new_n894), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1068), .A2(G50), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n263), .B1(new_n1062), .B2(G159), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1206), .A2(new_n1209), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n1201), .A2(new_n1203), .B1(new_n1205), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1198), .B1(new_n1216), .B2(new_n786), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n948), .B2(new_n784), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1177), .A2(new_n1197), .A3(new_n1218), .ZN(G378));
  OAI21_X1  g1019(.A(new_n772), .B1(G50), .B2(new_n882), .ZN(new_n1220));
  INV_X1    g1020(.A(G41), .ZN(new_n1221));
  AOI21_X1  g1021(.A(G50), .B1(new_n259), .B2(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n804), .A2(new_n807), .B1(new_n495), .B2(new_n793), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1070), .A2(G41), .A3(new_n351), .A4(new_n1081), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G58), .A2(new_n1068), .B1(new_n891), .B2(new_n338), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n1072), .C2(new_n226), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1223), .B(new_n1226), .C1(G97), .C2(new_n796), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT121), .Z(new_n1228));
  INV_X1    g1028(.A(KEYINPUT58), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1222), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n795), .A2(new_n903), .B1(new_n893), .B2(new_n811), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT122), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n794), .A2(G125), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n823), .A2(G128), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G150), .A2(new_n1062), .B1(new_n1208), .B2(new_n830), .ZN(new_n1235));
  AND4_X1   g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n390), .B(new_n1221), .C1(new_n809), .C2(new_n826), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n805), .B2(G124), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT59), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1240), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1230), .B1(new_n1229), .B2(new_n1228), .C1(new_n1238), .C2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1220), .B1(new_n1243), .B2(new_n786), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n312), .A2(new_n314), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n311), .A2(new_n921), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  OR3_X1    g1047(.A1(new_n331), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n331), .B2(new_n1245), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n783), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1244), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1253), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n980), .B2(G330), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n870), .B(new_n1253), .C1(new_n977), .C2(new_n979), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n964), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n864), .A2(new_n962), .A3(new_n970), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1261), .A2(new_n978), .B1(new_n976), .B2(KEYINPUT40), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1253), .B1(new_n1262), .B2(new_n870), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n951), .A2(new_n963), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n980), .A2(G330), .A3(new_n1257), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1260), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1256), .B1(new_n1267), .B2(new_n771), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1196), .A2(new_n1180), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1267), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT57), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1147), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1180), .A2(new_n1196), .B1(new_n1260), .B2(new_n1266), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT57), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1269), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(G375));
  OAI21_X1  g1077(.A(new_n771), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1103), .B1(new_n202), .B2(new_n881), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n786), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n899), .A2(new_n826), .B1(new_n894), .B2(new_n811), .ZN(new_n1281));
  OAI221_X1 g1081(.A(new_n351), .B1(new_n201), .B2(new_n809), .C1(new_n1072), .C2(new_n893), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n1281), .B(new_n1282), .C1(G50), .C2(new_n1062), .ZN(new_n1283));
  INV_X1    g1083(.A(G128), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n804), .A2(new_n1284), .B1(new_n903), .B2(new_n793), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n796), .B2(new_n1208), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n263), .B1(new_n809), .B2(new_n224), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1083), .B1(new_n811), .B2(new_n352), .C1(new_n899), .C2(new_n451), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1287), .B(new_n1288), .C1(G283), .C2(new_n823), .ZN(new_n1289));
  INV_X1    g1089(.A(G303), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n804), .A2(new_n1290), .B1(new_n495), .B2(new_n795), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(G294), .B2(new_n794), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1283), .A2(new_n1286), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1293));
  OAI221_X1 g1093(.A(new_n1279), .B1(new_n1280), .B2(new_n1293), .C1(new_n962), .C2(new_n784), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1278), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1194), .A2(new_n1179), .A3(new_n1183), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1195), .A2(new_n1023), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(G381));
  NOR2_X1   g1099(.A1(G375), .A2(G378), .ZN(new_n1300));
  NOR4_X1   g1100(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1300), .A2(new_n1079), .A3(new_n1298), .A4(new_n1301), .ZN(G407));
  INV_X1    g1102(.A(G213), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1303), .A2(G343), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(G407), .A2(G213), .A3(new_n1305), .ZN(G409));
  INV_X1    g1106(.A(new_n1295), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1188), .A2(KEYINPUT60), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1308), .A2(new_n1296), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1194), .A2(KEYINPUT60), .A3(new_n1179), .A4(new_n1183), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n727), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G384), .B(new_n1307), .C1(new_n1309), .C2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1311), .B1(new_n1308), .B2(new_n1296), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n910), .B1(new_n1313), .B2(new_n1295), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1304), .A2(G2897), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1312), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n727), .B1(new_n1274), .B2(KEYINPUT57), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1270), .A2(new_n1267), .A3(KEYINPUT57), .ZN(new_n1320));
  OAI211_X1 g1120(.A(G378), .B(new_n1268), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1177), .A2(new_n1197), .A3(new_n1218), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1260), .A2(KEYINPUT123), .A3(new_n1266), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT123), .B1(new_n1260), .B2(new_n1266), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1323), .A2(new_n1324), .A3(new_n1047), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1270), .A2(new_n1267), .A3(new_n1024), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1255), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1322), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1304), .B1(new_n1321), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT124), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1318), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1256), .B1(new_n1274), .B2(new_n1024), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT123), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1267), .A2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1260), .A2(new_n1266), .A3(KEYINPUT123), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n771), .A3(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G378), .B1(new_n1332), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1337), .B1(G378), .B2(new_n1276), .ZN(new_n1338));
  OAI21_X1  g1138(.A(KEYINPUT124), .B1(new_n1338), .B2(new_n1304), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1331), .A2(new_n1339), .ZN(new_n1340));
  AND2_X1   g1140(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1329), .A2(KEYINPUT63), .A3(new_n1341), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(G393), .B(new_n842), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1023), .B1(new_n1146), .B2(new_n767), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1020), .B(new_n1021), .C1(new_n1345), .C2(new_n771), .ZN(new_n1346));
  AOI21_X1  g1146(.A(G390), .B1(new_n1346), .B2(new_n1077), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1048), .A2(new_n1078), .A3(new_n1149), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1344), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT61), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1346), .A2(new_n1077), .A3(G390), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1149), .B1(new_n1048), .B2(new_n1078), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1351), .A2(new_n1352), .A3(new_n1343), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1349), .A2(new_n1350), .A3(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1321), .A2(new_n1328), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1304), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1355), .A2(new_n1356), .A3(new_n1341), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT63), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1354), .B1(new_n1357), .B2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1340), .A2(new_n1342), .A3(new_n1359), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1357), .A2(KEYINPUT62), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1350), .B1(new_n1329), .B2(new_n1318), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT62), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1363), .B1(new_n1329), .B2(new_n1341), .ZN(new_n1364));
  NOR3_X1   g1164(.A1(new_n1361), .A2(new_n1362), .A3(new_n1364), .ZN(new_n1365));
  AND2_X1   g1165(.A1(new_n1349), .A2(new_n1353), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1360), .B1(new_n1365), .B2(new_n1366), .ZN(G405));
  INV_X1    g1167(.A(KEYINPUT125), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT126), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1312), .A2(new_n1369), .A3(new_n1314), .ZN(new_n1370));
  AND3_X1   g1170(.A1(new_n1321), .A2(new_n1368), .A3(new_n1370), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1370), .B1(new_n1321), .B2(new_n1368), .ZN(new_n1372));
  OAI211_X1 g1172(.A(new_n1322), .B(G375), .C1(new_n1371), .C2(new_n1372), .ZN(new_n1373));
  INV_X1    g1173(.A(new_n1372), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1321), .A2(new_n1368), .A3(new_n1370), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(G375), .A2(new_n1322), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1374), .A2(new_n1375), .A3(new_n1376), .ZN(new_n1377));
  AND3_X1   g1177(.A1(new_n1373), .A2(new_n1377), .A3(new_n1366), .ZN(new_n1378));
  AOI21_X1  g1178(.A(new_n1366), .B1(new_n1373), .B2(new_n1377), .ZN(new_n1379));
  NOR2_X1   g1179(.A1(new_n1378), .A2(new_n1379), .ZN(G402));
endmodule


