//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT65), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  AOI22_X1  g031(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(G125), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(new_n465), .A3(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n458), .A2(new_n459), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n464), .A2(new_n466), .B1(new_n467), .B2(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n469), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n467), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  OAI211_X1 g055(.A(G138), .B(new_n467), .C1(new_n458), .C2(new_n459), .ZN(new_n481));
  OAI21_X1  g056(.A(G126), .B1(new_n458), .B2(new_n459), .ZN(new_n482));
  NAND2_X1  g057(.A1(G114), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n467), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(KEYINPUT4), .B(G138), .C1(new_n458), .C2(new_n459), .ZN(new_n487));
  NAND2_X1  g062(.A1(G102), .A2(G2104), .ZN(new_n488));
  AOI21_X1  g063(.A(G2105), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n486), .A2(KEYINPUT68), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(KEYINPUT68), .B1(new_n486), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(G164));
  NAND2_X1  g068(.A1(G75), .A2(G543), .ZN(new_n494));
  XOR2_X1   g069(.A(KEYINPUT5), .B(G543), .Z(new_n495));
  INV_X1    g070(.A(G62), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(G50), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G88), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G166));
  NAND2_X1  g080(.A1(G76), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT7), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(G63), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT6), .B(G651), .Z(new_n513));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n516));
  XOR2_X1   g091(.A(KEYINPUT70), .B(G51), .Z(new_n517));
  NAND4_X1  g092(.A1(new_n515), .A2(G543), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n509), .A2(new_n502), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n507), .B1(new_n506), .B2(new_n511), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n512), .A2(new_n518), .A3(new_n521), .A4(new_n522), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  NAND2_X1  g099(.A1(G77), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G64), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n495), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n527), .A2(G651), .B1(new_n520), .B2(G90), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(new_n513), .B2(new_n514), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G52), .A3(new_n516), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  NAND2_X1  g108(.A1(G68), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G56), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n495), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n536), .A2(G651), .B1(new_n520), .B2(G81), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n530), .A2(G43), .A3(new_n516), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT71), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT9), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n515), .A2(G543), .A3(new_n516), .ZN(new_n550));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n549), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n551), .B1(KEYINPUT73), .B2(KEYINPUT9), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n530), .A2(new_n516), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n495), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(new_n520), .B2(G91), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n552), .A2(new_n555), .A3(new_n559), .ZN(G299));
  XOR2_X1   g135(.A(new_n504), .B(KEYINPUT74), .Z(G303));
  NAND2_X1  g136(.A1(new_n520), .A2(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n563));
  INV_X1    g138(.A(G49), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n562), .B(new_n563), .C1(new_n550), .C2(new_n564), .ZN(G288));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  INV_X1    g141(.A(G61), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n495), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n509), .A2(KEYINPUT75), .A3(G61), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n509), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(new_n513), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G305));
  XNOR2_X1  g150(.A(KEYINPUT76), .B(G85), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n520), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G47), .ZN(new_n579));
  OAI221_X1 g154(.A(new_n577), .B1(new_n511), .B2(new_n578), .C1(new_n550), .C2(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  XNOR2_X1  g156(.A(KEYINPUT77), .B(KEYINPUT10), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT78), .ZN(new_n583));
  AND3_X1   g158(.A1(new_n509), .A2(new_n502), .A3(G92), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n495), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n515), .A2(G54), .A3(G543), .A4(new_n516), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT79), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n585), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n581), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n581), .B1(new_n595), .B2(G868), .ZN(G321));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G299), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n598), .B2(G168), .ZN(G297));
  XNOR2_X1  g175(.A(G297), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n473), .A2(G2104), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  AOI22_X1  g188(.A1(G123), .A2(new_n475), .B1(new_n473), .B2(G135), .ZN(new_n614));
  NOR3_X1   g189(.A1(new_n467), .A2(KEYINPUT81), .A3(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT81), .B1(new_n467), .B2(G111), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n616), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n614), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(G156));
  INV_X1    g195(.A(G14), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n630), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n621), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n627), .A2(new_n628), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n627), .A2(new_n628), .ZN(new_n640));
  AND3_X1   g215(.A1(new_n639), .A2(new_n633), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n633), .B1(new_n639), .B2(new_n640), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n638), .B1(new_n643), .B2(new_n635), .ZN(new_n644));
  NOR4_X1   g219(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT83), .A4(new_n636), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n637), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT85), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2084), .B(G2090), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT84), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT17), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n654), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n648), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n657), .B(new_n660), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n654), .A3(new_n648), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n662), .A2(new_n663), .A3(new_n659), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2096), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(new_n611), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n669), .A2(G2096), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(G2096), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(G2100), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  INV_X1    g251(.A(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n682), .A2(KEYINPUT19), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n682), .A2(KEYINPUT19), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n684), .A2(new_n685), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n683), .B2(new_n691), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n683), .A2(new_n691), .A3(new_n696), .ZN(new_n699));
  NAND4_X1  g274(.A1(new_n694), .A2(new_n695), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n699), .A2(new_n693), .A3(new_n688), .ZN(new_n701));
  OAI21_X1  g276(.A(G1986), .B1(new_n701), .B2(new_n697), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AND3_X1   g279(.A1(new_n700), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n704), .B1(new_n700), .B2(new_n702), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n679), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(new_n702), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(new_n703), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n700), .A2(new_n702), .A3(new_n704), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n709), .A2(new_n678), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  INV_X1    g288(.A(G28), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT30), .ZN(new_n715));
  AOI21_X1  g290(.A(G29), .B1(new_n714), .B2(KEYINPUT30), .ZN(new_n716));
  OR2_X1    g291(.A1(KEYINPUT31), .A2(G11), .ZN(new_n717));
  NAND2_X1  g292(.A1(KEYINPUT31), .A2(G11), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n715), .A2(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n473), .A2(G141), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n475), .A2(G129), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT26), .Z(new_n724));
  NAND3_X1  g299(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n721), .A2(new_n722), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(new_n720), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n720), .B2(G32), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  OAI221_X1 g305(.A(new_n719), .B1(new_n720), .B2(new_n618), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n720), .A2(G33), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT97), .B(KEYINPUT25), .ZN(new_n734));
  AND3_X1   g309(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n473), .A2(G139), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT3), .ZN(new_n738));
  INV_X1    g313(.A(G2104), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n742), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n736), .B(new_n737), .C1(new_n467), .C2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n733), .B1(new_n746), .B2(new_n720), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n732), .B1(G2072), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G16), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n540), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n749), .B2(G19), .ZN(new_n751));
  INV_X1    g326(.A(G1341), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G171), .A2(new_n749), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G5), .B2(new_n749), .ZN(new_n755));
  INV_X1    g330(.A(G1961), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n720), .A2(G35), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G162), .B2(new_n720), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT29), .B(G2090), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n749), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n749), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G1966), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n753), .A2(new_n757), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n748), .A2(new_n765), .ZN(new_n766));
  OAI22_X1  g341(.A1(new_n751), .A2(new_n752), .B1(new_n763), .B2(G1966), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n473), .A2(G140), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n475), .A2(G128), .ZN(new_n769));
  OR2_X1    g344(.A1(G104), .A2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n720), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2067), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n755), .B2(new_n756), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT24), .ZN(new_n781));
  INV_X1    g356(.A(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n781), .B2(new_n782), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G160), .B2(new_n720), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2084), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n747), .A2(G2072), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n749), .A2(G4), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n595), .B2(new_n749), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n786), .B(new_n787), .C1(G1348), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n766), .A2(new_n780), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(G299), .A2(G16), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n749), .A2(G20), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT23), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G1956), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G1348), .B2(new_n789), .ZN(new_n798));
  NOR2_X1   g373(.A1(G27), .A2(G29), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G164), .B2(G29), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2078), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n791), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT99), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n749), .A2(G23), .ZN(new_n804));
  INV_X1    g379(.A(G288), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n749), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT93), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT33), .B(G1976), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n807), .B(new_n808), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n749), .A2(G22), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G166), .B2(new_n749), .ZN(new_n811));
  INV_X1    g386(.A(G1971), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n749), .A2(G6), .ZN(new_n817));
  INV_X1    g392(.A(G305), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n749), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT92), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT32), .B(G1981), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OR3_X1    g397(.A1(new_n814), .A2(new_n816), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n816), .B1(new_n814), .B2(new_n822), .ZN(new_n824));
  MUX2_X1   g399(.A(G24), .B(G290), .S(G16), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1986), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n720), .A2(G25), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT89), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n475), .A2(G119), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT90), .ZN(new_n830));
  OR2_X1    g405(.A1(G95), .A2(G2105), .ZN(new_n831));
  INV_X1    g406(.A(G107), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n739), .B1(new_n832), .B2(G2105), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n473), .A2(G131), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n828), .B1(new_n835), .B2(G29), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT35), .B(G1991), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n826), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n823), .A2(new_n824), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(KEYINPUT96), .A2(KEYINPUT36), .ZN(new_n841));
  AND2_X1   g416(.A1(KEYINPUT96), .A2(KEYINPUT36), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(KEYINPUT94), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n823), .A2(new_n845), .A3(new_n824), .A4(new_n839), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(KEYINPUT36), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n844), .A2(KEYINPUT95), .A3(KEYINPUT36), .A4(new_n846), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n803), .B1(new_n849), .B2(new_n850), .ZN(G311));
  INV_X1    g426(.A(G311), .ZN(G150));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  INV_X1    g428(.A(G67), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n495), .B2(new_n854), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n855), .A2(G651), .B1(new_n520), .B2(G93), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n530), .A2(G55), .A3(new_n516), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n539), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n537), .A2(new_n856), .A3(new_n538), .A4(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT38), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n595), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n865), .A2(new_n866), .A3(G860), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n858), .A2(G860), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT37), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n473), .A2(G142), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT102), .ZN(new_n873));
  OR2_X1    g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  INV_X1    g449(.A(G118), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n739), .B1(new_n875), .B2(G2105), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n475), .A2(G130), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n609), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n609), .B1(new_n873), .B2(new_n877), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n879), .A2(new_n880), .A3(new_n835), .ZN(new_n881));
  INV_X1    g456(.A(new_n835), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n873), .A2(new_n877), .ZN(new_n883));
  INV_X1    g458(.A(new_n609), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n882), .B1(new_n885), .B2(new_n878), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n871), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n835), .B1(new_n879), .B2(new_n880), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n882), .A3(new_n878), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT103), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n726), .B(new_n772), .Z(new_n892));
  INV_X1    g467(.A(new_n481), .ZN(new_n893));
  INV_X1    g468(.A(G126), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n740), .B2(new_n741), .ZN(new_n895));
  INV_X1    g470(.A(new_n483), .ZN(new_n896));
  OAI21_X1  g471(.A(G2105), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n893), .B1(new_n897), .B2(KEYINPUT4), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT100), .B1(new_n898), .B2(new_n489), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n486), .A2(new_n900), .A3(new_n490), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n726), .B(new_n772), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n744), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n746), .B1(KEYINPUT98), .B2(KEYINPUT101), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n906), .A3(new_n903), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n891), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n912), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n890), .A3(new_n887), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G160), .B(new_n479), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(new_n618), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n888), .A2(new_n889), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n915), .B(new_n918), .C1(new_n922), .C2(new_n914), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g500(.A1(new_n858), .A2(new_n598), .ZN(new_n926));
  NAND2_X1  g501(.A1(G288), .A2(KEYINPUT105), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(G288), .A2(KEYINPUT105), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n818), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(G290), .B(new_n504), .ZN(new_n931));
  OR2_X1    g506(.A1(G288), .A2(KEYINPUT105), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(G305), .A3(new_n927), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n931), .B1(new_n930), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT42), .Z(new_n937));
  NAND2_X1  g512(.A1(G299), .A2(KEYINPUT104), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n552), .A2(new_n939), .A3(new_n555), .A4(new_n559), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n595), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n583), .A2(new_n584), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n583), .A2(new_n584), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT79), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT79), .B1(new_n589), .B2(new_n590), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n942), .B(new_n943), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(KEYINPUT104), .A3(G299), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT41), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n941), .A2(KEYINPUT41), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n604), .B(new_n861), .Z(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n941), .A2(new_n947), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n937), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n926), .B1(new_n957), .B2(new_n598), .ZN(G295));
  XOR2_X1   g533(.A(G295), .B(KEYINPUT106), .Z(G331));
  NAND2_X1  g534(.A1(G301), .A2(G286), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n510), .A2(new_n511), .ZN(new_n961));
  INV_X1    g536(.A(G89), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n522), .B1(new_n519), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n964), .A2(new_n528), .A3(new_n518), .A4(new_n531), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n861), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n859), .A2(new_n960), .A3(new_n860), .A4(new_n965), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n950), .A2(new_n951), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n968), .A2(new_n971), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n955), .A2(new_n967), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n974), .A3(new_n936), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n970), .A2(new_n974), .A3(new_n936), .A4(KEYINPUT109), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n977), .A2(new_n921), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n936), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n973), .A2(new_n967), .A3(new_n972), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n981), .A2(new_n951), .A3(new_n950), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n948), .A2(new_n969), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n970), .A2(new_n974), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n980), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n977), .A2(new_n988), .A3(new_n921), .A4(new_n978), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n986), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n979), .A2(KEYINPUT110), .A3(new_n991), .A4(new_n984), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n993));
  AOI21_X1  g568(.A(G37), .B1(new_n975), .B2(new_n976), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n994), .A2(new_n984), .A3(new_n991), .A4(new_n978), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n992), .A2(new_n993), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n990), .B1(new_n999), .B2(new_n1000), .ZN(G397));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n904), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n471), .A2(new_n467), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n465), .B1(new_n462), .B2(G2105), .ZN(new_n1008));
  AOI211_X1 g583(.A(KEYINPUT67), .B(new_n467), .C1(new_n460), .C2(new_n461), .ZN(new_n1009));
  OAI211_X1 g584(.A(G40), .B(new_n1007), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1002), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1010), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1004), .A2(KEYINPUT111), .A3(new_n1005), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1996), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(KEYINPUT112), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n1014), .B2(G1996), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n726), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n772), .B(new_n777), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n1016), .B2(new_n727), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1020), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n882), .A2(new_n837), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n882), .A2(new_n837), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1015), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(G290), .B(G1986), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1015), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT123), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G303), .A2(G8), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n1031), .B(KEYINPUT55), .Z(new_n1032));
  NAND4_X1  g607(.A1(new_n899), .A2(KEYINPUT45), .A3(new_n1003), .A4(new_n901), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1033), .A2(new_n1012), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT68), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n898), .B2(new_n489), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n486), .A2(KEYINPUT68), .A3(new_n490), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1035), .B1(new_n1039), .B2(KEYINPUT45), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1003), .B1(new_n491), .B2(new_n492), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(KEYINPUT113), .A3(new_n1005), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1034), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n812), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1384), .B1(new_n486), .B2(new_n490), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1010), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1039), .B2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n1044), .A2(new_n1045), .B1(G2090), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT114), .B1(new_n1043), .B2(new_n812), .ZN(new_n1052));
  OAI211_X1 g627(.A(G8), .B(new_n1032), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G305), .A2(G1981), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n572), .A2(new_n677), .A3(new_n574), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT49), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(KEYINPUT49), .A3(new_n1055), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n1012), .B2(new_n1046), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1012), .A2(new_n1046), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n805), .A2(G1976), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(G8), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT116), .B1(new_n1067), .B2(KEYINPUT52), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n805), .B2(G1976), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1067), .A2(KEYINPUT116), .A3(new_n1070), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1064), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G288), .A2(G1976), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1064), .A2(new_n1076), .B1(new_n677), .B2(new_n818), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1061), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1053), .A2(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1073), .B(new_n1072), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1032), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1003), .B1(new_n898), .B2(new_n489), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1047), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1010), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1041), .B2(KEYINPUT50), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(G2090), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n812), .B2(new_n1043), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1083), .B1(new_n1089), .B2(new_n1060), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1010), .B1(new_n1084), .B2(new_n1005), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n1041), .B2(new_n1005), .ZN(new_n1092));
  INV_X1    g667(.A(G1966), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1041), .A2(KEYINPUT50), .ZN(new_n1095));
  INV_X1    g670(.A(G2084), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1048), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G8), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(G286), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1053), .A2(new_n1082), .A3(new_n1090), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(G8), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1083), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1075), .A2(new_n1102), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1053), .A4(new_n1100), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1079), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(G299), .B(KEYINPUT57), .Z(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1034), .A2(new_n1040), .A3(new_n1042), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1087), .A2(new_n796), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1348), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1095), .B2(new_n1048), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1115), .B(new_n1048), .C1(new_n1039), .C2(new_n1049), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1114), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1065), .A2(G2067), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n946), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1111), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1113), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1050), .A2(KEYINPUT118), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1348), .B1(new_n1126), .B2(new_n1117), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n1120), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT120), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n1121), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n946), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n946), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1128), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1109), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1123), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1034), .A2(new_n1040), .A3(new_n1042), .A4(new_n1016), .ZN(new_n1144));
  XOR2_X1   g719(.A(KEYINPUT58), .B(G1341), .Z(new_n1145));
  NAND2_X1  g720(.A1(new_n1065), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1143), .B1(new_n1147), .B2(new_n540), .ZN(new_n1148));
  AOI211_X1 g723(.A(KEYINPUT59), .B(new_n539), .C1(new_n1144), .C2(new_n1146), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1142), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1111), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(new_n1113), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT119), .B(new_n1151), .C1(new_n1152), .C2(new_n1113), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1150), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1125), .B1(new_n1138), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(G286), .A2(G8), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT121), .Z(new_n1160));
  NAND3_X1  g735(.A1(new_n1099), .A2(KEYINPUT51), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1160), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1098), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT51), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1060), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(new_n1162), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1161), .A2(new_n1163), .A3(new_n1166), .ZN(new_n1167));
  AND4_X1   g742(.A1(new_n1053), .A2(new_n1167), .A3(new_n1082), .A4(new_n1090), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT53), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n1043), .B2(G2078), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n756), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1169), .A2(G2078), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1172), .B(new_n1091), .C1(new_n1041), .C2(new_n1005), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(G171), .ZN(new_n1175));
  AND4_X1   g750(.A1(G40), .A2(new_n1007), .A3(new_n463), .A4(new_n1172), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1006), .A2(new_n1033), .A3(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1170), .A2(new_n1171), .A3(G301), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT54), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1170), .A2(new_n1171), .A3(new_n1177), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(G301), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT54), .B1(new_n1174), .B2(G171), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1168), .B(new_n1180), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1030), .B(new_n1108), .C1(new_n1158), .C2(new_n1187), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1053), .A2(new_n1090), .A3(new_n1082), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n1167), .A2(KEYINPUT62), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1175), .B1(new_n1167), .B2(KEYINPUT62), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT124), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1188), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n595), .B1(new_n1129), .B2(KEYINPUT120), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1131), .A2(new_n1132), .A3(new_n946), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1197), .A2(new_n1130), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1152), .A2(new_n1113), .A3(new_n1151), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1124), .B1(new_n1198), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1186), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1053), .A2(new_n1167), .A3(new_n1082), .A4(new_n1090), .ZN(new_n1206));
  NOR3_X1   g781(.A1(new_n1205), .A2(new_n1206), .A3(new_n1179), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1030), .B1(new_n1208), .B2(new_n1108), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1029), .B1(new_n1194), .B2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n772), .A2(G2067), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1211), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1014), .A2(G1986), .A3(G290), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1213), .B(KEYINPUT48), .ZN(new_n1214));
  OAI22_X1  g789(.A1(new_n1212), .A2(new_n1014), .B1(new_n1027), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1021), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1015), .B1(new_n726), .B2(new_n1216), .ZN(new_n1217));
  AND3_X1   g792(.A1(new_n1017), .A2(KEYINPUT46), .A3(new_n1019), .ZN(new_n1218));
  AOI21_X1  g793(.A(KEYINPUT46), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT47), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n1223));
  OAI211_X1 g798(.A(KEYINPUT47), .B(new_n1217), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1224));
  AND3_X1   g799(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1223), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1226));
  NOR3_X1   g801(.A1(new_n1215), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1210), .A2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g803(.A1(new_n671), .A2(G319), .A3(new_n674), .ZN(new_n1230));
  AND3_X1   g804(.A1(new_n712), .A2(new_n1230), .A3(new_n646), .ZN(new_n1231));
  NAND2_X1  g805(.A1(new_n924), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g806(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n998), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g810(.A(KEYINPUT127), .ZN(new_n1237));
  NAND3_X1  g811(.A1(new_n998), .A2(KEYINPUT126), .A3(new_n1233), .ZN(new_n1238));
  NAND3_X1  g812(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g813(.A(KEYINPUT126), .B1(new_n998), .B2(new_n1233), .ZN(new_n1240));
  AOI22_X1  g814(.A1(new_n995), .A2(new_n996), .B1(new_n989), .B2(KEYINPUT43), .ZN(new_n1241));
  AOI211_X1 g815(.A(new_n1235), .B(new_n1232), .C1(new_n1241), .C2(new_n992), .ZN(new_n1242));
  OAI21_X1  g816(.A(KEYINPUT127), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  AND2_X1   g817(.A1(new_n1239), .A2(new_n1243), .ZN(G308));
  NAND2_X1  g818(.A1(new_n1236), .A2(new_n1238), .ZN(G225));
endmodule


