

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752;

  AND2_X1 U371 ( .A1(n568), .A2(n377), .ZN(n376) );
  XNOR2_X1 U372 ( .A(n543), .B(KEYINPUT32), .ZN(n621) );
  BUF_X1 U373 ( .A(n537), .Z(n647) );
  NAND2_X1 U374 ( .A1(n579), .A2(n500), .ZN(n502) );
  INV_X1 U375 ( .A(n532), .ZN(n649) );
  XNOR2_X1 U376 ( .A(n418), .B(n417), .ZN(n701) );
  XNOR2_X1 U377 ( .A(G146), .B(n736), .ZN(n415) );
  XNOR2_X1 U378 ( .A(n383), .B(KEYINPUT64), .ZN(n384) );
  NOR2_X1 U379 ( .A1(G953), .A2(G237), .ZN(n455) );
  INV_X2 U380 ( .A(G953), .ZN(n742) );
  OR2_X2 U381 ( .A1(n686), .A2(n603), .ZN(n689) );
  NOR2_X2 U382 ( .A1(n618), .A2(n720), .ZN(n620) );
  NOR2_X2 U383 ( .A1(n699), .A2(n720), .ZN(n700) );
  NOR2_X2 U384 ( .A1(n710), .A2(n720), .ZN(n711) );
  NOR2_X2 U385 ( .A1(n544), .A2(n400), .ZN(n401) );
  XNOR2_X2 U386 ( .A(n505), .B(n399), .ZN(n544) );
  OR2_X2 U387 ( .A1(n360), .A2(n358), .ZN(n511) );
  NAND2_X1 U388 ( .A1(n649), .A2(n484), .ZN(n513) );
  XNOR2_X1 U389 ( .A(G128), .B(G137), .ZN(n421) );
  BUF_X1 U390 ( .A(n716), .Z(n350) );
  AND2_X2 U391 ( .A1(n689), .A2(n604), .ZN(n349) );
  XNOR2_X2 U392 ( .A(n398), .B(n397), .ZN(n505) );
  AND2_X2 U393 ( .A1(n622), .A2(n751), .ZN(n551) );
  AND2_X4 U394 ( .A1(n349), .A2(n612), .ZN(n716) );
  XNOR2_X2 U395 ( .A(n563), .B(KEYINPUT31), .ZN(n639) );
  XNOR2_X2 U396 ( .A(n447), .B(n446), .ZN(n696) );
  XNOR2_X2 U397 ( .A(n410), .B(n409), .ZN(n447) );
  NOR2_X1 U398 ( .A1(n607), .A2(n606), .ZN(n682) );
  OR2_X1 U399 ( .A1(n558), .A2(n557), .ZN(n351) );
  XNOR2_X1 U400 ( .A(n492), .B(n491), .ZN(n676) );
  NOR2_X1 U401 ( .A1(n663), .A2(n370), .ZN(n369) );
  OR2_X2 U402 ( .A1(n581), .A2(n676), .ZN(n493) );
  NAND2_X1 U403 ( .A1(n371), .A2(n525), .ZN(n527) );
  NAND2_X1 U404 ( .A1(n362), .A2(n361), .ZN(n360) );
  NAND2_X1 U405 ( .A1(n420), .A2(n396), .ZN(n359) );
  XNOR2_X1 U406 ( .A(n432), .B(n431), .ZN(n532) );
  XNOR2_X1 U407 ( .A(n430), .B(n379), .ZN(n431) );
  INV_X1 U408 ( .A(KEYINPUT96), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n489), .B(KEYINPUT110), .ZN(n370) );
  XNOR2_X1 U410 ( .A(G137), .B(G134), .ZN(n386) );
  INV_X1 U411 ( .A(G140), .ZN(n411) );
  XNOR2_X1 U412 ( .A(G119), .B(KEYINPUT3), .ZN(n391) );
  XNOR2_X1 U413 ( .A(G113), .B(KEYINPUT85), .ZN(n390) );
  XNOR2_X1 U414 ( .A(n357), .B(KEYINPUT23), .ZN(n423) );
  INV_X1 U415 ( .A(KEYINPUT91), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n440), .B(n439), .ZN(n723) );
  XNOR2_X1 U417 ( .A(n472), .B(KEYINPUT16), .ZN(n439) );
  XNOR2_X1 U418 ( .A(n372), .B(n523), .ZN(n371) );
  AND2_X1 U419 ( .A1(n537), .A2(n649), .ZN(n538) );
  BUF_X1 U420 ( .A(n505), .Z(n645) );
  INV_X1 U421 ( .A(G469), .ZN(n419) );
  NAND2_X1 U422 ( .A1(n363), .A2(G902), .ZN(n361) );
  XOR2_X1 U423 ( .A(G116), .B(G122), .Z(n472) );
  AND2_X1 U424 ( .A1(n622), .A2(n556), .ZN(n557) );
  BUF_X1 U425 ( .A(n682), .Z(n741) );
  XOR2_X1 U426 ( .A(G104), .B(G113), .Z(n463) );
  XNOR2_X1 U427 ( .A(n521), .B(KEYINPUT33), .ZN(n678) );
  INV_X1 U428 ( .A(n666), .ZN(n367) );
  INV_X1 U429 ( .A(KEYINPUT89), .ZN(n503) );
  XNOR2_X1 U430 ( .A(n364), .B(n738), .ZN(n717) );
  NAND2_X1 U431 ( .A1(n611), .A2(n683), .ZN(n612) );
  AND2_X1 U432 ( .A1(n617), .A2(G953), .ZN(n720) );
  XOR2_X1 U433 ( .A(n421), .B(G119), .Z(n352) );
  XNOR2_X1 U434 ( .A(n374), .B(n569), .ZN(n686) );
  INV_X1 U435 ( .A(n420), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n419), .B(KEYINPUT70), .ZN(n420) );
  AND2_X1 U437 ( .A1(n621), .A2(n559), .ZN(n353) );
  XNOR2_X2 U438 ( .A(n387), .B(G131), .ZN(n736) );
  XNOR2_X1 U439 ( .A(n438), .B(KEYINPUT76), .ZN(n570) );
  NAND2_X1 U440 ( .A1(n351), .A2(n353), .ZN(n375) );
  NOR2_X2 U441 ( .A1(n544), .A2(n513), .ZN(n485) );
  NAND2_X1 U442 ( .A1(n376), .A2(n375), .ZN(n374) );
  NOR2_X2 U443 ( .A1(n623), .A2(n639), .ZN(n356) );
  XNOR2_X1 U444 ( .A(n356), .B(n355), .ZN(n354) );
  NAND2_X1 U445 ( .A1(n354), .A2(n566), .ZN(n567) );
  XNOR2_X2 U446 ( .A(n507), .B(KEYINPUT95), .ZN(n623) );
  XNOR2_X2 U447 ( .A(n511), .B(KEYINPUT1), .ZN(n537) );
  NOR2_X1 U448 ( .A1(n701), .A2(n359), .ZN(n358) );
  NAND2_X1 U449 ( .A1(n701), .A2(n363), .ZN(n362) );
  NOR2_X1 U450 ( .A1(n717), .A2(G902), .ZN(n432) );
  XNOR2_X1 U451 ( .A(n366), .B(n365), .ZN(n364) );
  XNOR2_X1 U452 ( .A(n424), .B(n352), .ZN(n365) );
  NAND2_X1 U453 ( .A1(n478), .A2(G221), .ZN(n366) );
  NAND2_X1 U454 ( .A1(n368), .A2(n367), .ZN(n492) );
  INV_X1 U455 ( .A(n370), .ZN(n368) );
  NAND2_X1 U456 ( .A1(n522), .A2(n678), .ZN(n372) );
  XNOR2_X1 U457 ( .A(n562), .B(n503), .ZN(n522) );
  XNOR2_X2 U458 ( .A(n373), .B(G143), .ZN(n473) );
  XNOR2_X2 U459 ( .A(G128), .B(KEYINPUT65), .ZN(n373) );
  NAND2_X1 U460 ( .A1(n554), .A2(n553), .ZN(n377) );
  AND2_X1 U461 ( .A1(n506), .A2(n645), .ZN(n378) );
  XOR2_X1 U462 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n379) );
  INV_X1 U463 ( .A(KEYINPUT77), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U465 ( .A(n393), .B(n440), .ZN(n394) );
  XNOR2_X1 U466 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U467 ( .A(n415), .B(n394), .ZN(n395) );
  NOR2_X2 U468 ( .A1(n437), .A2(n504), .ZN(n438) );
  XNOR2_X1 U469 ( .A(n712), .B(KEYINPUT120), .ZN(n713) );
  BUF_X1 U470 ( .A(n628), .Z(n633) );
  XNOR2_X1 U471 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U472 ( .A1(G237), .A2(G902), .ZN(n380) );
  XOR2_X1 U473 ( .A(KEYINPUT74), .B(n380), .Z(n449) );
  NAND2_X1 U474 ( .A1(n449), .A2(G214), .ZN(n382) );
  INV_X1 U475 ( .A(KEYINPUT87), .ZN(n381) );
  XNOR2_X1 U476 ( .A(n382), .B(n381), .ZN(n664) );
  INV_X1 U477 ( .A(n664), .ZN(n400) );
  XNOR2_X2 U478 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n383) );
  XNOR2_X2 U479 ( .A(n473), .B(n384), .ZN(n737) );
  XNOR2_X1 U480 ( .A(KEYINPUT67), .B(G101), .ZN(n385) );
  XNOR2_X2 U481 ( .A(n737), .B(n385), .ZN(n410) );
  INV_X1 U482 ( .A(n386), .ZN(n387) );
  XOR2_X1 U483 ( .A(KEYINPUT5), .B(G116), .Z(n389) );
  NAND2_X1 U484 ( .A1(n455), .A2(G210), .ZN(n388) );
  XNOR2_X1 U485 ( .A(n389), .B(n388), .ZN(n393) );
  INV_X1 U486 ( .A(n390), .ZN(n392) );
  XNOR2_X1 U487 ( .A(n392), .B(n391), .ZN(n440) );
  XNOR2_X1 U488 ( .A(n410), .B(n395), .ZN(n614) );
  INV_X1 U489 ( .A(G902), .ZN(n396) );
  NAND2_X1 U490 ( .A1(n614), .A2(n396), .ZN(n398) );
  INV_X1 U491 ( .A(G472), .ZN(n397) );
  INV_X1 U492 ( .A(KEYINPUT107), .ZN(n399) );
  XNOR2_X1 U493 ( .A(n401), .B(KEYINPUT30), .ZN(n407) );
  NAND2_X1 U494 ( .A1(G234), .A2(G237), .ZN(n402) );
  XNOR2_X1 U495 ( .A(n402), .B(KEYINPUT14), .ZN(n403) );
  NAND2_X1 U496 ( .A1(G952), .A2(n403), .ZN(n675) );
  NOR2_X1 U497 ( .A1(G953), .A2(n675), .ZN(n498) );
  AND2_X1 U498 ( .A1(G953), .A2(n403), .ZN(n404) );
  NAND2_X1 U499 ( .A1(G902), .A2(n404), .ZN(n496) );
  NOR2_X1 U500 ( .A1(G900), .A2(n496), .ZN(n405) );
  NOR2_X1 U501 ( .A1(n498), .A2(n405), .ZN(n483) );
  INV_X1 U502 ( .A(n483), .ZN(n406) );
  NAND2_X1 U503 ( .A1(n407), .A2(n406), .ZN(n437) );
  XNOR2_X1 U504 ( .A(G110), .B(G107), .ZN(n408) );
  XNOR2_X1 U505 ( .A(n408), .B(G104), .ZN(n721) );
  XNOR2_X1 U506 ( .A(n721), .B(KEYINPUT71), .ZN(n409) );
  XNOR2_X1 U507 ( .A(n447), .B(n411), .ZN(n418) );
  NAND2_X1 U508 ( .A1(G227), .A2(n742), .ZN(n413) );
  XOR2_X1 U509 ( .A(n416), .B(KEYINPUT90), .Z(n417) );
  XNOR2_X1 U510 ( .A(G110), .B(KEYINPUT24), .ZN(n422) );
  XNOR2_X1 U511 ( .A(n423), .B(n422), .ZN(n424) );
  NAND2_X1 U512 ( .A1(G234), .A2(n742), .ZN(n425) );
  XOR2_X1 U513 ( .A(KEYINPUT8), .B(n425), .Z(n478) );
  INV_X1 U514 ( .A(G146), .ZN(n426) );
  XNOR2_X1 U515 ( .A(n426), .B(G125), .ZN(n444) );
  XNOR2_X1 U516 ( .A(G140), .B(n444), .ZN(n427) );
  XNOR2_X1 U517 ( .A(n427), .B(KEYINPUT10), .ZN(n738) );
  XNOR2_X1 U518 ( .A(G902), .B(KEYINPUT15), .ZN(n448) );
  NAND2_X1 U519 ( .A1(n448), .A2(G234), .ZN(n429) );
  XNOR2_X1 U520 ( .A(KEYINPUT92), .B(KEYINPUT20), .ZN(n428) );
  XNOR2_X1 U521 ( .A(n429), .B(n428), .ZN(n433) );
  NAND2_X1 U522 ( .A1(n433), .A2(G217), .ZN(n430) );
  NAND2_X1 U523 ( .A1(n433), .A2(G221), .ZN(n434) );
  XNOR2_X1 U524 ( .A(n434), .B(KEYINPUT94), .ZN(n435) );
  XNOR2_X1 U525 ( .A(n435), .B(KEYINPUT21), .ZN(n650) );
  INV_X1 U526 ( .A(n650), .ZN(n436) );
  NAND2_X1 U527 ( .A1(n532), .A2(n436), .ZN(n560) );
  INV_X1 U528 ( .A(n560), .ZN(n646) );
  NAND2_X1 U529 ( .A1(n511), .A2(n646), .ZN(n504) );
  XNOR2_X1 U530 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n442) );
  NAND2_X1 U531 ( .A1(n742), .A2(G224), .ZN(n441) );
  XNOR2_X1 U532 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U533 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U534 ( .A(n723), .B(n445), .ZN(n446) );
  INV_X1 U535 ( .A(n448), .ZN(n604) );
  OR2_X2 U536 ( .A1(n696), .A2(n604), .ZN(n453) );
  NAND2_X1 U537 ( .A1(n449), .A2(G210), .ZN(n451) );
  INV_X1 U538 ( .A(KEYINPUT86), .ZN(n450) );
  XNOR2_X1 U539 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X2 U540 ( .A(n453), .B(n452), .ZN(n494) );
  BUF_X1 U541 ( .A(n494), .Z(n454) );
  INV_X1 U542 ( .A(n454), .ZN(n518) );
  XNOR2_X1 U543 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n468) );
  XOR2_X1 U544 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n457) );
  NAND2_X1 U545 ( .A1(G214), .A2(n455), .ZN(n456) );
  XNOR2_X1 U546 ( .A(n457), .B(n456), .ZN(n461) );
  XOR2_X1 U547 ( .A(KEYINPUT97), .B(KEYINPUT99), .Z(n459) );
  XNOR2_X1 U548 ( .A(G122), .B(KEYINPUT98), .ZN(n458) );
  XNOR2_X1 U549 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U550 ( .A(n461), .B(n460), .Z(n466) );
  XNOR2_X1 U551 ( .A(G143), .B(G131), .ZN(n462) );
  XNOR2_X1 U552 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U553 ( .A(n738), .B(n464), .ZN(n465) );
  XNOR2_X1 U554 ( .A(n466), .B(n465), .ZN(n707) );
  NOR2_X1 U555 ( .A1(G902), .A2(n707), .ZN(n467) );
  XNOR2_X1 U556 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U557 ( .A(n469), .B(G475), .ZN(n565) );
  INV_X1 U558 ( .A(n565), .ZN(n490) );
  XOR2_X1 U559 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n471) );
  XNOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT9), .ZN(n470) );
  XNOR2_X1 U561 ( .A(n471), .B(n470), .ZN(n477) );
  XOR2_X1 U562 ( .A(n472), .B(G107), .Z(n475) );
  XNOR2_X1 U563 ( .A(n473), .B(G134), .ZN(n474) );
  XNOR2_X1 U564 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U565 ( .A(n477), .B(n476), .Z(n480) );
  NAND2_X1 U566 ( .A1(G217), .A2(n478), .ZN(n479) );
  XNOR2_X1 U567 ( .A(n480), .B(n479), .ZN(n712) );
  NOR2_X1 U568 ( .A1(n712), .A2(G902), .ZN(n481) );
  XNOR2_X1 U569 ( .A(n481), .B(G478), .ZN(n564) );
  OR2_X1 U570 ( .A1(n490), .A2(n564), .ZN(n524) );
  NOR2_X1 U571 ( .A1(n518), .A2(n524), .ZN(n482) );
  NAND2_X1 U572 ( .A1(n570), .A2(n482), .ZN(n585) );
  XNOR2_X1 U573 ( .A(n585), .B(G143), .ZN(G45) );
  NOR2_X1 U574 ( .A1(n483), .A2(n650), .ZN(n484) );
  XNOR2_X1 U575 ( .A(n485), .B(KEYINPUT28), .ZN(n486) );
  NAND2_X1 U576 ( .A1(n486), .A2(n511), .ZN(n487) );
  XNOR2_X1 U577 ( .A(n487), .B(KEYINPUT108), .ZN(n581) );
  INV_X1 U578 ( .A(KEYINPUT38), .ZN(n488) );
  XNOR2_X1 U579 ( .A(n494), .B(n488), .ZN(n665) );
  NAND2_X1 U580 ( .A1(n665), .A2(n664), .ZN(n489) );
  NAND2_X1 U581 ( .A1(n490), .A2(n564), .ZN(n666) );
  INV_X1 U582 ( .A(KEYINPUT41), .ZN(n491) );
  XNOR2_X2 U583 ( .A(n493), .B(KEYINPUT42), .ZN(n575) );
  XNOR2_X1 U584 ( .A(n575), .B(G137), .ZN(G39) );
  NAND2_X1 U585 ( .A1(n494), .A2(n664), .ZN(n495) );
  XNOR2_X2 U586 ( .A(n495), .B(KEYINPUT19), .ZN(n579) );
  NOR2_X1 U587 ( .A1(G898), .A2(n496), .ZN(n497) );
  OR2_X1 U588 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U589 ( .A(n499), .B(KEYINPUT88), .ZN(n500) );
  INV_X1 U590 ( .A(KEYINPUT0), .ZN(n501) );
  XNOR2_X2 U591 ( .A(n502), .B(n501), .ZN(n562) );
  INV_X1 U592 ( .A(n504), .ZN(n506) );
  NAND2_X1 U593 ( .A1(n522), .A2(n378), .ZN(n507) );
  NAND2_X1 U594 ( .A1(n564), .A2(n565), .ZN(n509) );
  INV_X1 U595 ( .A(KEYINPUT103), .ZN(n508) );
  XNOR2_X1 U596 ( .A(n509), .B(n508), .ZN(n634) );
  INV_X1 U597 ( .A(n634), .ZN(n636) );
  NAND2_X1 U598 ( .A1(n623), .A2(n636), .ZN(n510) );
  XNOR2_X1 U599 ( .A(n510), .B(G104), .ZN(G6) );
  INV_X1 U600 ( .A(KEYINPUT6), .ZN(n512) );
  XNOR2_X1 U601 ( .A(n645), .B(n512), .ZN(n539) );
  NOR2_X1 U602 ( .A1(n634), .A2(n513), .ZN(n514) );
  NAND2_X1 U603 ( .A1(n514), .A2(n664), .ZN(n515) );
  NOR2_X1 U604 ( .A1(n539), .A2(n515), .ZN(n589) );
  INV_X1 U605 ( .A(n589), .ZN(n516) );
  OR2_X1 U606 ( .A1(n647), .A2(n516), .ZN(n517) );
  XNOR2_X1 U607 ( .A(n517), .B(KEYINPUT43), .ZN(n519) );
  NAND2_X1 U608 ( .A1(n519), .A2(n518), .ZN(n605) );
  XNOR2_X1 U609 ( .A(n605), .B(G140), .ZN(G42) );
  NOR2_X1 U610 ( .A1(n539), .A2(n560), .ZN(n520) );
  NAND2_X1 U611 ( .A1(n537), .A2(n520), .ZN(n521) );
  XOR2_X1 U612 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n523) );
  INV_X1 U613 ( .A(n524), .ZN(n525) );
  INV_X1 U614 ( .A(KEYINPUT35), .ZN(n526) );
  XNOR2_X2 U615 ( .A(n527), .B(n526), .ZN(n622) );
  NOR2_X1 U616 ( .A1(n666), .A2(n650), .ZN(n528) );
  NAND2_X1 U617 ( .A1(n562), .A2(n528), .ZN(n531) );
  INV_X1 U618 ( .A(KEYINPUT66), .ZN(n529) );
  XNOR2_X1 U619 ( .A(n529), .B(KEYINPUT22), .ZN(n530) );
  XNOR2_X1 U620 ( .A(n531), .B(n530), .ZN(n547) );
  NAND2_X1 U621 ( .A1(n539), .A2(n532), .ZN(n533) );
  NOR2_X1 U622 ( .A1(n647), .A2(n533), .ZN(n534) );
  NAND2_X1 U623 ( .A1(n547), .A2(n534), .ZN(n536) );
  INV_X1 U624 ( .A(KEYINPUT105), .ZN(n535) );
  XNOR2_X1 U625 ( .A(n536), .B(n535), .ZN(n751) );
  XNOR2_X1 U626 ( .A(n538), .B(KEYINPUT106), .ZN(n540) );
  AND2_X1 U627 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U628 ( .A(n541), .B(KEYINPUT78), .ZN(n542) );
  NAND2_X1 U629 ( .A1(n542), .A2(n547), .ZN(n543) );
  NAND2_X1 U630 ( .A1(n544), .A2(n649), .ZN(n545) );
  NOR2_X1 U631 ( .A1(n647), .A2(n545), .ZN(n546) );
  AND2_X1 U632 ( .A1(n547), .A2(n546), .ZN(n627) );
  INV_X1 U633 ( .A(KEYINPUT68), .ZN(n548) );
  NOR2_X1 U634 ( .A1(n627), .A2(n548), .ZN(n549) );
  AND2_X1 U635 ( .A1(n621), .A2(n549), .ZN(n550) );
  NAND2_X1 U636 ( .A1(n551), .A2(n550), .ZN(n554) );
  INV_X1 U637 ( .A(n751), .ZN(n552) );
  OR2_X1 U638 ( .A1(n552), .A2(KEYINPUT44), .ZN(n553) );
  NOR2_X1 U639 ( .A1(n622), .A2(KEYINPUT68), .ZN(n558) );
  INV_X1 U640 ( .A(KEYINPUT44), .ZN(n555) );
  AND2_X1 U641 ( .A1(n555), .A2(KEYINPUT68), .ZN(n556) );
  INV_X1 U642 ( .A(n627), .ZN(n559) );
  NOR2_X1 U643 ( .A1(n560), .A2(n645), .ZN(n561) );
  AND2_X1 U644 ( .A1(n647), .A2(n561), .ZN(n659) );
  NAND2_X1 U645 ( .A1(n659), .A2(n562), .ZN(n563) );
  OR2_X1 U646 ( .A1(n565), .A2(n564), .ZN(n629) );
  AND2_X1 U647 ( .A1(n634), .A2(n629), .ZN(n663) );
  INV_X1 U648 ( .A(n663), .ZN(n566) );
  XNOR2_X1 U649 ( .A(n567), .B(KEYINPUT104), .ZN(n568) );
  INV_X1 U650 ( .A(KEYINPUT45), .ZN(n569) );
  NAND2_X1 U651 ( .A1(n570), .A2(n665), .ZN(n571) );
  XNOR2_X2 U652 ( .A(n571), .B(KEYINPUT39), .ZN(n598) );
  NAND2_X1 U653 ( .A1(n598), .A2(n636), .ZN(n574) );
  INV_X1 U654 ( .A(KEYINPUT109), .ZN(n572) );
  XNOR2_X1 U655 ( .A(n572), .B(KEYINPUT40), .ZN(n573) );
  XNOR2_X1 U656 ( .A(n574), .B(n573), .ZN(n752) );
  NAND2_X1 U657 ( .A1(n752), .A2(n575), .ZN(n578) );
  INV_X1 U658 ( .A(KEYINPUT83), .ZN(n576) );
  XOR2_X1 U659 ( .A(n576), .B(KEYINPUT46), .Z(n577) );
  XNOR2_X1 U660 ( .A(n578), .B(n577), .ZN(n596) );
  INV_X1 U661 ( .A(n579), .ZN(n580) );
  NOR2_X1 U662 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U663 ( .A(n582), .B(KEYINPUT79), .ZN(n628) );
  NOR2_X1 U664 ( .A1(n663), .A2(n628), .ZN(n583) );
  XNOR2_X1 U665 ( .A(n583), .B(KEYINPUT47), .ZN(n587) );
  INV_X1 U666 ( .A(KEYINPUT81), .ZN(n584) );
  XNOR2_X1 U667 ( .A(n585), .B(n584), .ZN(n586) );
  NAND2_X1 U668 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U669 ( .A(n588), .B(KEYINPUT73), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n589), .A2(n454), .ZN(n591) );
  XNOR2_X1 U671 ( .A(KEYINPUT111), .B(KEYINPUT36), .ZN(n590) );
  XNOR2_X1 U672 ( .A(n591), .B(n590), .ZN(n592) );
  AND2_X1 U673 ( .A1(n592), .A2(n647), .ZN(n642) );
  INV_X1 U674 ( .A(n642), .ZN(n593) );
  AND2_X1 U675 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U677 ( .A(n597), .B(KEYINPUT48), .ZN(n607) );
  INV_X1 U678 ( .A(n629), .ZN(n638) );
  NAND2_X1 U679 ( .A1(n598), .A2(n638), .ZN(n644) );
  NAND2_X1 U680 ( .A1(n644), .A2(KEYINPUT2), .ZN(n599) );
  XNOR2_X1 U681 ( .A(n599), .B(KEYINPUT80), .ZN(n601) );
  INV_X1 U682 ( .A(n605), .ZN(n600) );
  OR2_X1 U683 ( .A1(n601), .A2(n600), .ZN(n602) );
  OR2_X1 U684 ( .A1(n607), .A2(n602), .ZN(n603) );
  NAND2_X1 U685 ( .A1(n644), .A2(n605), .ZN(n606) );
  XNOR2_X1 U686 ( .A(n682), .B(KEYINPUT75), .ZN(n608) );
  INV_X1 U687 ( .A(n608), .ZN(n610) );
  INV_X1 U688 ( .A(n686), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n716), .A2(G472), .ZN(n616) );
  XOR2_X1 U691 ( .A(KEYINPUT84), .B(KEYINPUT62), .Z(n613) );
  XNOR2_X1 U692 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U693 ( .A(n616), .B(n615), .ZN(n618) );
  INV_X1 U694 ( .A(G952), .ZN(n617) );
  XOR2_X1 U695 ( .A(KEYINPUT112), .B(KEYINPUT63), .Z(n619) );
  XNOR2_X1 U696 ( .A(n620), .B(n619), .ZN(G57) );
  XNOR2_X1 U697 ( .A(n621), .B(G119), .ZN(G21) );
  XNOR2_X1 U698 ( .A(n622), .B(G122), .ZN(G24) );
  NAND2_X1 U699 ( .A1(n623), .A2(n638), .ZN(n625) );
  XOR2_X1 U700 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n624) );
  XNOR2_X1 U701 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U702 ( .A(G107), .B(n626), .ZN(G9) );
  XOR2_X1 U703 ( .A(G110), .B(n627), .Z(G12) );
  NOR2_X1 U704 ( .A1(n629), .A2(n633), .ZN(n631) );
  XNOR2_X1 U705 ( .A(KEYINPUT29), .B(KEYINPUT113), .ZN(n630) );
  XNOR2_X1 U706 ( .A(n631), .B(n630), .ZN(n632) );
  XOR2_X1 U707 ( .A(G128), .B(n632), .Z(G30) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U709 ( .A(G146), .B(n635), .Z(G48) );
  NAND2_X1 U710 ( .A1(n639), .A2(n636), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n637), .B(G113), .ZN(G15) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n640), .B(KEYINPUT114), .ZN(n641) );
  XNOR2_X1 U714 ( .A(G116), .B(n641), .ZN(G18) );
  XNOR2_X1 U715 ( .A(G125), .B(n642), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U717 ( .A(G134), .B(n644), .ZN(G36) );
  INV_X1 U718 ( .A(n645), .ZN(n656) );
  NOR2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U720 ( .A(KEYINPUT50), .B(n648), .Z(n654) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n651), .B(KEYINPUT115), .ZN(n652) );
  XNOR2_X1 U723 ( .A(KEYINPUT49), .B(n652), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U725 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U726 ( .A(n657), .B(KEYINPUT116), .ZN(n658) );
  NOR2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(KEYINPUT117), .ZN(n661) );
  XNOR2_X1 U729 ( .A(KEYINPUT51), .B(n661), .ZN(n662) );
  NOR2_X1 U730 ( .A1(n662), .A2(n676), .ZN(n672) );
  INV_X1 U731 ( .A(n678), .ZN(n670) );
  NOR2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n667) );
  NOR2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U734 ( .A1(n369), .A2(n668), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U737 ( .A(n673), .B(KEYINPUT52), .ZN(n674) );
  NOR2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n680) );
  INV_X1 U739 ( .A(n676), .ZN(n677) );
  AND2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U742 ( .A1(n681), .A2(n742), .ZN(n692) );
  INV_X1 U743 ( .A(n741), .ZN(n684) );
  INV_X1 U744 ( .A(KEYINPUT2), .ZN(n683) );
  NAND2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U746 ( .A(KEYINPUT82), .B(n685), .Z(n688) );
  NOR2_X1 U747 ( .A1(n609), .A2(KEYINPUT2), .ZN(n687) );
  NOR2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n690) );
  AND2_X1 U749 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U750 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U751 ( .A(KEYINPUT53), .B(n693), .ZN(G75) );
  NAND2_X1 U752 ( .A1(n716), .A2(G210), .ZN(n698) );
  XOR2_X1 U753 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n694) );
  XNOR2_X1 U754 ( .A(n694), .B(KEYINPUT55), .ZN(n695) );
  XNOR2_X1 U755 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U756 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U757 ( .A(n700), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U758 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n703) );
  XNOR2_X1 U759 ( .A(n701), .B(KEYINPUT119), .ZN(n702) );
  XNOR2_X1 U760 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U761 ( .A1(n716), .A2(G469), .ZN(n704) );
  XOR2_X1 U762 ( .A(n705), .B(n704), .Z(n706) );
  NOR2_X1 U763 ( .A1(n720), .A2(n706), .ZN(G54) );
  NAND2_X1 U764 ( .A1(n716), .A2(G475), .ZN(n709) );
  XOR2_X1 U765 ( .A(n707), .B(KEYINPUT59), .Z(n708) );
  XNOR2_X1 U766 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n711), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U768 ( .A1(n350), .A2(G478), .ZN(n714) );
  NOR2_X1 U769 ( .A1(n720), .A2(n715), .ZN(G63) );
  NAND2_X1 U770 ( .A1(n350), .A2(G217), .ZN(n718) );
  XNOR2_X1 U771 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U772 ( .A1(n720), .A2(n719), .ZN(G66) );
  NOR2_X1 U773 ( .A1(G898), .A2(n742), .ZN(n725) );
  XOR2_X1 U774 ( .A(G101), .B(n721), .Z(n722) );
  XNOR2_X1 U775 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n727) );
  XNOR2_X1 U777 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n726) );
  XNOR2_X1 U778 ( .A(n727), .B(n726), .ZN(n735) );
  NAND2_X1 U779 ( .A1(n609), .A2(n742), .ZN(n733) );
  XOR2_X1 U780 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n729) );
  NAND2_X1 U781 ( .A1(G224), .A2(G953), .ZN(n728) );
  XNOR2_X1 U782 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U783 ( .A1(G898), .A2(n730), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n731), .B(KEYINPUT122), .ZN(n732) );
  NAND2_X1 U785 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U786 ( .A(n735), .B(n734), .Z(G69) );
  XOR2_X1 U787 ( .A(n737), .B(n736), .Z(n739) );
  XNOR2_X1 U788 ( .A(n739), .B(n738), .ZN(n745) );
  XNOR2_X1 U789 ( .A(n745), .B(KEYINPUT125), .ZN(n740) );
  XNOR2_X1 U790 ( .A(n741), .B(n740), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U792 ( .A(n744), .B(KEYINPUT126), .ZN(n750) );
  XNOR2_X1 U793 ( .A(G227), .B(n745), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G900), .ZN(n747) );
  XOR2_X1 U795 ( .A(KEYINPUT127), .B(n747), .Z(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(G953), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n750), .A2(n749), .ZN(G72) );
  XNOR2_X1 U798 ( .A(G101), .B(n751), .ZN(G3) );
  XNOR2_X1 U799 ( .A(n752), .B(G131), .ZN(G33) );
endmodule

