//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n187));
  XNOR2_X1  g001(.A(G128), .B(G143), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT14), .A3(G122), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G122), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  OAI211_X1 g008(.A(G107), .B(new_n192), .C1(new_n194), .C2(KEYINPUT14), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n190), .B(new_n195), .C1(G107), .C2(new_n194), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(KEYINPUT13), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G128), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n197), .B(G134), .C1(KEYINPUT13), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n193), .B(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n188), .A2(new_n189), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n196), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT9), .B(G234), .Z(new_n206));
  INV_X1    g020(.A(G953), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(G217), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n205), .B(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G902), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G478), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n211), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G475), .ZN(new_n215));
  NOR2_X1   g029(.A1(G237), .A2(G953), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n216), .A2(G214), .B1(KEYINPUT86), .B2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G237), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n218), .A2(new_n207), .A3(G214), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT86), .B(G143), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT18), .A2(G131), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT87), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n219), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n218), .A2(new_n207), .A3(G214), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT86), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(new_n198), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT87), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT18), .A4(G131), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n222), .ZN(new_n232));
  INV_X1    g046(.A(G140), .ZN(new_n233));
  OAI211_X1 g047(.A(KEYINPUT74), .B(G125), .C1(new_n233), .C2(KEYINPUT75), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT74), .A2(G125), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT75), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G140), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT75), .B1(new_n233), .B2(G125), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT88), .ZN(new_n241));
  INV_X1    g055(.A(G125), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G140), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n233), .A2(G125), .ZN(new_n244));
  INV_X1    g058(.A(G146), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n239), .A2(new_n247), .A3(G146), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n241), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n231), .A2(new_n232), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT89), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT89), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n231), .A2(new_n252), .A3(new_n249), .A4(new_n232), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G131), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n228), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT17), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT16), .B1(new_n233), .B2(G125), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(new_n239), .B2(KEYINPUT16), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n245), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT16), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n233), .A2(KEYINPUT75), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n263), .A2(new_n235), .B1(new_n243), .B2(KEYINPUT75), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n262), .B1(new_n264), .B2(new_n234), .ZN(new_n265));
  OAI21_X1  g079(.A(G146), .B1(new_n265), .B2(new_n259), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n228), .A2(KEYINPUT17), .A3(G131), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n258), .A2(new_n261), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n254), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G113), .B(G122), .ZN(new_n270));
  INV_X1    g084(.A(G104), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n254), .A2(new_n272), .A3(new_n268), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n215), .B1(new_n276), .B2(new_n210), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n239), .A2(KEYINPUT19), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n243), .A2(new_n244), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n279), .B1(KEYINPUT19), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(G146), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n260), .A2(new_n245), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n256), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n239), .A2(new_n247), .A3(G146), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n247), .B1(new_n239), .B2(G146), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n288), .A2(new_n246), .B1(new_n223), .B2(new_n230), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n252), .B1(new_n289), .B2(new_n232), .ZN(new_n290));
  INV_X1    g104(.A(new_n253), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n285), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT90), .A3(new_n273), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT90), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n284), .B1(new_n251), .B2(new_n253), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(new_n272), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n296), .A3(new_n275), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT20), .ZN(new_n298));
  NOR2_X1   g112(.A1(G475), .A2(G902), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n298), .B1(new_n297), .B2(new_n299), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n214), .B(new_n278), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n207), .A2(G952), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n303), .B1(G234), .B2(G237), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XOR2_X1   g119(.A(KEYINPUT21), .B(G898), .Z(new_n306));
  NAND2_X1  g120(.A1(G234), .A2(G237), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(G902), .A3(G953), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n305), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n187), .B1(new_n302), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n297), .A2(new_n299), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT20), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n277), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n315), .A2(KEYINPUT91), .A3(new_n309), .A4(new_n214), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G116), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n191), .B2(G119), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n318), .A2(KEYINPUT67), .A3(G116), .ZN(new_n322));
  OAI211_X1 g136(.A(KEYINPUT5), .B(new_n319), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n319), .A2(KEYINPUT5), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(G113), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT67), .B1(new_n318), .B2(G116), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(new_n191), .A3(G119), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n326), .A2(new_n327), .B1(G116), .B2(new_n318), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT2), .B(G113), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(new_n271), .B2(G107), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n201), .A3(G104), .ZN(new_n335));
  INV_X1    g149(.A(G101), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n271), .A2(G107), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n333), .A2(new_n335), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n271), .A2(G107), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n201), .A2(G104), .ZN(new_n340));
  OAI21_X1  g154(.A(G101), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT85), .B1(new_n342), .B2(KEYINPUT84), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT8), .ZN(new_n345));
  XOR2_X1   g159(.A(G110), .B(G122), .Z(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n332), .A2(new_n344), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n343), .B1(KEYINPUT85), .B2(new_n342), .ZN(new_n349));
  OAI221_X1 g163(.A(new_n348), .B1(new_n345), .B2(new_n347), .C1(new_n332), .C2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n338), .A2(new_n341), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n325), .A2(new_n331), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n333), .A2(new_n335), .A3(new_n337), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G101), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n356), .A3(G101), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n328), .B(new_n329), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n352), .B(new_n347), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT81), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n328), .B(new_n330), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n355), .A3(new_n357), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n363), .A2(new_n364), .A3(new_n352), .A4(new_n347), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n198), .A2(G146), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n245), .A2(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G128), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT64), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n245), .A2(KEYINPUT64), .A3(G143), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n367), .A3(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT0), .B(G128), .Z(new_n376));
  AOI22_X1  g190(.A1(KEYINPUT0), .A2(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OR3_X1    g191(.A1(new_n369), .A2(KEYINPUT1), .A3(new_n370), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n368), .A2(KEYINPUT1), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G128), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  MUX2_X1   g196(.A(new_n377), .B(new_n382), .S(new_n242), .Z(new_n383));
  OR2_X1    g197(.A1(new_n383), .A2(KEYINPUT7), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n350), .A2(new_n366), .A3(new_n384), .ZN(new_n385));
  XOR2_X1   g199(.A(KEYINPUT82), .B(G224), .Z(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n207), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n383), .A2(new_n387), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(KEYINPUT7), .ZN(new_n390));
  AOI21_X1  g204(.A(G902), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n347), .B1(new_n363), .B2(new_n352), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n392), .A2(KEYINPUT6), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n361), .B2(new_n365), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n389), .A2(new_n388), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n397), .B1(new_n396), .B2(new_n398), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n391), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G210), .B1(G237), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n391), .B(new_n402), .C1(new_n399), .C2(new_n400), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G214), .B1(G237), .B2(G902), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G469), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n369), .A2(KEYINPUT1), .A3(new_n370), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n379), .A2(G128), .B1(new_n367), .B2(new_n368), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n351), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n382), .B2(new_n351), .ZN(new_n413));
  INV_X1    g227(.A(G137), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT65), .B1(new_n414), .B2(G134), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT65), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n189), .A3(G137), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT11), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n189), .B2(G137), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(KEYINPUT11), .A3(G134), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n418), .A2(new_n255), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n420), .A2(new_n421), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n255), .B1(new_n424), .B2(new_n418), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n413), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT12), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT12), .B1(new_n413), .B2(new_n427), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT10), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n412), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n382), .A2(KEYINPUT10), .A3(new_n351), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n377), .A2(new_n355), .A3(new_n357), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n434), .A2(new_n426), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n207), .A2(G227), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT80), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n427), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n441), .B1(new_n445), .B2(new_n437), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n409), .B(new_n210), .C1(new_n443), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(G469), .A2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n441), .ZN(new_n449));
  INV_X1    g263(.A(new_n437), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n449), .B1(new_n432), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n442), .B1(new_n427), .B2(new_n444), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n453), .A3(G469), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n447), .A2(new_n448), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n206), .A2(new_n210), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G221), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT79), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n408), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT66), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n414), .B2(G134), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n414), .A2(G134), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n189), .A2(KEYINPUT66), .A3(G137), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G131), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n422), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n422), .A2(KEYINPUT68), .A3(new_n468), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n382), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n377), .B1(new_n423), .B2(new_n425), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n422), .A2(new_n468), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n382), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n474), .A2(new_n477), .A3(new_n462), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n362), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n382), .A2(new_n472), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT68), .B1(new_n422), .B2(new_n468), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n474), .B(new_n359), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n216), .A2(G210), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(new_n336), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n484), .B(new_n485), .Z(new_n486));
  NAND3_X1  g300(.A1(new_n479), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT31), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n482), .A2(KEYINPUT28), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT28), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n473), .A2(new_n490), .A3(new_n359), .A4(new_n474), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n474), .A2(new_n477), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n362), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n486), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n479), .A2(new_n498), .A3(new_n482), .A4(new_n486), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n488), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G472), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n210), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n495), .A2(new_n486), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n479), .A2(new_n482), .A3(new_n496), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT29), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n359), .B1(new_n473), .B2(new_n474), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n489), .B2(new_n491), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT29), .A3(new_n486), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n210), .ZN(new_n511));
  OAI21_X1  g325(.A(G472), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n500), .A2(KEYINPUT32), .A3(new_n501), .A4(new_n210), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT32), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n502), .A2(KEYINPUT69), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n504), .A2(new_n512), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n207), .A2(G221), .A3(G234), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT76), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT22), .B(G137), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT77), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT71), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n524), .B1(new_n318), .B2(G128), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n318), .A2(G128), .ZN(new_n526));
  MUX2_X1   g340(.A(new_n525), .B(new_n524), .S(new_n526), .Z(new_n527));
  XOR2_X1   g341(.A(KEYINPUT24), .B(G110), .Z(new_n528));
  NAND3_X1  g342(.A1(new_n370), .A2(KEYINPUT23), .A3(G119), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n530), .B1(new_n318), .B2(G128), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n529), .B1(new_n531), .B2(new_n526), .ZN(new_n532));
  OAI22_X1  g346(.A1(new_n527), .A2(new_n528), .B1(G110), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n266), .A3(new_n246), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(KEYINPUT72), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT72), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n536), .B(new_n529), .C1(new_n531), .C2(new_n526), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(G110), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT73), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n535), .A2(KEYINPUT73), .A3(G110), .A4(new_n537), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n527), .A2(new_n528), .ZN(new_n543));
  AOI211_X1 g357(.A(G146), .B(new_n259), .C1(new_n239), .C2(KEYINPUT16), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n543), .B1(new_n283), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n523), .B(new_n534), .C1(new_n542), .C2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n266), .A2(new_n261), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n548), .A2(new_n543), .A3(new_n540), .A4(new_n541), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n523), .B1(new_n549), .B2(new_n534), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n522), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n534), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT77), .ZN(new_n553));
  INV_X1    g367(.A(new_n522), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n551), .A2(new_n210), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT78), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(KEYINPUT25), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G217), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(G234), .B2(new_n210), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n551), .A2(new_n555), .A3(new_n210), .A4(new_n558), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n551), .A2(new_n555), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n562), .A2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n317), .A2(new_n461), .A3(new_n518), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  NAND2_X1  g385(.A1(new_n500), .A2(new_n210), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G472), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n502), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n574), .A2(new_n568), .A3(new_n460), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n575), .B(KEYINPUT92), .Z(new_n576));
  INV_X1    g390(.A(new_n407), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n404), .B2(new_n405), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n278), .B1(new_n300), .B2(new_n301), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n205), .A2(new_n208), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT33), .B1(new_n580), .B2(KEYINPUT93), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(new_n209), .ZN(new_n582));
  OAI21_X1  g396(.A(G478), .B1(new_n582), .B2(G902), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n211), .A2(G478), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(new_n310), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n576), .A2(new_n578), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT34), .B(G104), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G6));
  INV_X1    g404(.A(new_n214), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n591), .B(new_n278), .C1(new_n300), .C2(new_n301), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n309), .B(KEYINPUT94), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n408), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n576), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT95), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT35), .B(G107), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G9));
  NOR2_X1   g412(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n552), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n566), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n564), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  OR3_X1    g417(.A1(new_n603), .A2(new_n574), .A3(KEYINPUT96), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT96), .B1(new_n603), .B2(new_n574), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n317), .A2(new_n461), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G110), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n606), .B(new_n608), .ZN(G12));
  AOI221_X4 g423(.A(new_n577), .B1(new_n564), .B2(new_n601), .C1(new_n404), .C2(new_n405), .ZN(new_n610));
  INV_X1    g424(.A(new_n460), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n304), .B(KEYINPUT98), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(G900), .B2(new_n308), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n592), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n518), .A2(new_n610), .A3(new_n611), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G128), .ZN(G30));
  NOR2_X1   g432(.A1(new_n315), .A2(new_n214), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n614), .B(KEYINPUT39), .Z(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n455), .A2(new_n459), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n619), .B1(new_n624), .B2(KEYINPUT40), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n622), .A2(new_n623), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n622), .A2(new_n623), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n602), .A2(new_n577), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n496), .B1(new_n479), .B2(new_n482), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n482), .A2(new_n496), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n210), .B1(new_n633), .B2(new_n508), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n504), .A2(new_n515), .A3(new_n517), .A4(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n406), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n638), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n406), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n630), .A2(new_n631), .A3(new_n636), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G143), .ZN(G45));
  NAND3_X1  g458(.A1(new_n518), .A2(new_n610), .A3(new_n611), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n579), .A2(new_n585), .A3(new_n614), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n579), .A2(KEYINPUT101), .A3(new_n585), .A4(new_n614), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(new_n245), .ZN(G48));
  NAND3_X1  g466(.A1(new_n587), .A2(new_n518), .A3(new_n569), .ZN(new_n653));
  INV_X1    g467(.A(new_n446), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n654), .B1(new_n432), .B2(new_n442), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n210), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(G469), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n447), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n458), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n578), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT41), .B(G113), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT102), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G15));
  AOI211_X1 g478(.A(new_n577), .B(new_n593), .C1(new_n404), .C2(new_n405), .ZN(new_n665));
  INV_X1    g479(.A(new_n592), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n518), .A2(new_n665), .A3(new_n569), .A4(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n660), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n191), .ZN(G18));
  AND3_X1   g483(.A1(new_n578), .A2(new_n602), .A3(new_n659), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n317), .A3(new_n518), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT103), .ZN(new_n672));
  AOI211_X1 g486(.A(new_n514), .B(new_n516), .C1(new_n502), .C2(KEYINPUT69), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n517), .A2(new_n515), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI22_X1  g489(.A1(new_n675), .A2(new_n512), .B1(new_n311), .B2(new_n316), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n670), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G119), .ZN(G21));
  AOI21_X1  g494(.A(KEYINPUT105), .B1(new_n572), .B2(G472), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n682));
  AOI211_X1 g496(.A(new_n682), .B(new_n501), .C1(new_n500), .C2(new_n210), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n488), .B(new_n499), .C1(new_n486), .C2(new_n509), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n501), .A3(new_n210), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n685), .A2(KEYINPUT104), .A3(new_n501), .A4(new_n210), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n569), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n660), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n315), .A2(new_n214), .A3(new_n593), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G122), .ZN(G24));
  NAND4_X1  g511(.A1(new_n670), .A2(new_n648), .A3(new_n649), .A4(new_n691), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT106), .B(G125), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G27));
  NOR3_X1   g514(.A1(new_n406), .A2(new_n577), .A3(new_n460), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n518), .A3(new_n569), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n648), .A2(new_n704), .A3(new_n649), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n502), .A2(new_n516), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n512), .A3(new_n513), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n707), .A2(new_n569), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n648), .A2(new_n708), .A3(new_n701), .A4(new_n649), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n703), .A2(new_n705), .B1(new_n709), .B2(KEYINPUT42), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G131), .ZN(G33));
  AOI21_X1  g525(.A(new_n568), .B1(new_n675), .B2(new_n512), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n713), .B1(new_n592), .B2(new_n615), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n315), .A2(KEYINPUT107), .A3(new_n591), .A4(new_n614), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n712), .A2(KEYINPUT108), .A3(new_n716), .A4(new_n701), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n715), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n702), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n574), .A2(new_n602), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n315), .A2(new_n585), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT43), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n315), .A2(new_n729), .A3(new_n585), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n723), .B1(new_n726), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n724), .B(KEYINPUT110), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(KEYINPUT44), .A3(new_n728), .A4(new_n730), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n428), .B(new_n429), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n441), .B1(new_n736), .B2(new_n437), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n735), .B1(new_n737), .B2(new_n452), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n451), .A2(new_n453), .A3(KEYINPUT45), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(G469), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(KEYINPUT46), .A3(new_n448), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n447), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT46), .B1(new_n740), .B2(new_n448), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n459), .B(new_n621), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT109), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n406), .A2(new_n577), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n732), .A2(new_n734), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT111), .B(G137), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G39));
  OAI21_X1  g563(.A(new_n459), .B1(new_n742), .B2(new_n743), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT47), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n752), .B(new_n459), .C1(new_n742), .C2(new_n743), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n650), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n518), .A2(new_n569), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n746), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G140), .ZN(G42));
  INV_X1    g572(.A(new_n642), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n658), .A2(KEYINPUT49), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n658), .A2(KEYINPUT49), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n569), .A3(new_n761), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n762), .A2(new_n577), .A3(new_n727), .ZN(new_n763));
  INV_X1    g577(.A(new_n636), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n759), .A2(new_n763), .A3(new_n459), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n648), .A2(new_n691), .A3(new_n649), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n578), .A2(new_n602), .A3(new_n659), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n617), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n651), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n564), .A2(new_n601), .A3(new_n614), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n460), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n636), .A2(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n619), .A3(new_n578), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n769), .A2(new_n770), .A3(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n698), .B(new_n617), .C1(new_n650), .C2(new_n645), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT52), .B1(new_n780), .B2(new_n777), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n712), .B(new_n694), .C1(new_n587), .C2(new_n594), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n677), .B1(new_n676), .B2(new_n670), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n677), .A2(new_n670), .A3(new_n317), .A4(new_n518), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n786), .B(new_n696), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n586), .A2(new_n592), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n665), .A3(new_n575), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n606), .A2(new_n570), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n606), .A2(new_n570), .A3(new_n792), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT112), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n789), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n770), .B1(new_n769), .B2(new_n778), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n518), .A2(new_n214), .A3(new_n315), .A4(new_n614), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n766), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n602), .A3(new_n701), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n721), .A2(new_n800), .A3(new_n710), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n768), .A2(new_n651), .A3(new_n777), .A4(KEYINPUT52), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n797), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n785), .A2(new_n796), .A3(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n721), .A2(new_n800), .A3(new_n710), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n779), .A3(new_n781), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n795), .A2(new_n793), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n660), .B1(new_n667), .B2(new_n653), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n678), .B2(new_n672), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n696), .A3(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n784), .B(new_n783), .C1(new_n806), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n804), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT54), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n731), .A2(new_n613), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n693), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n639), .A2(new_n577), .A3(new_n641), .A4(new_n659), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT117), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT50), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  OAI211_X1 g633(.A(KEYINPUT117), .B(new_n819), .C1(new_n815), .C2(new_n816), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n746), .A2(new_n659), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n569), .A3(new_n304), .A4(new_n764), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n823), .A2(new_n579), .A3(new_n585), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n814), .A2(new_n602), .A3(new_n691), .A4(new_n822), .ZN(new_n825));
  INV_X1    g639(.A(new_n746), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n658), .A2(new_n459), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(KEYINPUT116), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(KEYINPUT116), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n754), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n827), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n821), .A2(new_n824), .A3(new_n825), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n823), .A2(new_n586), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n303), .A2(KEYINPUT118), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n303), .A2(KEYINPUT118), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n814), .A2(new_n708), .A3(new_n822), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT48), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT48), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n814), .A2(new_n842), .A3(new_n708), .A4(new_n822), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n814), .A2(new_n694), .A3(new_n693), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n839), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n839), .A2(new_n844), .A3(KEYINPUT119), .A4(new_n845), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n754), .B1(new_n459), .B2(new_n658), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n834), .B1(new_n827), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n821), .A2(new_n852), .A3(new_n824), .A4(new_n825), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n835), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT120), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n809), .A2(new_n856), .A3(new_n696), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n789), .A2(KEYINPUT115), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n784), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n803), .A3(new_n807), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n784), .B1(new_n806), .B2(new_n810), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n835), .A2(new_n850), .A3(new_n864), .A4(new_n853), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n813), .A2(new_n855), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(G952), .A2(G953), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n765), .B1(new_n866), .B2(new_n867), .ZN(G75));
  NAND2_X1  g682(.A1(new_n860), .A2(new_n861), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(G210), .A3(G902), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n396), .B(new_n398), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT55), .Z(new_n873));
  AND3_X1   g687(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n870), .B2(new_n871), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n207), .A2(G952), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(G51));
  NAND2_X1  g691(.A1(new_n448), .A2(KEYINPUT57), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n448), .A2(KEYINPUT57), .ZN(new_n879));
  INV_X1    g693(.A(new_n863), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n862), .B1(new_n860), .B2(new_n861), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n878), .B(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n655), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n856), .B1(new_n809), .B2(new_n696), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n789), .A2(KEYINPUT115), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT53), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n805), .A2(new_n807), .A3(new_n779), .A4(new_n781), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT53), .B1(new_n803), .B2(new_n796), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n890), .A2(new_n210), .A3(new_n740), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n876), .B1(new_n883), .B2(new_n891), .ZN(G54));
  NAND4_X1  g706(.A1(new_n869), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n893));
  INV_X1    g707(.A(new_n297), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n895), .A2(new_n896), .A3(new_n876), .ZN(G60));
  INV_X1    g711(.A(new_n876), .ZN(new_n898));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT59), .Z(new_n900));
  NOR2_X1   g714(.A1(new_n582), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n880), .B2(new_n881), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n813), .B2(new_n863), .ZN(new_n903));
  INV_X1    g717(.A(new_n582), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n898), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(G63));
  NAND2_X1  g720(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT121), .Z(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT60), .Z(new_n913));
  OAI211_X1 g727(.A(new_n600), .B(new_n913), .C1(new_n888), .C2(new_n889), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n898), .ZN(new_n915));
  INV_X1    g729(.A(new_n913), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n860), .B2(new_n861), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n565), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n907), .B(new_n910), .C1(new_n915), .C2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n565), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n890), .B2(new_n916), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n876), .B1(new_n917), .B2(new_n600), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n922), .A3(new_n908), .A4(new_n909), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n919), .A2(new_n923), .ZN(G66));
  AOI21_X1  g738(.A(new_n207), .B1(new_n306), .B2(new_n386), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n810), .B2(new_n207), .ZN(new_n926));
  INV_X1    g740(.A(new_n396), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(G898), .B2(new_n207), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n926), .B(new_n928), .Z(G69));
  AOI21_X1  g743(.A(new_n207), .B1(G227), .B2(G900), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n930), .A2(KEYINPUT126), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n475), .A2(new_n478), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(new_n281), .Z(new_n933));
  NOR2_X1   g747(.A1(new_n826), .A2(new_n624), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n712), .A3(new_n791), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(KEYINPUT124), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(KEYINPUT124), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n747), .B(new_n757), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n768), .B2(new_n651), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n518), .A2(new_n610), .A3(new_n611), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n648), .A2(new_n649), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n943), .A2(KEYINPUT123), .A3(new_n617), .A4(new_n698), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n940), .A2(new_n944), .A3(new_n643), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n940), .A2(new_n944), .A3(new_n643), .A4(KEYINPUT62), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n938), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n933), .B1(new_n949), .B2(G953), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(KEYINPUT125), .B(new_n933), .C1(new_n949), .C2(G953), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n930), .A2(KEYINPUT126), .ZN(new_n955));
  AND4_X1   g769(.A1(new_n710), .A2(new_n747), .A3(new_n757), .A4(new_n721), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n940), .A2(new_n944), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n745), .A2(new_n578), .A3(new_n619), .A4(new_n708), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n956), .A2(new_n957), .A3(new_n207), .A4(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n933), .ZN(new_n960));
  NAND2_X1  g774(.A1(G900), .A2(G953), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n931), .A2(new_n954), .A3(new_n955), .A4(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n952), .B2(new_n953), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n931), .B1(new_n965), .B2(new_n955), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n963), .A2(new_n966), .ZN(G72));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  NAND3_X1  g783(.A1(new_n956), .A2(new_n958), .A3(new_n957), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n810), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n506), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n972), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n949), .A2(new_n796), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n969), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n876), .B1(new_n978), .B2(new_n632), .ZN(new_n979));
  INV_X1    g793(.A(new_n632), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n812), .A2(new_n506), .A3(new_n980), .A4(new_n969), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n976), .A2(new_n979), .A3(new_n981), .ZN(G57));
endmodule


