//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT2), .ZN(new_n187));
  INV_X1    g001(.A(G113), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(KEYINPUT64), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n190), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT2), .A2(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT2), .A3(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G116), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G119), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n199), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n203), .A3(new_n199), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n198), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n191), .A2(new_n189), .B1(new_n194), .B2(new_n196), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n201), .A2(new_n203), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT0), .B(G128), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT11), .ZN(new_n222));
  INV_X1    g036(.A(G134), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(G137), .ZN(new_n224));
  INV_X1    g038(.A(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT11), .A3(G134), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(G137), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n224), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(new_n226), .A3(new_n228), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n221), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n215), .B2(G146), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n215), .A2(G146), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n213), .A2(G143), .ZN(new_n235));
  OAI211_X1 g049(.A(G128), .B(new_n233), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n214), .B(new_n216), .C1(KEYINPUT1), .C2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n223), .A2(G137), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n225), .A2(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(G131), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND4_X1   g055(.A1(new_n229), .A2(new_n236), .A3(new_n238), .A4(new_n241), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n232), .A2(new_n242), .A3(KEYINPUT30), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT30), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n231), .A2(new_n229), .ZN(new_n245));
  INV_X1    g059(.A(new_n221), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n236), .A2(new_n229), .A3(new_n241), .A4(new_n238), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n212), .B1(new_n243), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n247), .A2(new_n207), .A3(new_n211), .A4(new_n248), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT67), .B(KEYINPUT31), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n250), .A2(new_n251), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n256), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n212), .B1(new_n232), .B2(new_n242), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n251), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n232), .A2(new_n242), .ZN(new_n263));
  INV_X1    g077(.A(new_n212), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT28), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n259), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT30), .B1(new_n232), .B2(new_n242), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n247), .A2(new_n244), .A3(new_n248), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n212), .A2(new_n232), .A3(new_n242), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n269), .A2(new_n270), .A3(new_n259), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT31), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n258), .B(new_n266), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(G472), .A2(G902), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT32), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n274), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n276), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n247), .A2(new_n248), .B1(new_n207), .B2(new_n211), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT28), .B1(new_n270), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n251), .A2(new_n260), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n256), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n259), .B1(new_n269), .B2(new_n270), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n265), .B1(new_n262), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n259), .A2(new_n288), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT69), .B(G902), .Z(new_n295));
  NAND3_X1  g109(.A1(new_n289), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G472), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n273), .A2(KEYINPUT70), .A3(new_n277), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n280), .A2(new_n282), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n300), .A2(KEYINPUT16), .A3(G140), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT16), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n302), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n213), .ZN(new_n309));
  XNOR2_X1  g123(.A(G125), .B(G140), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n301), .B1(new_n310), .B2(KEYINPUT16), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G146), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n200), .B2(G128), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n237), .A2(KEYINPUT23), .A3(G119), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n315), .B(new_n316), .C1(G119), .C2(new_n237), .ZN(new_n317));
  XNOR2_X1  g131(.A(G119), .B(G128), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT24), .B(G110), .Z(new_n319));
  AOI22_X1  g133(.A1(new_n317), .A2(G110), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n306), .A2(G146), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n311), .B2(G146), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT72), .B(G110), .Z(new_n324));
  OAI22_X1  g138(.A1(new_n317), .A2(new_n324), .B1(new_n318), .B2(new_n319), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(KEYINPUT73), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT73), .B1(new_n323), .B2(new_n325), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n321), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G221), .A3(G234), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT74), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT22), .B(G137), .Z(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n334), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n323), .A2(new_n325), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n326), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n336), .B1(new_n340), .B2(new_n321), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n295), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n329), .A2(new_n334), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n340), .A2(new_n321), .A3(new_n336), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT25), .A3(new_n295), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G217), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n295), .B2(G234), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n351), .B(KEYINPUT71), .Z(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n351), .A2(G902), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n349), .A2(new_n353), .B1(new_n354), .B2(new_n347), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n299), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G469), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(new_n231), .B2(new_n229), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n236), .A2(new_n238), .ZN(new_n361));
  INV_X1    g175(.A(G104), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G107), .ZN(new_n363));
  INV_X1    g177(.A(G101), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G107), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT76), .A3(G104), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n366), .A2(KEYINPUT76), .A3(KEYINPUT3), .A4(G104), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n365), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n366), .A2(G104), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n362), .A2(G107), .ZN(new_n373));
  OAI21_X1  g187(.A(G101), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n361), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n365), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT3), .B1(new_n373), .B2(KEYINPUT76), .ZN(new_n378));
  INV_X1    g192(.A(new_n370), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n380), .A2(new_n374), .B1(new_n238), .B2(new_n236), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n360), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT12), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT12), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n360), .B(new_n384), .C1(new_n376), .C2(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n372), .B1(new_n369), .B2(new_n370), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n380), .B(KEYINPUT4), .C1(new_n387), .C2(new_n364), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n363), .B1(new_n378), .B2(new_n379), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n364), .A2(KEYINPUT4), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n221), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT10), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n380), .A2(new_n374), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n361), .ZN(new_n395));
  INV_X1    g209(.A(new_n245), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n371), .A2(new_n375), .ZN(new_n397));
  INV_X1    g211(.A(new_n361), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT10), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n395), .A3(new_n396), .A4(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G110), .B(G140), .ZN(new_n401));
  INV_X1    g215(.A(G227), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G953), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n401), .B(new_n403), .Z(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n386), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n392), .A2(new_n395), .A3(new_n399), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n245), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n404), .B1(new_n408), .B2(new_n400), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n358), .B(new_n295), .C1(new_n406), .C2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G902), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n358), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n383), .A2(new_n400), .A3(new_n385), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n404), .B(KEYINPUT75), .Z(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n408), .A2(new_n400), .A3(new_n404), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n410), .B(new_n413), .C1(new_n358), .C2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT9), .B(G234), .ZN(new_n420));
  OAI21_X1  g234(.A(G221), .B1(new_n420), .B2(G902), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G478), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT15), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n202), .A2(G122), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n366), .B1(new_n426), .B2(KEYINPUT14), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n202), .A2(G122), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n427), .B(new_n429), .Z(new_n430));
  XNOR2_X1  g244(.A(G128), .B(G143), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT90), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n432), .A2(new_n223), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n223), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n223), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(KEYINPUT13), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n215), .A2(G128), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n437), .B(G134), .C1(KEYINPUT13), .C2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT89), .B(G107), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n429), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n429), .A2(new_n440), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n436), .A2(new_n439), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n420), .A2(new_n350), .A3(G953), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n435), .A2(new_n443), .A3(new_n445), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n425), .B1(new_n449), .B2(new_n295), .ZN(new_n450));
  INV_X1    g264(.A(new_n295), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n451), .B(new_n424), .C1(new_n447), .C2(new_n448), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n306), .A2(KEYINPUT84), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n304), .A2(new_n305), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(G146), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n458));
  INV_X1    g272(.A(new_n322), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(KEYINPUT18), .A2(G131), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n252), .A2(G143), .A3(G214), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(G143), .B1(new_n252), .B2(G214), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G237), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n330), .A3(G214), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n215), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(KEYINPUT18), .A3(G131), .A4(new_n462), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n460), .A2(new_n470), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n304), .A2(new_n305), .A3(new_n455), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n455), .B1(new_n304), .B2(new_n305), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n472), .A2(new_n473), .A3(new_n213), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT85), .B1(new_n474), .B2(new_n322), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n468), .A2(new_n227), .A3(new_n462), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT86), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT17), .ZN(new_n478));
  OAI21_X1  g292(.A(G131), .B1(new_n463), .B2(new_n464), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT86), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n468), .A2(new_n480), .A3(new_n227), .A4(new_n462), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(KEYINPUT17), .B(G131), .C1(new_n463), .C2(new_n464), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n309), .A2(new_n312), .A3(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n471), .A2(new_n475), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G113), .B(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n362), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n485), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n411), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT88), .B(G475), .Z(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(G475), .A2(G902), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n475), .A2(new_n460), .A3(new_n470), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n454), .A2(KEYINPUT19), .A3(new_n456), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n306), .A2(KEYINPUT19), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n213), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n312), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT87), .ZN(new_n500));
  INV_X1    g314(.A(new_n487), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n484), .A2(new_n482), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n493), .A3(new_n487), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n487), .B1(new_n493), .B2(new_n498), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(new_n500), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n492), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(KEYINPUT20), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT20), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n499), .A2(new_n501), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT87), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n504), .A3(new_n502), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n510), .B1(new_n513), .B2(new_n492), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n453), .B(new_n491), .C1(new_n509), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n330), .A2(G952), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(G234), .B2(G237), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n330), .B(new_n295), .C1(G234), .C2(G237), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT21), .B(G898), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n422), .A2(new_n515), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(G110), .B(G122), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT8), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n201), .A2(new_n203), .A3(new_n199), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT5), .B1(new_n525), .B2(new_n204), .ZN(new_n526));
  INV_X1    g340(.A(new_n201), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT5), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n188), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n526), .A2(new_n529), .B1(new_n210), .B2(new_n208), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n530), .A2(new_n397), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n531), .A2(KEYINPUT81), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n529), .B1(new_n528), .B2(new_n209), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n397), .A2(new_n211), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(new_n531), .B2(KEYINPUT81), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n524), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n221), .A2(G125), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n398), .B2(G125), .ZN(new_n538));
  INV_X1    g352(.A(G224), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT7), .B1(new_n539), .B2(G953), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n538), .B(new_n540), .Z(new_n541));
  NAND2_X1  g355(.A1(new_n389), .A2(new_n390), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n388), .A2(new_n212), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n530), .A2(new_n397), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n522), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n411), .B1(new_n536), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n207), .A2(new_n211), .B1(new_n389), .B2(new_n390), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n548), .A2(new_n388), .B1(new_n530), .B2(new_n397), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n549), .A2(KEYINPUT6), .A3(new_n522), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT79), .B1(new_n549), .B2(new_n522), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT6), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n549), .B2(new_n522), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n543), .A2(new_n544), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT79), .ZN(new_n555));
  INV_X1    g369(.A(new_n522), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT80), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n551), .A2(new_n553), .A3(new_n557), .A4(KEYINPUT80), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n550), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n539), .A2(G953), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n538), .B(new_n563), .Z(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n547), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G210), .B1(G237), .B2(G902), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT82), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n550), .ZN(new_n569));
  AOI211_X1 g383(.A(KEYINPUT79), .B(new_n522), .C1(new_n543), .C2(new_n544), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n545), .A2(KEYINPUT6), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT80), .B1(new_n572), .B2(new_n551), .ZN(new_n573));
  INV_X1    g387(.A(new_n561), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n569), .B(new_n565), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n547), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n567), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT82), .ZN(new_n578));
  INV_X1    g392(.A(new_n567), .ZN(new_n579));
  AOI211_X1 g393(.A(new_n550), .B(new_n564), .C1(new_n560), .C2(new_n561), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n547), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n568), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT83), .ZN(new_n583));
  OAI21_X1  g397(.A(G214), .B1(G237), .B2(G902), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n584), .B(KEYINPUT78), .Z(new_n585));
  AND3_X1   g399(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n583), .B1(new_n582), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n357), .B(new_n521), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n347), .A2(new_n354), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT25), .B1(new_n347), .B2(new_n295), .ZN(new_n592));
  AOI211_X1 g406(.A(new_n343), .B(new_n451), .C1(new_n345), .C2(new_n346), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n353), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n419), .A2(new_n591), .A3(new_n594), .A4(new_n421), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n273), .A2(new_n295), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n596), .A2(G472), .B1(new_n273), .B2(new_n274), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n590), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n421), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n416), .A2(new_n417), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n412), .B1(new_n601), .B2(G469), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n600), .B1(new_n602), .B2(new_n410), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n603), .A2(new_n597), .A3(KEYINPUT91), .A4(new_n355), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n547), .B(new_n579), .C1(new_n562), .C2(new_n565), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n567), .B1(new_n575), .B2(new_n576), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n584), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n491), .B1(new_n509), .B2(new_n514), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT92), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n610), .B1(new_n448), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n449), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n447), .B(new_n448), .C1(new_n611), .C2(new_n610), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n451), .A2(new_n423), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n449), .A2(new_n295), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n423), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  NOR4_X1   g435(.A1(new_n605), .A2(new_n520), .A3(new_n608), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n584), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n579), .B1(new_n580), .B2(new_n547), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n626), .B2(new_n577), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT93), .ZN(new_n628));
  INV_X1    g442(.A(new_n490), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n488), .B2(new_n411), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n508), .A2(KEYINPUT20), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n513), .A2(new_n510), .A3(new_n492), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n453), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n628), .B1(new_n635), .B2(new_n520), .ZN(new_n636));
  INV_X1    g450(.A(new_n520), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n633), .A2(KEYINPUT93), .A3(new_n637), .A4(new_n634), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n627), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n605), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT35), .B(G107), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  INV_X1    g456(.A(KEYINPUT36), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n334), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT94), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n329), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n644), .B(KEYINPUT94), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n329), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n349), .A2(new_n353), .B1(new_n354), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n598), .A2(new_n652), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n521), .B(new_n653), .C1(new_n586), .C2(new_n587), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n354), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n594), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n299), .A2(new_n603), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n517), .B1(new_n518), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n633), .A2(new_n634), .A3(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n608), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n237), .ZN(G30));
  OR2_X1    g479(.A1(new_n582), .A2(KEYINPUT38), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n582), .A2(KEYINPUT38), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n269), .A2(new_n270), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n259), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n251), .A2(new_n261), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n411), .B1(new_n671), .B2(new_n256), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n280), .A2(new_n282), .A3(new_n298), .A4(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n633), .A2(new_n453), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n658), .A2(new_n625), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n661), .B(KEYINPUT39), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n603), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n675), .B(new_n676), .C1(new_n678), .C2(KEYINPUT40), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(KEYINPUT40), .B2(new_n678), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n668), .A2(new_n674), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  AOI22_X1  g496(.A1(new_n615), .A2(new_n616), .B1(new_n423), .B2(new_n618), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n633), .A2(new_n683), .A3(new_n661), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n684), .B(new_n584), .C1(new_n606), .C2(new_n607), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT95), .B1(new_n685), .B2(new_n659), .ZN(new_n686));
  INV_X1    g500(.A(new_n659), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT95), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(new_n627), .A3(new_n688), .A4(new_n684), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  OAI21_X1  g505(.A(new_n295), .B1(new_n406), .B2(new_n409), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n421), .A3(new_n410), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT96), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n693), .A2(KEYINPUT96), .A3(new_n421), .A4(new_n410), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n299), .A2(new_n696), .A3(new_n355), .A4(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n621), .A2(new_n520), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n627), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT41), .B(G113), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT97), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n700), .B(new_n702), .ZN(G15));
  NAND4_X1  g517(.A1(new_n698), .A2(new_n627), .A3(new_n638), .A4(new_n636), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  AND2_X1   g519(.A1(new_n696), .A2(new_n697), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n515), .A2(new_n652), .A3(new_n520), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n627), .A2(new_n706), .A3(new_n707), .A4(new_n299), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  AND3_X1   g523(.A1(new_n696), .A2(new_n637), .A3(new_n697), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n291), .A2(new_n292), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n256), .B1(new_n711), .B2(KEYINPUT98), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT98), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n291), .A2(new_n292), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n258), .B1(new_n271), .B2(new_n272), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n275), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n596), .A2(G472), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n594), .A2(new_n591), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n710), .A2(new_n627), .A3(new_n675), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NAND2_X1  g537(.A1(new_n596), .A2(G472), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n716), .B1(new_n712), .B2(new_n714), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n658), .B(new_n724), .C1(new_n275), .C2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n609), .A2(new_n620), .A3(new_n662), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n627), .A3(new_n706), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT99), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n728), .A2(new_n627), .A3(KEYINPUT99), .A4(new_n706), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n625), .B1(new_n566), .B2(new_n567), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n568), .A2(new_n736), .A3(new_n581), .A4(new_n603), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n296), .A2(G472), .B1(new_n273), .B2(new_n277), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n720), .B1(new_n282), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n684), .A3(KEYINPUT42), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n735), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n568), .A2(new_n736), .A3(new_n581), .A4(new_n603), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n743), .A2(new_n740), .A3(KEYINPUT100), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n356), .A3(new_n727), .ZN(new_n745));
  OAI22_X1  g559(.A1(new_n742), .A2(new_n744), .B1(new_n745), .B2(KEYINPUT42), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NOR2_X1   g561(.A1(new_n743), .A2(new_n356), .ZN(new_n748));
  INV_X1    g562(.A(new_n663), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  AND2_X1   g565(.A1(new_n601), .A2(KEYINPUT45), .ZN(new_n752));
  OAI21_X1  g566(.A(G469), .B1(new_n601), .B2(KEYINPUT45), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n412), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(KEYINPUT46), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n410), .B1(new_n755), .B2(KEYINPUT46), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n421), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n677), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n568), .A2(new_n736), .A3(new_n581), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n652), .A2(new_n597), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT101), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n620), .A2(new_n633), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT43), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n762), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n764), .A2(new_n766), .A3(new_n762), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n761), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  XNOR2_X1  g584(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n758), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(KEYINPUT102), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n758), .B2(new_n775), .ZN(new_n776));
  OR4_X1    g590(.A1(new_n299), .A2(new_n760), .A3(new_n355), .A4(new_n727), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n303), .ZN(G42));
  NAND2_X1  g593(.A1(new_n696), .A2(new_n697), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n760), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT114), .ZN(new_n782));
  INV_X1    g596(.A(new_n517), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n674), .A2(new_n720), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(new_n633), .A3(new_n683), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n693), .A2(new_n410), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT111), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT111), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n600), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n776), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n760), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n355), .B(new_n724), .C1(new_n275), .C2(new_n725), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n766), .A2(KEYINPUT110), .A3(new_n783), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT110), .B1(new_n766), .B2(new_n783), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n718), .A2(new_n652), .A3(new_n719), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n795), .A2(new_n796), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n782), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n801), .B1(new_n782), .B2(new_n800), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n787), .A2(new_n798), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n666), .A2(new_n625), .A3(new_n667), .A4(new_n706), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n797), .B1(new_n807), .B2(KEYINPUT112), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n807), .A2(KEYINPUT112), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n806), .B(KEYINPUT50), .C1(new_n808), .C2(new_n809), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT109), .B1(new_n805), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT51), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n817));
  OAI211_X1 g631(.A(KEYINPUT109), .B(new_n817), .C1(new_n805), .C2(new_n814), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n739), .B1(new_n802), .B2(new_n803), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT48), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n609), .A2(new_n782), .A3(new_n620), .A4(new_n784), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n608), .A2(new_n780), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n516), .B(new_n822), .C1(new_n823), .C2(new_n797), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n820), .B2(new_n824), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n816), .B(new_n818), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n664), .B1(new_n686), .B2(new_n689), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n584), .B(new_n675), .C1(new_n606), .C2(new_n607), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n422), .A2(new_n658), .A3(new_n661), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n674), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n829), .A2(new_n733), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT105), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n829), .A2(new_n733), .A3(KEYINPUT52), .A4(new_n833), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n834), .A2(KEYINPUT105), .A3(new_n835), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n704), .A2(new_n700), .A3(new_n722), .A4(new_n708), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT103), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n599), .A2(new_n604), .A3(new_n637), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n635), .A2(KEYINPUT104), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT104), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n633), .A2(new_n847), .A3(new_n634), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n846), .A2(new_n621), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n586), .B2(new_n587), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n588), .A2(new_n654), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n799), .A2(new_n603), .A3(new_n684), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n515), .A2(new_n661), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n299), .A3(new_n603), .A4(new_n658), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n793), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n750), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n745), .A2(KEYINPUT42), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n737), .A2(new_n741), .A3(new_n735), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT100), .B1(new_n743), .B2(new_n740), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n858), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n844), .A2(new_n852), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n828), .B1(new_n841), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT107), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n836), .A2(new_n838), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n707), .A2(new_n299), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n696), .A2(new_n637), .A3(new_n697), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n794), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n823), .A2(new_n868), .B1(new_n831), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n843), .A3(new_n700), .A4(new_n704), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n842), .A2(KEYINPUT103), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n749), .A2(new_n748), .B1(new_n856), .B2(new_n793), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n746), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n867), .A2(new_n875), .A3(new_n852), .ZN(new_n876));
  XNOR2_X1  g690(.A(KEYINPUT106), .B(KEYINPUT53), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n866), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(new_n873), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n746), .A2(new_n874), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n588), .A2(new_n654), .A3(new_n851), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n877), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n882), .A2(KEYINPUT107), .A3(new_n867), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n865), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n842), .A2(new_n828), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n880), .A2(new_n881), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n839), .A3(new_n840), .ZN(new_n889));
  AOI211_X1 g703(.A(KEYINPUT108), .B(new_n883), .C1(new_n882), .C2(new_n867), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT108), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n876), .B2(new_n877), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n886), .B1(KEYINPUT54), .B2(new_n893), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n827), .A2(new_n894), .B1(G952), .B2(G953), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n585), .A2(new_n421), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(new_n355), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  OR4_X1    g713(.A1(new_n668), .A2(new_n674), .A3(new_n765), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n895), .A2(new_n900), .ZN(G75));
  NOR2_X1   g715(.A1(new_n562), .A2(new_n565), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n580), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  INV_X1    g718(.A(new_n889), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n836), .A2(new_n838), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n877), .B1(new_n906), .B2(new_n864), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT108), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n876), .A2(new_n891), .A3(new_n877), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n295), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n579), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n330), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n893), .A2(new_n451), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n567), .ZN(new_n918));
  NOR2_X1   g732(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n919));
  AND2_X1   g733(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n904), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n914), .A2(new_n922), .ZN(G51));
  NAND3_X1  g737(.A1(new_n893), .A2(new_n451), .A3(new_n754), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n412), .B(KEYINPUT57), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT54), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n908), .A2(new_n909), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n928), .B1(new_n929), .B2(new_n889), .ZN(new_n930));
  AOI211_X1 g744(.A(KEYINPUT54), .B(new_n905), .C1(new_n908), .C2(new_n909), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n406), .A2(new_n409), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n915), .B1(new_n926), .B2(new_n934), .ZN(G54));
  NAND4_X1  g749(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .A4(new_n513), .ZN(new_n936));
  INV_X1    g750(.A(new_n513), .ZN(new_n937));
  NAND2_X1  g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n917), .B2(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n936), .A2(new_n939), .A3(new_n916), .ZN(G60));
  NOR2_X1   g754(.A1(new_n930), .A2(new_n931), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n615), .B(KEYINPUT120), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT59), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n916), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n894), .B2(new_n944), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(G63));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT121), .Z(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT60), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n893), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n651), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n916), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n347), .B1(new_n893), .B2(new_n952), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT122), .ZN(new_n958));
  INV_X1    g772(.A(new_n952), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n910), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n960), .B2(new_n347), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n956), .A2(KEYINPUT122), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(KEYINPUT61), .B(new_n916), .C1(new_n953), .C2(new_n954), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n957), .B1(new_n963), .B2(new_n964), .ZN(G66));
  OAI21_X1  g779(.A(G953), .B1(new_n519), .B2(new_n539), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n879), .A2(new_n881), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(G953), .ZN(new_n968));
  INV_X1    g782(.A(new_n562), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(G898), .B2(new_n330), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n968), .B(new_n970), .ZN(G69));
  NOR2_X1   g785(.A1(new_n849), .A2(new_n759), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n748), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n769), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT123), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n681), .A2(new_n733), .A3(new_n829), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n778), .B1(new_n976), .B2(KEYINPUT62), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n975), .B(new_n977), .C1(KEYINPUT62), .C2(new_n976), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n330), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n267), .A2(new_n268), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n495), .A2(new_n496), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n330), .A2(G900), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n776), .A2(new_n777), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n758), .A2(new_n759), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n831), .A3(new_n739), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n985), .A2(new_n750), .A3(new_n769), .A4(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n746), .A2(new_n733), .A3(new_n829), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT125), .B1(new_n988), .B2(new_n991), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n984), .B1(new_n995), .B2(new_n330), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n983), .B1(new_n996), .B2(new_n982), .ZN(new_n997));
  OAI21_X1  g811(.A(G953), .B1(new_n402), .B2(new_n660), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT124), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n997), .B(new_n999), .ZN(G72));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT126), .ZN(new_n1003));
  INV_X1    g817(.A(new_n967), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1003), .B1(new_n978), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n915), .B1(new_n1005), .B2(new_n670), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n669), .A2(new_n259), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n993), .A2(new_n967), .A3(new_n994), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n1008), .A2(new_n1003), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n670), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(new_n1007), .A3(new_n1002), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT127), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1010), .B1(new_n885), .B2(new_n1013), .ZN(G57));
endmodule


