//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(KEYINPUT69), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT68), .B(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G137), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n461), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n460), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n466), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  OAI221_X1 g051(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT70), .Z(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT68), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n465), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n465), .A2(new_n479), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(G124), .A2(new_n485), .B1(new_n487), .B2(G136), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n478), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT71), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n471), .A2(new_n472), .A3(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(new_n483), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT4), .A2(G138), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n466), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n493), .B(new_n497), .C1(new_n498), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G651), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n507), .A2(new_n509), .B1(new_n506), .B2(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n507), .A2(new_n509), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n506), .A2(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(G543), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n513), .A2(G62), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT73), .Z(new_n524));
  OAI21_X1  g099(.A(G651), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n516), .A2(new_n521), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n515), .A2(G89), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n513), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT74), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n513), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G51), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n519), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n531), .B1(new_n539), .B2(KEYINPUT75), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n520), .A2(G51), .B1(new_n534), .B2(new_n536), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G168));
  XNOR2_X1  g119(.A(KEYINPUT76), .B(G52), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n510), .A2(G543), .A3(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI221_X1 g123(.A(new_n546), .B1(new_n547), .B2(new_n508), .C1(new_n514), .C2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(new_n515), .A2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n520), .A2(G43), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n508), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT78), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT77), .B(KEYINPUT8), .Z(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(new_n563), .ZN(G188));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n565));
  AND2_X1   g140(.A1(KEYINPUT5), .A2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(KEYINPUT5), .A2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(G65), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n565), .B1(new_n570), .B2(G651), .ZN(new_n571));
  AOI211_X1 g146(.A(KEYINPUT80), .B(new_n508), .C1(new_n568), .C2(new_n569), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(new_n514), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n519), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n510), .A2(new_n577), .A3(G53), .A4(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(KEYINPUT79), .A3(new_n578), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n574), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  XNOR2_X1  g159(.A(new_n549), .B(KEYINPUT81), .ZN(G301));
  NAND2_X1  g160(.A1(new_n539), .A2(KEYINPUT75), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n541), .A2(new_n542), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n586), .A2(new_n587), .A3(new_n531), .ZN(G286));
  NAND3_X1  g163(.A1(new_n510), .A2(G87), .A3(new_n513), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n510), .A2(G49), .A3(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  NAND3_X1  g167(.A1(new_n510), .A2(G86), .A3(new_n513), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n517), .A2(G48), .A3(G543), .A4(new_n518), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n511), .B2(new_n512), .ZN(new_n596));
  AND2_X1   g171(.A1(G73), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(new_n515), .A2(G85), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n520), .A2(G47), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n508), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(new_n513), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n520), .A2(G54), .B1(new_n608), .B2(G651), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n611));
  OR3_X1    g186(.A1(new_n514), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n514), .B2(new_n610), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n609), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n549), .B(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n615), .B1(new_n617), .B2(G868), .ZN(G321));
  XNOR2_X1  g193(.A(G321), .B(KEYINPUT83), .ZN(G284));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n583), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(G868), .B2(new_n583), .ZN(G280));
  INV_X1    g197(.A(new_n614), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g204(.A1(new_n479), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2100), .Z(new_n633));
  OAI221_X1 g208(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  INV_X1    g210(.A(G135), .ZN(new_n636));
  OAI221_X1 g211(.A(new_n634), .B1(new_n484), .B2(new_n635), .C1(new_n636), .C2(new_n486), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n633), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  XOR2_X1   g217(.A(KEYINPUT15), .B(G2435), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT85), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2427), .B(G2430), .Z(new_n646));
  OAI21_X1  g221(.A(KEYINPUT14), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT87), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n645), .A2(new_n646), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n649), .B2(new_n653), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n642), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n656), .ZN(new_n658));
  INV_X1    g233(.A(new_n642), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(new_n654), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G14), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n657), .B2(new_n660), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT88), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  OR3_X1    g262(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n691), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(KEYINPUT94), .ZN(new_n697));
  NAND2_X1  g272(.A1(G288), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n590), .A2(new_n589), .A3(KEYINPUT94), .A4(new_n591), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G23), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT95), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT33), .B(G1976), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n707), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n702), .A2(G22), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G166), .B2(new_n702), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1971), .ZN(new_n712));
  MUX2_X1   g287(.A(G6), .B(G305), .S(G16), .Z(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT32), .B(G1981), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n708), .A2(new_n709), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n708), .A2(new_n719), .A3(new_n709), .A4(new_n716), .ZN(new_n720));
  MUX2_X1   g295(.A(G24), .B(G290), .S(G16), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT93), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT92), .B(G1986), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G25), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT90), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n485), .A2(G119), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT91), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n466), .A2(G107), .ZN(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n487), .A2(G131), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  XOR2_X1   g311(.A(new_n735), .B(new_n736), .Z(new_n737));
  NAND4_X1  g312(.A1(new_n718), .A2(new_n720), .A3(new_n724), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT36), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n725), .A2(G35), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G162), .B2(new_n725), .ZN(new_n741));
  INV_X1    g316(.A(G2090), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT102), .B(KEYINPUT29), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n702), .A2(G19), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n556), .B2(new_n702), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G1341), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n702), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n623), .B2(new_n702), .ZN(new_n751));
  INV_X1    g326(.A(G1348), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n725), .A2(G26), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT28), .Z(new_n755));
  OAI221_X1 g330(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n756));
  INV_X1    g331(.A(G128), .ZN(new_n757));
  INV_X1    g332(.A(G140), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n756), .B1(new_n484), .B2(new_n757), .C1(new_n758), .C2(new_n486), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n755), .B1(new_n759), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2067), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n749), .A2(new_n753), .A3(new_n761), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n745), .A2(new_n746), .B1(KEYINPUT96), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n725), .A2(G33), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n765));
  NAND2_X1  g340(.A1(G103), .A2(G2104), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n483), .B2(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n487), .A2(G139), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n471), .A2(new_n472), .A3(G127), .ZN(new_n770));
  NAND2_X1  g345(.A1(G115), .A2(G2104), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n466), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT97), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n769), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n764), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT99), .ZN(new_n780));
  AND2_X1   g355(.A1(KEYINPUT24), .A2(G34), .ZN(new_n781));
  NOR2_X1   g356(.A1(KEYINPUT24), .A2(G34), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n725), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT98), .ZN(new_n784));
  INV_X1    g359(.A(G160), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n725), .ZN(new_n786));
  INV_X1    g361(.A(G2084), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n702), .A2(G5), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G171), .B2(new_n702), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(G1961), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n725), .A2(G32), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n487), .A2(G141), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n485), .A2(G129), .ZN(new_n794));
  NAND3_X1  g369(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT26), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n797), .A2(new_n798), .B1(G105), .B2(new_n468), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n793), .A2(new_n794), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n792), .B1(new_n801), .B2(new_n725), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT27), .B(G1996), .Z(new_n803));
  AOI211_X1 g378(.A(new_n788), .B(new_n791), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n780), .B1(new_n804), .B2(KEYINPUT101), .ZN(new_n805));
  NOR2_X1   g380(.A1(G164), .A2(new_n725), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G27), .B2(new_n725), .ZN(new_n807));
  INV_X1    g382(.A(G2078), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT31), .B(G11), .Z(new_n811));
  NOR2_X1   g386(.A1(new_n637), .A2(new_n725), .ZN(new_n812));
  INV_X1    g387(.A(G28), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT30), .ZN(new_n814));
  AOI21_X1  g389(.A(G29), .B1(new_n813), .B2(KEYINPUT30), .ZN(new_n815));
  AOI211_X1 g390(.A(new_n811), .B(new_n812), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n786), .A2(new_n787), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n809), .A2(new_n810), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n802), .A2(new_n803), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n819), .A2(KEYINPUT100), .B1(G1961), .B2(new_n790), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n777), .A2(new_n778), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n820), .B(new_n821), .C1(KEYINPUT100), .C2(new_n819), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n805), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n702), .A2(G21), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G168), .B2(new_n702), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G1966), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n825), .A2(G1966), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n804), .A2(KEYINPUT101), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n823), .A2(new_n826), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n702), .A2(G20), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT23), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n583), .B2(new_n702), .ZN(new_n833));
  INV_X1    g408(.A(G1956), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n763), .A2(new_n829), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n739), .A2(new_n837), .ZN(G311));
  NAND2_X1  g413(.A1(new_n739), .A2(new_n837), .ZN(G150));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n624), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n515), .A2(G93), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n520), .A2(G55), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(new_n508), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n842), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n555), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n841), .B(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n849), .A2(new_n850), .A3(G860), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(G860), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n851), .A2(new_n853), .ZN(G145));
  INV_X1    g429(.A(KEYINPUT105), .ZN(new_n855));
  INV_X1    g430(.A(new_n734), .ZN(new_n856));
  OAI221_X1 g431(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n857));
  INV_X1    g432(.A(G130), .ZN(new_n858));
  INV_X1    g433(.A(G142), .ZN(new_n859));
  OAI221_X1 g434(.A(new_n857), .B1(new_n484), .B2(new_n858), .C1(new_n859), .C2(new_n486), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT104), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n631), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n860), .A2(KEYINPUT104), .ZN(new_n863));
  INV_X1    g438(.A(new_n631), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(KEYINPUT104), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n856), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n862), .A2(new_n866), .A3(new_n856), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n855), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n871), .A2(KEYINPUT105), .A3(new_n867), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n776), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n759), .A2(new_n503), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n759), .A2(new_n503), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n875), .A2(new_n800), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n800), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n776), .B(KEYINPUT103), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR3_X1    g457(.A1(new_n870), .A2(new_n872), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n785), .B(new_n637), .ZN(new_n884));
  XNOR2_X1  g459(.A(G162), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n871), .A2(new_n867), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(new_n882), .A3(new_n855), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n870), .A2(new_n872), .A3(new_n882), .ZN(new_n891));
  INV_X1    g466(.A(new_n888), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n885), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g470(.A(G303), .B(G290), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n700), .B(G305), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n847), .B(new_n626), .Z(new_n901));
  NAND2_X1  g476(.A1(G299), .A2(new_n614), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n583), .A2(new_n623), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n902), .A2(KEYINPUT41), .A3(new_n903), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT41), .B1(new_n902), .B2(new_n903), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n905), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n900), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n912), .A2(new_n900), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G868), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n846), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(G295));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n917), .ZN(G331));
  OAI21_X1  g494(.A(new_n549), .B1(new_n540), .B2(new_n543), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(G301), .B2(G286), .ZN(new_n921));
  INV_X1    g496(.A(new_n847), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n847), .B(new_n920), .C1(G286), .C2(G301), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT108), .B1(new_n925), .B2(new_n904), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n923), .B(new_n924), .C1(new_n906), .C2(new_n907), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n898), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n890), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n898), .B1(new_n926), .B2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT110), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n927), .ZN(new_n932));
  INV_X1    g507(.A(new_n898), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n890), .A4(new_n928), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(KEYINPUT43), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n931), .A2(new_n936), .A3(KEYINPUT111), .A4(KEYINPUT43), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n929), .A2(new_n930), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n940), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n934), .A2(new_n943), .A3(new_n890), .A4(new_n928), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n928), .A2(new_n890), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n949), .A2(KEYINPUT109), .A3(new_n943), .A4(new_n934), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n948), .B(new_n950), .C1(new_n943), .C2(new_n942), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n941), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n945), .A2(new_n952), .ZN(G397));
  INV_X1    g528(.A(new_n475), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n954), .A2(G40), .A3(new_n469), .A4(new_n467), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(G2084), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n497), .B1(new_n502), .B2(new_n498), .ZN(new_n959));
  INV_X1    g534(.A(new_n493), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n957), .B(new_n958), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT113), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n957), .B1(new_n503), .B2(new_n958), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n480), .A2(new_n482), .A3(new_n501), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n499), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n496), .B1(new_n966), .B2(new_n465), .ZN(new_n967));
  AOI21_X1  g542(.A(G1384), .B1(new_n967), .B2(new_n493), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n968), .A2(KEYINPUT113), .A3(new_n957), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT117), .B(new_n956), .C1(new_n964), .C2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n972), .B(G1384), .C1(new_n967), .C2(new_n493), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT45), .B1(new_n503), .B2(new_n958), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n973), .A2(new_n974), .A3(new_n955), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n971), .B1(new_n975), .B2(G1966), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n503), .A2(new_n958), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n972), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n470), .A2(new_n979), .A3(new_n475), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n958), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1966), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(KEYINPUT116), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n970), .A2(new_n976), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n977), .A2(KEYINPUT50), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(KEYINPUT113), .A3(new_n961), .ZN(new_n987));
  OR3_X1    g562(.A1(new_n968), .A2(KEYINPUT113), .A3(new_n957), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT117), .B1(new_n989), .B2(new_n956), .ZN(new_n990));
  OAI21_X1  g565(.A(G286), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n982), .A2(KEYINPUT116), .A3(new_n983), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT116), .B1(new_n982), .B2(new_n983), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n956), .B1(new_n964), .B2(new_n969), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n994), .A2(G168), .A3(new_n997), .A4(new_n970), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n991), .A2(new_n998), .A3(G8), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT51), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n1001), .A3(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT62), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1000), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n975), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n955), .B1(new_n987), .B2(new_n988), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT122), .B(G1961), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1007), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT123), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT123), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(new_n1007), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n982), .B2(G2078), .ZN(new_n1017));
  AOI21_X1  g592(.A(G301), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n742), .B(new_n980), .C1(new_n964), .C2(new_n969), .ZN(new_n1019));
  INV_X1    g594(.A(G1971), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n982), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G8), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G303), .A2(G8), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT114), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n1026), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n593), .A2(new_n598), .A3(new_n1035), .A4(new_n594), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT49), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1029), .B1(new_n980), .B2(new_n968), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT115), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1039), .A2(new_n1044), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n698), .A2(G1976), .A3(new_n699), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1040), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1048), .A2(new_n1040), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1049), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n986), .A2(new_n980), .A3(new_n961), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1021), .B1(G2090), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1026), .B1(new_n1056), .B2(G8), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1018), .A2(new_n1033), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1004), .A2(new_n1006), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n980), .B1(new_n968), .B2(new_n957), .ZN(new_n1061));
  INV_X1    g636(.A(new_n961), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n834), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1055), .A2(KEYINPUT119), .A3(new_n834), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n574), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n579), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n583), .B2(new_n1069), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n982), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1067), .A2(new_n1072), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n980), .A2(new_n968), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G2067), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1008), .B2(G1348), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(new_n614), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1072), .B1(new_n1067), .B2(new_n1076), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1077), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1075), .B(new_n1071), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n1085), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT119), .B1(new_n1055), .B2(new_n834), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1076), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1071), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(KEYINPUT61), .A3(new_n1077), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1082), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(KEYINPUT60), .B(new_n1081), .C1(new_n1008), .C2(G1348), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n623), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1089), .A2(new_n1094), .A3(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT120), .B(G1996), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n975), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n975), .A2(KEYINPUT121), .A3(new_n1100), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n1078), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n556), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1097), .A2(new_n623), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(KEYINPUT59), .A3(new_n556), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1086), .B1(new_n1099), .B2(new_n1113), .ZN(new_n1114));
  AND4_X1   g689(.A1(new_n1031), .A2(new_n1022), .A3(G8), .A4(new_n1026), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1031), .B1(new_n1030), .B2(new_n1026), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1058), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n980), .B1(new_n964), .B2(new_n969), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1009), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n470), .A2(KEYINPUT124), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT125), .B(G2078), .Z(new_n1123));
  NAND4_X1  g698(.A1(new_n954), .A2(KEYINPUT53), .A3(G40), .A4(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n470), .A2(KEYINPUT124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(new_n978), .A3(new_n981), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1121), .A2(new_n1017), .A3(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(new_n617), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1119), .B1(new_n1018), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1013), .B1(new_n1121), .B2(new_n1007), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1014), .ZN(new_n1132));
  OAI211_X1 g707(.A(G301), .B(new_n1017), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1015), .A2(KEYINPUT126), .A3(G301), .A4(new_n1017), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1119), .B1(new_n1128), .B2(G171), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1114), .A2(new_n1118), .A3(new_n1130), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n994), .A2(new_n997), .A3(new_n970), .ZN(new_n1142));
  NOR2_X1   g717(.A1(G286), .A2(new_n1029), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1030), .A2(new_n1026), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT63), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g721(.A(G1976), .B(G288), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1036), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1040), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1057), .A2(KEYINPUT63), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1054), .B1(new_n1033), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1140), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1033), .A2(new_n1152), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1141), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1156), .A2(KEYINPUT118), .A3(new_n1149), .A4(new_n1146), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1060), .A2(new_n1139), .A3(new_n1154), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n856), .A2(new_n736), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n800), .B(G1996), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n759), .B(G2067), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n856), .A2(new_n736), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1160), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(G290), .A2(G1986), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT112), .ZN(new_n1167));
  NAND2_X1  g742(.A1(G290), .A2(G1986), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n978), .A2(new_n955), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1158), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1170), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1173), .A2(G1996), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT46), .Z(new_n1175));
  OAI21_X1  g750(.A(new_n1170), .B1(new_n1162), .B2(new_n800), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT47), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1165), .A2(new_n1173), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1167), .A2(new_n1173), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1179), .B1(KEYINPUT48), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(KEYINPUT48), .B2(new_n1180), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1163), .A2(new_n1159), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n759), .A2(G2067), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1170), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1178), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1172), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g762(.A(G319), .ZN(new_n1189));
  NOR2_X1   g763(.A1(G227), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g764(.A(new_n1190), .B1(new_n663), .B2(new_n664), .ZN(new_n1191));
  AOI21_X1  g765(.A(G229), .B1(new_n1191), .B2(KEYINPUT127), .ZN(new_n1192));
  OR2_X1    g766(.A1(new_n1191), .A2(KEYINPUT127), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n894), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1194), .A2(new_n951), .ZN(G225));
  INV_X1    g769(.A(G225), .ZN(G308));
endmodule


