//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G68), .A2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G58), .C2(G232), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G1), .B2(G20), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n206), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n210), .B(new_n222), .C1(new_n224), .C2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  INV_X1    g0031(.A(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n213), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  INV_X1    g0039(.A(G107), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n212), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n223), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G68), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n250), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G68), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT74), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT74), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n206), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n254), .B1(new_n263), .B2(KEYINPUT7), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT7), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n262), .A2(new_n265), .A3(new_n206), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n253), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n249), .B1(new_n267), .B2(KEYINPUT16), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT3), .B1(new_n256), .B2(new_n258), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(KEYINPUT7), .B(new_n206), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n261), .A2(new_n270), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n265), .B1(new_n273), .B2(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n253), .B1(new_n275), .B2(G68), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(KEYINPUT16), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n268), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(new_n223), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n232), .A2(G1698), .ZN(new_n283));
  OR2_X1    g0083(.A1(G223), .A2(G1698), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n259), .A2(new_n261), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G87), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT66), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(new_n280), .B2(new_n223), .ZN(new_n291));
  AND2_X1   g0091(.A1(G1), .A2(G13), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(KEYINPUT66), .A3(new_n293), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n229), .B(new_n289), .C1(new_n291), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  AOI211_X1 g0096(.A(new_n296), .B(new_n288), .C1(new_n291), .C2(new_n294), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n287), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G13), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n303), .A2(new_n206), .A3(G1), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n248), .B1(new_n205), .B2(G20), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n302), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n298), .A2(G190), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n279), .A2(new_n300), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT17), .ZN(new_n311));
  INV_X1    g0111(.A(new_n261), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT74), .B(G33), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(KEYINPUT3), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT7), .B1(new_n314), .B2(G20), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(G68), .A3(new_n266), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(KEYINPUT16), .A3(new_n252), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n248), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n308), .B1(new_n318), .B2(new_n277), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT17), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n300), .A4(new_n309), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n311), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n302), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n206), .A2(G33), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT15), .B(G87), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n248), .B1(new_n202), .B2(new_n304), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT69), .B1(new_n307), .B2(G77), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n307), .A2(KEYINPUT69), .A3(G77), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n296), .B1(new_n291), .B2(new_n294), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n289), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n289), .B1(new_n291), .B2(new_n294), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G244), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n333), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT68), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n273), .A2(G238), .A3(G1698), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n240), .B2(new_n273), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n261), .A2(new_n270), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n341), .A2(new_n229), .A3(G1698), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n281), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT68), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n333), .B(new_n344), .C1(new_n335), .C2(new_n336), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n338), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n331), .B1(new_n346), .B2(G200), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n338), .A2(new_n343), .A3(G190), .A4(new_n345), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n251), .A2(G150), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n350), .B1(new_n201), .B2(new_n206), .C1(new_n301), .C2(new_n325), .ZN(new_n351));
  INV_X1    g0151(.A(G50), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n351), .A2(new_n248), .B1(new_n352), .B2(new_n304), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n307), .A2(G50), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT9), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n353), .A2(KEYINPUT9), .A3(new_n354), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n261), .A2(new_n270), .A3(G223), .A4(G1698), .ZN(new_n359));
  INV_X1    g0159(.A(G1698), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n261), .A2(new_n270), .A3(G222), .A4(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n361), .C1(new_n273), .C2(new_n202), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n281), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n334), .A2(G226), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n333), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G200), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n363), .A2(G190), .A3(new_n333), .A4(new_n364), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n357), .A2(new_n358), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT10), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n355), .A2(new_n356), .B1(new_n365), .B2(G200), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT10), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n358), .A4(new_n367), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT67), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT67), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G179), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n355), .B1(new_n365), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G169), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n365), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n349), .A2(new_n373), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT75), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n298), .A2(G169), .ZN(new_n386));
  NOR4_X1   g0186(.A1(new_n287), .A2(new_n295), .A3(new_n297), .A4(new_n379), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n298), .A2(new_n378), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n389), .B(KEYINPUT75), .C1(G169), .C2(new_n298), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n319), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT18), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n319), .A2(new_n388), .A3(new_n390), .A4(KEYINPUT18), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n323), .A2(new_n384), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n261), .A2(new_n270), .A3(G226), .A4(new_n360), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n261), .A2(new_n270), .A3(G232), .A4(G1698), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n255), .A2(new_n217), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT70), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT70), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n397), .A2(new_n398), .A3(new_n403), .A4(new_n400), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n281), .A3(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(G238), .A2(new_n334), .B1(new_n332), .B2(new_n289), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT13), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT71), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT13), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n410), .A3(new_n406), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n407), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(G200), .A3(new_n413), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n325), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT72), .ZN(new_n416));
  INV_X1    g0216(.A(new_n251), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n352), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n248), .ZN(new_n419));
  XOR2_X1   g0219(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n418), .A2(new_n248), .A3(new_n420), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n304), .A2(new_n254), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT12), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n307), .A2(G68), .B1(new_n424), .B2(new_n425), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n422), .A2(new_n423), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n408), .A2(G190), .A3(new_n411), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n414), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n412), .A2(G169), .A3(new_n413), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n408), .A2(G179), .A3(new_n411), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n412), .A2(new_n437), .A3(G169), .A4(new_n413), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n433), .B1(new_n439), .B2(new_n429), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n346), .A2(new_n381), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n331), .C1(new_n346), .C2(new_n379), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n396), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n305), .B(new_n249), .C1(G1), .C2(new_n255), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G107), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n304), .B(new_n240), .C1(KEYINPUT86), .C2(KEYINPUT25), .ZN(new_n448));
  NAND2_X1  g0248(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n206), .A2(G107), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT84), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(KEYINPUT23), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT22), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n261), .A2(new_n270), .A3(new_n206), .A4(G87), .ZN(new_n457));
  XOR2_X1   g0257(.A(KEYINPUT84), .B(KEYINPUT23), .Z(new_n458));
  AOI22_X1  g0258(.A1(new_n456), .A2(new_n457), .B1(new_n458), .B2(new_n451), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n313), .A2(new_n212), .ZN(new_n460));
  INV_X1    g0260(.A(G87), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n314), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n455), .B(new_n459), .C1(new_n463), .C2(G20), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT24), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n259), .A2(new_n261), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n256), .A2(new_n258), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G116), .ZN(new_n468));
  AOI21_X1  g0268(.A(G20), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT24), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n455), .A4(new_n459), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT85), .B1(new_n473), .B2(new_n248), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT85), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n475), .B(new_n249), .C1(new_n465), .C2(new_n472), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n447), .B(new_n450), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n218), .A2(G1698), .ZN(new_n478));
  OR2_X1    g0278(.A1(G250), .A2(G1698), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n259), .A2(new_n261), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G294), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n313), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n281), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT5), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G41), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n205), .A2(G45), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT79), .B1(new_n484), .B2(G41), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT79), .ZN(new_n488));
  INV_X1    g0288(.A(G41), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT5), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n486), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n332), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n485), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n291), .A2(new_n294), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(G264), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n483), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n381), .ZN(new_n497));
  INV_X1    g0297(.A(new_n496), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n374), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n477), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n336), .A2(G1698), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n259), .A2(new_n261), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT77), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT4), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT77), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n259), .A2(new_n505), .A3(new_n261), .A4(new_n501), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n273), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n273), .A2(G250), .A3(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n281), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT78), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n493), .A2(G257), .A3(new_n494), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n492), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n282), .B1(new_n507), .B2(new_n511), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT78), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n515), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n513), .A2(G190), .A3(new_n518), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT80), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n517), .B1(new_n512), .B2(new_n281), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(KEYINPUT80), .A3(G190), .ZN(new_n526));
  AOI22_X1  g0326(.A1(G200), .A2(new_n521), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n305), .A2(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n445), .A2(new_n217), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n217), .A2(new_n240), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n240), .A2(KEYINPUT6), .A3(G97), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n206), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n417), .A2(new_n202), .ZN(new_n536));
  AOI211_X1 g0336(.A(new_n535), .B(new_n536), .C1(new_n275), .C2(G107), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT76), .B1(new_n537), .B2(new_n249), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n275), .B2(G107), .ZN(new_n539));
  INV_X1    g0339(.A(new_n535), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT76), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(new_n248), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n528), .B(new_n529), .C1(new_n538), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n527), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n528), .B1(new_n538), .B2(new_n543), .ZN(new_n546));
  INV_X1    g0346(.A(new_n529), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n381), .B1(new_n519), .B2(new_n517), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n519), .A2(KEYINPUT78), .ZN(new_n550));
  AOI211_X1 g0350(.A(new_n514), .B(new_n282), .C1(new_n507), .C2(new_n511), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n550), .A2(new_n551), .A3(new_n517), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n378), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n500), .A2(new_n545), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n457), .A2(new_n456), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n458), .A2(new_n451), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n469), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n471), .B1(new_n559), .B2(new_n455), .ZN(new_n560));
  NOR4_X1   g0360(.A1(new_n469), .A2(new_n558), .A3(KEYINPUT24), .A4(new_n454), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n248), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n475), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n473), .A2(KEYINPUT85), .A3(new_n248), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n563), .A2(new_n564), .B1(G107), .B2(new_n446), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n496), .A2(G200), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n498), .A2(G190), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n565), .A2(new_n450), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n510), .B(new_n206), .C1(G33), .C2(new_n217), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n569), .B(new_n248), .C1(new_n206), .C2(G116), .ZN(new_n570));
  XOR2_X1   g0370(.A(new_n570), .B(KEYINPUT20), .Z(new_n571));
  NAND2_X1  g0371(.A1(new_n446), .A2(G116), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(G116), .C2(new_n305), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OR2_X1    g0374(.A1(new_n360), .A2(G264), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n218), .A2(new_n360), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n259), .A2(new_n261), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n341), .A2(G303), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n281), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n493), .A2(G270), .A3(new_n494), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n580), .A2(new_n492), .A3(G179), .A4(new_n581), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n574), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n492), .A3(new_n581), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G200), .ZN(new_n585));
  INV_X1    g0385(.A(G190), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n574), .B(new_n585), .C1(new_n586), .C2(new_n584), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n573), .A2(G169), .A3(new_n584), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n573), .A2(KEYINPUT21), .A3(G169), .A4(new_n584), .ZN(new_n591));
  AND4_X1   g0391(.A1(new_n583), .A2(new_n587), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n494), .A2(G250), .A3(new_n486), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n494), .A2(KEYINPUT81), .A3(G250), .A4(new_n486), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n290), .A2(new_n205), .A3(G45), .A4(G274), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n336), .A2(G1698), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(G238), .B2(G1698), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n468), .B1(new_n262), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n281), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n597), .A2(G190), .A3(new_n598), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT83), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n597), .A2(new_n598), .A3(new_n602), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G200), .ZN(new_n606));
  INV_X1    g0406(.A(new_n326), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n305), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n445), .A2(new_n461), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n314), .A2(new_n206), .A3(G68), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n325), .A2(new_n217), .ZN(new_n611));
  XNOR2_X1  g0411(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(G20), .B1(new_n612), .B2(new_n399), .ZN(new_n614));
  NOR3_X1   g0414(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n610), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n608), .B(new_n609), .C1(new_n616), .C2(new_n248), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n595), .A2(new_n596), .B1(new_n281), .B2(new_n601), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT83), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(G190), .A4(new_n598), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n604), .A2(new_n606), .A3(new_n617), .A4(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n608), .B1(new_n616), .B2(new_n248), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n326), .B2(new_n445), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n605), .A2(new_n381), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n618), .A2(new_n378), .A3(new_n598), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n568), .A2(new_n592), .A3(new_n627), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n444), .A2(new_n555), .A3(new_n628), .ZN(G372));
  NAND2_X1  g0429(.A1(new_n323), .A2(new_n432), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n439), .A2(new_n429), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n631), .B2(new_n442), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n386), .A2(new_n387), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n319), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(new_n392), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n373), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(new_n383), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n624), .A2(KEYINPUT87), .A3(new_n625), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT87), .B1(new_n624), .B2(new_n625), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n623), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n606), .A2(KEYINPUT88), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n606), .A2(KEYINPUT88), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n642), .A2(new_n617), .A3(new_n603), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n546), .A2(new_n547), .B1(new_n552), .B2(new_n378), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n549), .A4(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n549), .A3(new_n627), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n641), .A2(KEYINPUT89), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT89), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n652), .B(new_n623), .C1(new_n639), .C2(new_n640), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n650), .A2(KEYINPUT26), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n583), .A2(new_n590), .A3(new_n591), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n500), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n549), .A2(new_n648), .B1(new_n527), .B2(new_n544), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n646), .A2(new_n568), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n649), .B(new_n654), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n638), .B1(new_n444), .B2(new_n662), .ZN(G369));
  NOR2_X1   g0463(.A1(new_n303), .A2(G20), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n205), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n573), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n592), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n656), .B2(new_n671), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(G330), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n477), .A2(new_n670), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n568), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n500), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n500), .A2(new_n670), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n670), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n655), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(new_n679), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n207), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n615), .A2(new_n212), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n225), .B2(new_n690), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n661), .A2(new_n683), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(KEYINPUT29), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT26), .B1(new_n645), .B2(new_n554), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n651), .A2(new_n653), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n648), .A2(new_n627), .A3(new_n647), .A4(new_n549), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n657), .A2(new_n658), .A3(new_n568), .A4(new_n646), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n670), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT29), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n698), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n568), .A2(new_n592), .A3(new_n627), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n658), .A3(new_n500), .A4(new_n683), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n483), .A2(new_n495), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n582), .A2(new_n712), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n597), .A2(new_n598), .A3(new_n602), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n714), .A3(new_n525), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n605), .A2(new_n378), .A3(new_n584), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n521), .A2(new_n496), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n715), .A2(new_n716), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT91), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(KEYINPUT90), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT90), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n715), .A2(new_n725), .A3(new_n716), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n724), .A2(new_n717), .A3(new_n719), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n670), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n723), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI211_X1 g0530(.A(KEYINPUT91), .B(KEYINPUT31), .C1(new_n727), .C2(new_n670), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n711), .B(new_n722), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n709), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n695), .B1(new_n735), .B2(G1), .ZN(G364));
  AOI21_X1  g0536(.A(new_n205), .B1(new_n664), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n689), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n674), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G330), .B2(new_n673), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n292), .B1(new_n206), .B2(G169), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT93), .Z(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n206), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT92), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT94), .Z(new_n748));
  NOR2_X1   g0548(.A1(new_n225), .A2(G45), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n245), .B2(G45), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n314), .A2(new_n688), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n750), .A2(new_n751), .B1(new_n212), .B2(new_n688), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n273), .A2(G355), .A3(new_n207), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n206), .A2(G190), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(new_n374), .A3(G200), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT97), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n760), .A2(KEYINPUT98), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(KEYINPUT98), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G107), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n374), .A2(G20), .A3(G190), .A4(G200), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT96), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT96), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G87), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n765), .A2(new_n273), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT99), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n379), .A2(new_n299), .A3(new_n755), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n378), .A2(new_n206), .A3(new_n586), .A4(G200), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n775), .A2(G77), .B1(G58), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n379), .A2(G20), .A3(G200), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(new_n586), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n777), .B1(new_n352), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G179), .A2(G200), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n206), .B1(new_n781), .B2(G190), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n217), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n755), .A2(new_n781), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT95), .B(KEYINPUT32), .Z(new_n787));
  XNOR2_X1  g0587(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n780), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n778), .A2(G190), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n773), .B(new_n789), .C1(new_n254), .C2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G326), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n341), .B1(new_n481), .B2(new_n782), .C1(new_n779), .C2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n784), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(G329), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n764), .A2(G283), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n776), .A2(G322), .ZN(new_n798));
  INV_X1    g0598(.A(G303), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n769), .A2(new_n799), .B1(new_n774), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(new_n790), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n792), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n743), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n754), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n807), .B(new_n739), .C1(new_n673), .C2(new_n746), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n741), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  NAND2_X1  g0610(.A1(new_n331), .A2(new_n670), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n349), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n442), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n442), .A2(new_n670), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n696), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(new_n733), .ZN(new_n818));
  INV_X1    g0618(.A(new_n739), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n763), .A2(new_n254), .ZN(new_n821));
  INV_X1    g0621(.A(G58), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n314), .B1(new_n822), .B2(new_n782), .C1(new_n769), .C2(new_n352), .ZN(new_n823));
  INV_X1    g0623(.A(new_n779), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(G137), .B1(G150), .B2(new_n790), .ZN(new_n825));
  INV_X1    g0625(.A(G143), .ZN(new_n826));
  INV_X1    g0626(.A(new_n776), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n827), .C1(new_n785), .C2(new_n774), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT34), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n821), .B(new_n823), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n829), .B2(new_n828), .C1(new_n831), .C2(new_n784), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n774), .A2(new_n212), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n341), .B1(new_n784), .B2(new_n800), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n783), .B(new_n834), .C1(new_n824), .C2(G303), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n827), .A2(new_n481), .B1(new_n240), .B2(new_n769), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G283), .B2(new_n790), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n835), .B(new_n837), .C1(new_n461), .C2(new_n763), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n832), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n744), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n743), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT100), .Z(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n839), .A2(new_n806), .B1(new_n202), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n844), .B(new_n739), .C1(new_n816), .C2(new_n840), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n820), .A2(new_n845), .ZN(G384));
  INV_X1    g0646(.A(new_n668), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n319), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n310), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n391), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n267), .A2(KEYINPUT16), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n308), .B1(new_n852), .B2(new_n318), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n847), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n633), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n310), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n323), .A2(new_n395), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n859), .B2(new_n854), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n858), .B(KEYINPUT38), .C1(new_n859), .C2(new_n854), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT40), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT31), .B1(new_n727), .B2(new_n670), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n711), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n429), .A2(new_n670), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT104), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n871), .B(new_n872), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n631), .A2(new_n432), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n631), .B2(new_n432), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n874), .A2(new_n875), .A3(new_n815), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n864), .A2(new_n865), .A3(new_n870), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n848), .B1(new_n635), .B2(new_n323), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n310), .A2(new_n634), .A3(new_n848), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n850), .A2(new_n391), .B1(new_n879), .B2(KEYINPUT37), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n861), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n863), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n882), .A2(new_n870), .A3(new_n876), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n877), .B1(new_n883), .B2(new_n865), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n870), .A2(new_n443), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(G330), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n874), .A2(new_n875), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n661), .A2(new_n683), .A3(new_n816), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT103), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n889), .A2(new_n890), .A3(new_n814), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n889), .B2(new_n814), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n888), .B(new_n864), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n636), .A2(new_n668), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n882), .A2(KEYINPUT39), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n631), .A2(new_n670), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n893), .A2(new_n894), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n887), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n443), .B1(new_n697), .B2(new_n706), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n638), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n901), .B(new_n903), .Z(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n205), .B2(new_n664), .ZN(new_n905));
  OAI21_X1  g0705(.A(G77), .B1(new_n822), .B2(new_n254), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n906), .A2(new_n225), .B1(G50), .B2(new_n254), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(G1), .A3(new_n303), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n533), .A2(new_n534), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT101), .Z(new_n910));
  AOI21_X1  g0710(.A(new_n212), .B1(new_n910), .B2(KEYINPUT35), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(new_n224), .C1(KEYINPUT35), .C2(new_n910), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT102), .B(KEYINPUT36), .Z(new_n913));
  XNOR2_X1  g0713(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n905), .A2(new_n908), .A3(new_n914), .ZN(G367));
  INV_X1    g0715(.A(KEYINPUT44), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n658), .B1(new_n544), .B2(new_n683), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n648), .A2(new_n549), .A3(new_n670), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n916), .B1(new_n686), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n685), .A2(new_n679), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n921), .A2(KEYINPUT44), .A3(new_n917), .A4(new_n918), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n685), .A2(new_n679), .A3(new_n919), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT45), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(KEYINPUT108), .A3(new_n682), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n682), .A2(KEYINPUT108), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n682), .A2(KEYINPUT108), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n923), .A2(new_n926), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n680), .B(new_n684), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(new_n674), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n734), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n936));
  XOR2_X1   g0736(.A(new_n689), .B(new_n936), .Z(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n737), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n680), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n940), .A2(new_n655), .A3(new_n683), .A4(new_n919), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n554), .B1(new_n917), .B2(new_n500), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n683), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n617), .A2(new_n683), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n651), .A2(new_n653), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n645), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n952), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n946), .A2(new_n954), .A3(new_n950), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(KEYINPUT105), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT106), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n681), .A2(new_n919), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n953), .A2(new_n955), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n959), .A2(new_n960), .B1(KEYINPUT105), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n956), .A2(new_n958), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT106), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n961), .A2(KEYINPUT105), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n939), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n236), .A2(new_n688), .A3(new_n314), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n969), .B(new_n748), .C1(new_n688), .C2(new_n607), .ZN(new_n970));
  INV_X1    g0770(.A(G283), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n760), .A2(new_n217), .B1(new_n971), .B2(new_n774), .ZN(new_n972));
  INV_X1    g0772(.A(new_n782), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n314), .B(new_n972), .C1(G107), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n795), .A2(G317), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n791), .A2(new_n481), .B1(new_n799), .B2(new_n827), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G311), .B2(new_n824), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n770), .A2(G116), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT46), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n974), .A2(new_n975), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n779), .A2(new_n826), .B1(new_n254), .B2(new_n782), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n341), .B(new_n981), .C1(G137), .C2(new_n795), .ZN(new_n982));
  INV_X1    g0782(.A(G150), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n827), .A2(new_n983), .B1(new_n352), .B2(new_n774), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n790), .B2(G159), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n982), .B(new_n985), .C1(new_n822), .C2(new_n769), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n760), .A2(new_n202), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n980), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n970), .B1(new_n989), .B2(new_n806), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n990), .B(new_n739), .C1(new_n746), .C2(new_n949), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n968), .A2(new_n991), .ZN(G387));
  NAND2_X1  g0792(.A1(new_n302), .A2(new_n352), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n692), .B1(new_n254), .B2(new_n202), .C1(new_n993), .C2(KEYINPUT50), .ZN(new_n994));
  AOI211_X1 g0794(.A(G45), .B(new_n994), .C1(KEYINPUT50), .C2(new_n993), .ZN(new_n995));
  INV_X1    g0795(.A(G45), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n751), .B1(new_n233), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n273), .A2(new_n691), .A3(new_n207), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n240), .B2(new_n688), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n739), .B1(new_n1000), .B2(new_n748), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT109), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n784), .A2(new_n793), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n760), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n314), .B1(new_n1005), .B2(G116), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n790), .A2(G311), .B1(G317), .B2(new_n776), .ZN(new_n1007));
  XOR2_X1   g0807(.A(KEYINPUT110), .B(G322), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1007), .B1(new_n799), .B2(new_n774), .C1(new_n779), .C2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT48), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n971), .B2(new_n782), .C1(new_n481), .C2(new_n769), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(KEYINPUT111), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(KEYINPUT111), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT49), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1012), .A2(KEYINPUT111), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT49), .B1(new_n1018), .B2(new_n1013), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1004), .B(new_n1006), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n769), .A2(new_n202), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n779), .A2(new_n785), .B1(new_n254), .B2(new_n774), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n314), .B1(new_n983), .B2(new_n784), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n782), .A2(new_n326), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n790), .A2(new_n302), .B1(G50), .B2(new_n776), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1021), .B(new_n1027), .C1(G97), .C2(new_n764), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1020), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1002), .B1(new_n1030), .B2(new_n806), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(KEYINPUT112), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT112), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1033), .B(new_n1002), .C1(new_n1030), .C2(new_n806), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n1032), .A2(new_n1034), .B1(new_n940), .B2(new_n746), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT113), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT113), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n940), .B2(new_n746), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1036), .A2(new_n1038), .B1(new_n738), .B2(new_n934), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n735), .A2(new_n934), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n735), .A2(new_n934), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n689), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1039), .A2(new_n1042), .ZN(G393));
  INV_X1    g0843(.A(KEYINPUT115), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n919), .A2(new_n746), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n207), .A2(new_n217), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1046), .B(new_n748), .C1(new_n242), .C2(new_n751), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n779), .A2(new_n983), .B1(new_n785), .B2(new_n827), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n769), .A2(new_n254), .B1(new_n774), .B2(new_n301), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n973), .A2(G77), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n314), .C1(new_n826), .C2(new_n784), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1049), .B(new_n1053), .C1(new_n461), .C2(new_n763), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n791), .A2(new_n352), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n795), .A2(new_n1008), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G283), .A2(new_n770), .B1(new_n775), .B2(G294), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n341), .B1(new_n782), .B2(new_n212), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n790), .B2(G303), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n765), .A2(new_n1056), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n824), .A2(G317), .B1(G311), .B2(new_n776), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1054), .A2(new_n1055), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1047), .B1(new_n1064), .B2(new_n806), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1045), .A2(new_n739), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n932), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1044), .B(new_n1066), .C1(new_n1067), .C2(new_n737), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n737), .B1(new_n928), .B2(new_n931), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1066), .ZN(new_n1070));
  OAI21_X1  g0870(.A(KEYINPUT115), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n690), .B1(new_n1067), .B2(new_n1041), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n932), .A2(new_n735), .A3(new_n934), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1068), .A2(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G390));
  NAND3_X1  g0875(.A1(new_n870), .A2(new_n876), .A3(G330), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT116), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n870), .A2(new_n876), .A3(KEYINPUT116), .A4(G330), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n898), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n897), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n814), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n704), .B2(new_n813), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n888), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n882), .A2(new_n1083), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1081), .B1(new_n1084), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n897), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n889), .A2(new_n814), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT103), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n889), .A2(new_n890), .A3(new_n814), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1087), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1092), .B1(new_n1096), .B2(new_n898), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n722), .B1(new_n730), .B2(new_n731), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n628), .A2(new_n555), .A3(new_n670), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n876), .B(G330), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT117), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT117), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n732), .A2(new_n1102), .A3(G330), .A4(new_n876), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1090), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1097), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1091), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n738), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT121), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n1111), .A3(new_n738), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n728), .A2(new_n729), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n866), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n443), .B(G330), .C1(new_n1099), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT118), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT118), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n870), .A2(new_n1118), .A3(G330), .A4(new_n443), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n902), .A2(new_n638), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(G330), .B1(new_n1099), .B2(new_n1115), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n816), .B1(new_n1122), .B2(KEYINPUT119), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT119), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n870), .B2(G330), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1087), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1104), .A2(new_n1126), .A3(new_n1086), .ZN(new_n1127));
  OAI211_X1 g0927(.A(G330), .B(new_n816), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1087), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(KEYINPUT120), .B(new_n1121), .C1(new_n1127), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT120), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1121), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1108), .B1(new_n1133), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1122), .A2(KEYINPUT119), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n870), .A2(new_n1124), .A3(G330), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n1140), .A3(new_n816), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1087), .A2(new_n1141), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1142), .A2(new_n1086), .B1(new_n1131), .B2(new_n1130), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT120), .B1(new_n1143), .B2(new_n1121), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1135), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1144), .A2(new_n1145), .A3(new_n1107), .A4(new_n1091), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1138), .A2(new_n1146), .A3(new_n689), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n273), .B1(new_n795), .B2(G294), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n771), .A2(new_n1051), .A3(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n779), .A2(new_n971), .B1(new_n212), .B2(new_n827), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(G97), .C2(new_n775), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n254), .B2(new_n763), .C1(new_n240), .C2(new_n791), .ZN(new_n1152));
  INV_X1    g0952(.A(G137), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n791), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n769), .A2(new_n983), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT53), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n273), .B1(new_n785), .B2(new_n782), .C1(new_n827), .C2(new_n831), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G125), .B2(new_n795), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT54), .B(G143), .Z(new_n1159));
  AOI22_X1  g0959(.A1(new_n824), .A2(G128), .B1(new_n775), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1005), .A2(G50), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1156), .A2(new_n1158), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1152), .B1(new_n1154), .B2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(new_n806), .B1(new_n301), .B2(new_n843), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n739), .B(new_n1164), .C1(new_n897), .C2(new_n840), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1113), .A2(new_n1147), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(G378));
  NAND2_X1  g0967(.A1(new_n373), .A2(new_n383), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n355), .A2(new_n847), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT55), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT56), .Z(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n744), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n843), .A2(new_n352), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1021), .B1(new_n824), .B2(G116), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n254), .B2(new_n782), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n790), .A2(G97), .B1(G107), .B2(new_n776), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n326), .B2(new_n774), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n760), .A2(new_n822), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n262), .B(new_n489), .C1(new_n971), .C2(new_n784), .ZN(new_n1180));
  NOR4_X1   g0980(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT58), .Z(new_n1182));
  OAI22_X1  g0982(.A1(new_n774), .A2(new_n1153), .B1(new_n983), .B2(new_n782), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n770), .A2(new_n1159), .ZN(new_n1184));
  INV_X1    g0984(.A(G128), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1184), .B1(new_n1185), .B2(new_n827), .C1(new_n791), .C2(new_n831), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1183), .B(new_n1186), .C1(G125), .C2(new_n824), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT59), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G33), .B1(new_n795), .B2(G124), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G41), .B1(new_n1005), .B2(G159), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n489), .B1(new_n258), .B2(new_n260), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n352), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1182), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n819), .B1(new_n1196), .B2(new_n806), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1173), .A2(new_n1174), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n884), .A2(G330), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n900), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n884), .A2(G330), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1202), .A2(new_n893), .A3(new_n894), .A4(new_n899), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1172), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1201), .A2(new_n1203), .A3(new_n1172), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1199), .B1(new_n1208), .B2(new_n738), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1121), .B(KEYINPUT122), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1138), .A2(new_n1210), .B1(new_n1207), .B2(new_n1206), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n689), .B1(new_n1211), .B2(KEYINPUT57), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1144), .A2(new_n1145), .B1(new_n1107), .B2(new_n1091), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1210), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1208), .B(KEYINPUT57), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1209), .B1(new_n1212), .B2(new_n1216), .ZN(G375));
  NAND2_X1  g1017(.A1(new_n1087), .A2(new_n744), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n827), .A2(new_n971), .B1(new_n217), .B2(new_n769), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G107), .B2(new_n775), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n341), .B1(new_n784), .B2(new_n799), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1024), .B(new_n1221), .C1(new_n790), .C2(G116), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n202), .B2(new_n763), .C1(new_n481), .C2(new_n779), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n314), .B1(new_n352), .B2(new_n782), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1225), .B(new_n1179), .C1(G132), .C2(new_n824), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n769), .A2(new_n785), .B1(new_n774), .B2(new_n983), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n827), .A2(new_n1153), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n790), .C2(new_n1159), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1226), .B(new_n1229), .C1(new_n1185), .C2(new_n784), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n743), .B1(new_n1224), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n254), .B2(new_n843), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1218), .A2(new_n739), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1143), .B2(new_n737), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1143), .A2(new_n1121), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1144), .A2(new_n1145), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1237), .B2(new_n938), .ZN(G381));
  NAND4_X1  g1038(.A1(new_n1113), .A2(new_n1209), .A3(new_n1147), .A4(new_n1165), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1208), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n690), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1239), .B1(new_n1215), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1039), .A2(new_n809), .A3(new_n1042), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1244), .A2(G381), .A3(G384), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1074), .A2(new_n968), .A3(new_n991), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT123), .ZN(G407));
  NAND2_X1  g1048(.A1(new_n1243), .A2(new_n669), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(G213), .A3(new_n1249), .ZN(G409));
  NAND2_X1  g1050(.A1(G375), .A2(G378), .ZN(new_n1251));
  INV_X1    g1051(.A(G213), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1252), .A2(G343), .ZN(new_n1253));
  AND4_X1   g1053(.A1(new_n1147), .A2(new_n1113), .A3(new_n1209), .A4(new_n1165), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1211), .A2(new_n937), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1253), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT60), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n1236), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n689), .B1(new_n1260), .B2(KEYINPUT60), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G384), .B(new_n1235), .C1(new_n1259), .C2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G384), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1261), .B1(new_n1237), .B2(KEYINPUT60), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1234), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1251), .A2(new_n1256), .A3(new_n1267), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1253), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1147), .A2(new_n1165), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1273), .A2(new_n1255), .A3(new_n1113), .A4(new_n1209), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1209), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1242), .B2(new_n1215), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1272), .B(new_n1274), .C1(new_n1276), .C2(new_n1166), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1262), .A2(new_n1265), .A3(KEYINPUT125), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1253), .A2(G2897), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1266), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1266), .A2(new_n1281), .A3(new_n1279), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1277), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G387), .A2(G390), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1244), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n809), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT126), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G393), .A2(G396), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT126), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1244), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1074), .A2(new_n968), .A3(new_n991), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1287), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1074), .B1(new_n968), .B2(new_n991), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1293), .B1(new_n1246), .B2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1286), .A2(new_n1296), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n689), .A3(new_n1215), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1166), .B1(new_n1301), .B2(new_n1209), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1240), .A2(new_n938), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1272), .B1(new_n1239), .B2(new_n1303), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1302), .A2(new_n1304), .A3(new_n1266), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT124), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1305), .A2(new_n1306), .A3(KEYINPUT63), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT63), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT124), .B1(new_n1268), .B2(new_n1308), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1251), .A2(new_n1256), .A3(KEYINPUT63), .A4(new_n1267), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1298), .A2(new_n1296), .ZN(new_n1312));
  AND4_X1   g1112(.A1(new_n1271), .A2(new_n1285), .A3(new_n1311), .A4(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT127), .B1(new_n1310), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1306), .B1(new_n1305), .B2(KEYINPUT63), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1268), .A2(KEYINPUT124), .A3(new_n1308), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1285), .A2(new_n1312), .A3(new_n1311), .A4(new_n1271), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1299), .B1(new_n1314), .B2(new_n1320), .ZN(G405));
  NOR2_X1   g1121(.A1(new_n1302), .A2(new_n1243), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(new_n1266), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1323), .B(new_n1312), .ZN(G402));
endmodule


