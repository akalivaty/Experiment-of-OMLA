

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U546 ( .A1(n756), .A2(n754), .ZN(n743) );
  AND2_X1 U547 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U548 ( .A(n759), .B(KEYINPUT100), .ZN(n772) );
  NAND2_X1 U549 ( .A1(n707), .A2(n706), .ZN(n762) );
  NOR2_X1 U550 ( .A1(n673), .A2(n672), .ZN(n706) );
  NOR2_X1 U551 ( .A1(G164), .A2(G1384), .ZN(n707) );
  NOR2_X1 U552 ( .A1(G651), .A2(n614), .ZN(n639) );
  NOR2_X1 U553 ( .A1(G2104), .A2(G2105), .ZN(n509) );
  XOR2_X2 U554 ( .A(KEYINPUT17), .B(n509), .Z(n875) );
  NAND2_X1 U555 ( .A1(G138), .A2(n875), .ZN(n512) );
  INV_X1 U556 ( .A(G2105), .ZN(n513) );
  AND2_X1 U557 ( .A1(G2104), .A2(n513), .ZN(n510) );
  XNOR2_X2 U558 ( .A(n510), .B(KEYINPUT64), .ZN(n876) );
  NAND2_X1 U559 ( .A1(G102), .A2(n876), .ZN(n511) );
  NAND2_X1 U560 ( .A1(n512), .A2(n511), .ZN(n517) );
  NOR2_X1 U561 ( .A1(G2104), .A2(n513), .ZN(n879) );
  NAND2_X1 U562 ( .A1(G126), .A2(n879), .ZN(n515) );
  AND2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  NAND2_X1 U564 ( .A1(G114), .A2(n881), .ZN(n514) );
  NAND2_X1 U565 ( .A1(n515), .A2(n514), .ZN(n516) );
  NOR2_X1 U566 ( .A1(n517), .A2(n516), .ZN(G164) );
  INV_X1 U567 ( .A(G651), .ZN(n520) );
  NOR2_X1 U568 ( .A1(G543), .A2(n520), .ZN(n518) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n518), .Z(n638) );
  NAND2_X1 U570 ( .A1(G65), .A2(n638), .ZN(n522) );
  XNOR2_X1 U571 ( .A(G543), .B(KEYINPUT0), .ZN(n519) );
  XNOR2_X1 U572 ( .A(n519), .B(KEYINPUT65), .ZN(n614) );
  NOR2_X1 U573 ( .A1(n614), .A2(n520), .ZN(n634) );
  NAND2_X1 U574 ( .A1(G78), .A2(n634), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n526) );
  NOR2_X1 U576 ( .A1(G651), .A2(G543), .ZN(n632) );
  NAND2_X1 U577 ( .A1(G91), .A2(n632), .ZN(n524) );
  NAND2_X1 U578 ( .A1(G53), .A2(n639), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n524), .A2(n523), .ZN(n525) );
  OR2_X1 U580 ( .A1(n526), .A2(n525), .ZN(G299) );
  XOR2_X1 U581 ( .A(G2451), .B(G2454), .Z(n528) );
  XNOR2_X1 U582 ( .A(G2430), .B(KEYINPUT104), .ZN(n527) );
  XNOR2_X1 U583 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U584 ( .A(n529), .B(G2446), .Z(n531) );
  XNOR2_X1 U585 ( .A(G1341), .B(G1348), .ZN(n530) );
  XNOR2_X1 U586 ( .A(n531), .B(n530), .ZN(n535) );
  XOR2_X1 U587 ( .A(G2438), .B(G2427), .Z(n533) );
  XNOR2_X1 U588 ( .A(G2443), .B(G2435), .ZN(n532) );
  XNOR2_X1 U589 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U590 ( .A(n535), .B(n534), .Z(n536) );
  AND2_X1 U591 ( .A1(G14), .A2(n536), .ZN(G401) );
  NAND2_X1 U592 ( .A1(G64), .A2(n638), .ZN(n538) );
  NAND2_X1 U593 ( .A1(G52), .A2(n639), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n543) );
  NAND2_X1 U595 ( .A1(G77), .A2(n634), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G90), .A2(n632), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n541), .Z(n542) );
  NOR2_X1 U599 ( .A1(n543), .A2(n542), .ZN(G171) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U601 ( .A1(n876), .A2(G101), .ZN(n544) );
  XOR2_X1 U602 ( .A(KEYINPUT23), .B(n544), .Z(n546) );
  NAND2_X1 U603 ( .A1(n879), .A2(G125), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n673) );
  NAND2_X1 U605 ( .A1(G137), .A2(n875), .ZN(n548) );
  NAND2_X1 U606 ( .A1(G113), .A2(n881), .ZN(n547) );
  NAND2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n671) );
  NOR2_X1 U608 ( .A1(n673), .A2(n671), .ZN(G160) );
  NAND2_X1 U609 ( .A1(n632), .A2(G89), .ZN(n549) );
  XNOR2_X1 U610 ( .A(n549), .B(KEYINPUT4), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G76), .A2(n634), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U613 ( .A(n552), .B(KEYINPUT5), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G63), .A2(n638), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G51), .A2(n639), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n555), .Z(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U619 ( .A(n558), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U623 ( .A(G223), .ZN(n816) );
  NAND2_X1 U624 ( .A1(n816), .A2(G567), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  NAND2_X1 U626 ( .A1(G56), .A2(n638), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT14), .B(n561), .Z(n568) );
  NAND2_X1 U628 ( .A1(n634), .A2(G68), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT69), .B(n562), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n632), .A2(G81), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT12), .B(n563), .Z(n564) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT13), .ZN(n567) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n639), .A2(G43), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n969) );
  XOR2_X1 U637 ( .A(G860), .B(KEYINPUT70), .Z(n584) );
  NOR2_X1 U638 ( .A1(n969), .A2(n584), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n571), .B(KEYINPUT71), .ZN(G153) );
  INV_X1 U640 ( .A(G171), .ZN(G301) );
  NAND2_X1 U641 ( .A1(G868), .A2(G301), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G66), .A2(n638), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G79), .A2(n634), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G92), .A2(n632), .ZN(n575) );
  NAND2_X1 U646 ( .A1(G54), .A2(n639), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U649 ( .A(KEYINPUT15), .B(n578), .Z(n960) );
  OR2_X1 U650 ( .A1(n960), .A2(G868), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(G284) );
  INV_X1 U652 ( .A(G868), .ZN(n581) );
  NOR2_X1 U653 ( .A1(G286), .A2(n581), .ZN(n583) );
  NOR2_X1 U654 ( .A1(G868), .A2(G299), .ZN(n582) );
  NOR2_X1 U655 ( .A1(n583), .A2(n582), .ZN(G297) );
  NAND2_X1 U656 ( .A1(n584), .A2(G559), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n585), .A2(n960), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n586), .B(KEYINPUT72), .ZN(n587) );
  XNOR2_X1 U659 ( .A(KEYINPUT16), .B(n587), .ZN(G148) );
  NOR2_X1 U660 ( .A1(G868), .A2(n969), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G868), .A2(n960), .ZN(n588) );
  NOR2_X1 U662 ( .A1(G559), .A2(n588), .ZN(n589) );
  NOR2_X1 U663 ( .A1(n590), .A2(n589), .ZN(G282) );
  XOR2_X1 U664 ( .A(G2100), .B(KEYINPUT76), .Z(n602) );
  NAND2_X1 U665 ( .A1(G123), .A2(n879), .ZN(n591) );
  XOR2_X1 U666 ( .A(KEYINPUT73), .B(n591), .Z(n592) );
  XNOR2_X1 U667 ( .A(n592), .B(KEYINPUT18), .ZN(n594) );
  NAND2_X1 U668 ( .A1(G135), .A2(n875), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U670 ( .A(KEYINPUT74), .B(n595), .ZN(n598) );
  NAND2_X1 U671 ( .A1(G99), .A2(n876), .ZN(n596) );
  XNOR2_X1 U672 ( .A(KEYINPUT75), .B(n596), .ZN(n597) );
  NOR2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n881), .A2(G111), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n909) );
  XOR2_X1 U676 ( .A(G2096), .B(n909), .Z(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(G156) );
  NAND2_X1 U678 ( .A1(G61), .A2(n638), .ZN(n604) );
  NAND2_X1 U679 ( .A1(G86), .A2(n632), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n634), .A2(G73), .ZN(n605) );
  XOR2_X1 U682 ( .A(KEYINPUT2), .B(n605), .Z(n606) );
  NOR2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n639), .A2(G48), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(G305) );
  NAND2_X1 U686 ( .A1(G49), .A2(n639), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G74), .A2(G651), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U689 ( .A(KEYINPUT80), .B(n612), .ZN(n613) );
  NOR2_X1 U690 ( .A1(n638), .A2(n613), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n614), .A2(G87), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(G288) );
  AND2_X1 U693 ( .A1(n638), .A2(G60), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G72), .A2(n634), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G85), .A2(n632), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n639), .A2(G47), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(G290) );
  NAND2_X1 U700 ( .A1(G75), .A2(n634), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G88), .A2(n632), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(KEYINPUT82), .B(n625), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G62), .A2(n638), .ZN(n626) );
  XNOR2_X1 U705 ( .A(KEYINPUT81), .B(n626), .ZN(n627) );
  NOR2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n639), .A2(G50), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(G303) );
  INV_X1 U709 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U710 ( .A(G299), .B(G305), .ZN(n631) );
  XNOR2_X1 U711 ( .A(n631), .B(G288), .ZN(n649) );
  NAND2_X1 U712 ( .A1(n632), .A2(G93), .ZN(n633) );
  XOR2_X1 U713 ( .A(KEYINPUT77), .B(n633), .Z(n636) );
  NAND2_X1 U714 ( .A1(n634), .A2(G80), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U716 ( .A(KEYINPUT78), .B(n637), .ZN(n643) );
  NAND2_X1 U717 ( .A1(G67), .A2(n638), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G55), .A2(n639), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U721 ( .A(KEYINPUT79), .B(n644), .Z(n825) );
  XNOR2_X1 U722 ( .A(n825), .B(KEYINPUT19), .ZN(n646) );
  XNOR2_X1 U723 ( .A(G290), .B(G166), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n646), .B(n645), .ZN(n647) );
  XOR2_X1 U725 ( .A(n647), .B(n969), .Z(n648) );
  XNOR2_X1 U726 ( .A(n649), .B(n648), .ZN(n896) );
  NAND2_X1 U727 ( .A1(n960), .A2(G559), .ZN(n823) );
  XNOR2_X1 U728 ( .A(n896), .B(n823), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n650), .A2(G868), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n651), .B(KEYINPUT83), .ZN(n653) );
  NOR2_X1 U731 ( .A1(n825), .A2(G868), .ZN(n652) );
  NOR2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U733 ( .A(KEYINPUT84), .B(n654), .Z(G295) );
  NAND2_X1 U734 ( .A1(G2078), .A2(G2084), .ZN(n655) );
  XOR2_X1 U735 ( .A(KEYINPUT20), .B(n655), .Z(n656) );
  NAND2_X1 U736 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U737 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n658), .A2(G2072), .ZN(G158) );
  XOR2_X1 U739 ( .A(KEYINPUT66), .B(G57), .Z(G237) );
  XNOR2_X1 U740 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U741 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  XNOR2_X1 U742 ( .A(KEYINPUT67), .B(G132), .ZN(G219) );
  NAND2_X1 U743 ( .A1(G108), .A2(G120), .ZN(n659) );
  NOR2_X1 U744 ( .A1(G237), .A2(n659), .ZN(n660) );
  NAND2_X1 U745 ( .A1(G69), .A2(n660), .ZN(n822) );
  NAND2_X1 U746 ( .A1(G567), .A2(n822), .ZN(n666) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n661) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n661), .Z(n662) );
  NOR2_X1 U749 ( .A1(G218), .A2(n662), .ZN(n663) );
  NAND2_X1 U750 ( .A1(G96), .A2(n663), .ZN(n821) );
  NAND2_X1 U751 ( .A1(G2106), .A2(n821), .ZN(n664) );
  XOR2_X1 U752 ( .A(KEYINPUT85), .B(n664), .Z(n665) );
  NAND2_X1 U753 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U754 ( .A(KEYINPUT86), .B(n667), .Z(G319) );
  INV_X1 U755 ( .A(G319), .ZN(n669) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n668) );
  NOR2_X1 U757 ( .A1(n669), .A2(n668), .ZN(n820) );
  NAND2_X1 U758 ( .A1(n820), .A2(G36), .ZN(G176) );
  XNOR2_X1 U759 ( .A(G1986), .B(G290), .ZN(n964) );
  INV_X1 U760 ( .A(G40), .ZN(n670) );
  OR2_X1 U761 ( .A1(n671), .A2(n670), .ZN(n672) );
  INV_X1 U762 ( .A(n706), .ZN(n674) );
  NOR2_X1 U763 ( .A1(n707), .A2(n674), .ZN(n810) );
  NAND2_X1 U764 ( .A1(n964), .A2(n810), .ZN(n798) );
  NAND2_X1 U765 ( .A1(G140), .A2(n875), .ZN(n676) );
  NAND2_X1 U766 ( .A1(G104), .A2(n876), .ZN(n675) );
  NAND2_X1 U767 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U768 ( .A(KEYINPUT34), .B(n677), .ZN(n682) );
  NAND2_X1 U769 ( .A1(G128), .A2(n879), .ZN(n679) );
  NAND2_X1 U770 ( .A1(G116), .A2(n881), .ZN(n678) );
  NAND2_X1 U771 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U772 ( .A(KEYINPUT35), .B(n680), .Z(n681) );
  NOR2_X1 U773 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U774 ( .A(KEYINPUT36), .B(n683), .ZN(n872) );
  XOR2_X1 U775 ( .A(G2067), .B(KEYINPUT37), .Z(n684) );
  XNOR2_X1 U776 ( .A(KEYINPUT87), .B(n684), .ZN(n799) );
  NOR2_X1 U777 ( .A1(n872), .A2(n799), .ZN(n925) );
  NAND2_X1 U778 ( .A1(n810), .A2(n925), .ZN(n807) );
  NAND2_X1 U779 ( .A1(G107), .A2(n881), .ZN(n685) );
  XNOR2_X1 U780 ( .A(n685), .B(KEYINPUT88), .ZN(n687) );
  NAND2_X1 U781 ( .A1(n879), .A2(G119), .ZN(n686) );
  NAND2_X1 U782 ( .A1(n687), .A2(n686), .ZN(n691) );
  NAND2_X1 U783 ( .A1(G131), .A2(n875), .ZN(n689) );
  NAND2_X1 U784 ( .A1(G95), .A2(n876), .ZN(n688) );
  NAND2_X1 U785 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U786 ( .A1(n691), .A2(n690), .ZN(n889) );
  XNOR2_X1 U787 ( .A(KEYINPUT89), .B(G1991), .ZN(n936) );
  NOR2_X1 U788 ( .A1(n889), .A2(n936), .ZN(n701) );
  NAND2_X1 U789 ( .A1(G129), .A2(n879), .ZN(n693) );
  NAND2_X1 U790 ( .A1(G117), .A2(n881), .ZN(n692) );
  NAND2_X1 U791 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U792 ( .A(KEYINPUT90), .B(n694), .ZN(n697) );
  NAND2_X1 U793 ( .A1(G105), .A2(n876), .ZN(n695) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n695), .Z(n696) );
  NOR2_X1 U795 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U796 ( .A1(n875), .A2(G141), .ZN(n698) );
  NAND2_X1 U797 ( .A1(n699), .A2(n698), .ZN(n871) );
  AND2_X1 U798 ( .A1(n871), .A2(G1996), .ZN(n700) );
  NOR2_X1 U799 ( .A1(n701), .A2(n700), .ZN(n905) );
  XNOR2_X1 U800 ( .A(KEYINPUT91), .B(n810), .ZN(n702) );
  NOR2_X1 U801 ( .A1(n905), .A2(n702), .ZN(n803) );
  INV_X1 U802 ( .A(n803), .ZN(n703) );
  NAND2_X1 U803 ( .A1(n807), .A2(n703), .ZN(n796) );
  NAND2_X1 U804 ( .A1(G8), .A2(n762), .ZN(n789) );
  NOR2_X1 U805 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XOR2_X1 U806 ( .A(n704), .B(KEYINPUT24), .Z(n705) );
  NOR2_X1 U807 ( .A1(n789), .A2(n705), .ZN(n794) );
  NOR2_X1 U808 ( .A1(n709), .A2(G1961), .ZN(n711) );
  XOR2_X1 U809 ( .A(G2078), .B(KEYINPUT25), .Z(n937) );
  INV_X1 U810 ( .A(KEYINPUT93), .ZN(n708) );
  XNOR2_X1 U811 ( .A(n709), .B(n708), .ZN(n719) );
  INV_X1 U812 ( .A(n719), .ZN(n715) );
  NOR2_X1 U813 ( .A1(n937), .A2(n715), .ZN(n710) );
  NOR2_X1 U814 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U815 ( .A(n712), .B(KEYINPUT94), .Z(n747) );
  AND2_X1 U816 ( .A1(G171), .A2(n747), .ZN(n713) );
  XOR2_X1 U817 ( .A(KEYINPUT95), .B(n713), .Z(n741) );
  NAND2_X1 U818 ( .A1(n719), .A2(G2072), .ZN(n714) );
  XOR2_X1 U819 ( .A(KEYINPUT27), .B(n714), .Z(n717) );
  NAND2_X1 U820 ( .A1(G1956), .A2(n715), .ZN(n716) );
  NAND2_X1 U821 ( .A1(n717), .A2(n716), .ZN(n729) );
  NAND2_X1 U822 ( .A1(G299), .A2(n729), .ZN(n718) );
  XOR2_X1 U823 ( .A(KEYINPUT28), .B(n718), .Z(n737) );
  NAND2_X1 U824 ( .A1(G2067), .A2(n719), .ZN(n721) );
  NAND2_X1 U825 ( .A1(G1348), .A2(n762), .ZN(n720) );
  NAND2_X1 U826 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U827 ( .A(n722), .B(KEYINPUT96), .ZN(n728) );
  INV_X1 U828 ( .A(G1996), .ZN(n932) );
  NOR2_X1 U829 ( .A1(n762), .A2(n932), .ZN(n723) );
  XOR2_X1 U830 ( .A(n723), .B(KEYINPUT26), .Z(n725) );
  NAND2_X1 U831 ( .A1(n762), .A2(G1341), .ZN(n724) );
  NAND2_X1 U832 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U833 ( .A1(n969), .A2(n726), .ZN(n731) );
  NOR2_X1 U834 ( .A1(n960), .A2(n731), .ZN(n727) );
  NOR2_X1 U835 ( .A1(n728), .A2(n727), .ZN(n735) );
  NOR2_X1 U836 ( .A1(G299), .A2(n729), .ZN(n730) );
  XNOR2_X1 U837 ( .A(n730), .B(KEYINPUT97), .ZN(n733) );
  NAND2_X1 U838 ( .A1(n731), .A2(n960), .ZN(n732) );
  NAND2_X1 U839 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U840 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U841 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U842 ( .A(KEYINPUT29), .B(n738), .ZN(n739) );
  INV_X1 U843 ( .A(n739), .ZN(n740) );
  NOR2_X1 U844 ( .A1(n741), .A2(n740), .ZN(n752) );
  NOR2_X1 U845 ( .A1(G2084), .A2(n762), .ZN(n756) );
  NOR2_X1 U846 ( .A1(G1966), .A2(n789), .ZN(n742) );
  XNOR2_X1 U847 ( .A(KEYINPUT92), .B(n742), .ZN(n754) );
  XNOR2_X1 U848 ( .A(KEYINPUT98), .B(n743), .ZN(n744) );
  NAND2_X1 U849 ( .A1(n744), .A2(G8), .ZN(n745) );
  XNOR2_X1 U850 ( .A(KEYINPUT30), .B(n745), .ZN(n746) );
  NOR2_X1 U851 ( .A1(G168), .A2(n746), .ZN(n749) );
  NOR2_X1 U852 ( .A1(G171), .A2(n747), .ZN(n748) );
  NOR2_X1 U853 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U854 ( .A(n750), .B(KEYINPUT31), .ZN(n751) );
  NOR2_X1 U855 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U856 ( .A(n753), .B(KEYINPUT99), .ZN(n761) );
  INV_X1 U857 ( .A(n754), .ZN(n755) );
  AND2_X1 U858 ( .A1(n761), .A2(n755), .ZN(n758) );
  NAND2_X1 U859 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U860 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U861 ( .A1(G286), .A2(G8), .ZN(n760) );
  NAND2_X1 U862 ( .A1(n761), .A2(n760), .ZN(n769) );
  INV_X1 U863 ( .A(G8), .ZN(n767) );
  NOR2_X1 U864 ( .A1(G1971), .A2(n789), .ZN(n764) );
  NOR2_X1 U865 ( .A1(G2090), .A2(n762), .ZN(n763) );
  NOR2_X1 U866 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U867 ( .A1(n765), .A2(G303), .ZN(n766) );
  OR2_X1 U868 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U869 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U870 ( .A(KEYINPUT32), .B(n770), .ZN(n771) );
  NAND2_X1 U871 ( .A1(n772), .A2(n771), .ZN(n788) );
  NOR2_X1 U872 ( .A1(G1976), .A2(G288), .ZN(n780) );
  NOR2_X1 U873 ( .A1(G1971), .A2(G303), .ZN(n773) );
  NOR2_X1 U874 ( .A1(n780), .A2(n773), .ZN(n958) );
  INV_X1 U875 ( .A(KEYINPUT33), .ZN(n777) );
  AND2_X1 U876 ( .A1(n958), .A2(n777), .ZN(n774) );
  AND2_X1 U877 ( .A1(n788), .A2(n774), .ZN(n779) );
  NAND2_X1 U878 ( .A1(G1976), .A2(G288), .ZN(n965) );
  INV_X1 U879 ( .A(n789), .ZN(n775) );
  NAND2_X1 U880 ( .A1(n965), .A2(n775), .ZN(n776) );
  AND2_X1 U881 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U882 ( .A1(n779), .A2(n778), .ZN(n785) );
  XOR2_X1 U883 ( .A(G1981), .B(G305), .Z(n955) );
  INV_X1 U884 ( .A(n955), .ZN(n783) );
  NAND2_X1 U885 ( .A1(n780), .A2(KEYINPUT33), .ZN(n781) );
  NOR2_X1 U886 ( .A1(n789), .A2(n781), .ZN(n782) );
  NOR2_X1 U887 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U888 ( .A1(n785), .A2(n784), .ZN(n792) );
  NOR2_X1 U889 ( .A1(G2090), .A2(G303), .ZN(n786) );
  NAND2_X1 U890 ( .A1(G8), .A2(n786), .ZN(n787) );
  NAND2_X1 U891 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U892 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U893 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U894 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U895 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U896 ( .A1(n798), .A2(n797), .ZN(n813) );
  NAND2_X1 U897 ( .A1(n872), .A2(n799), .ZN(n922) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n871), .ZN(n916) );
  AND2_X1 U899 ( .A1(n936), .A2(n889), .ZN(n908) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n800) );
  XOR2_X1 U901 ( .A(n800), .B(KEYINPUT101), .Z(n801) );
  NOR2_X1 U902 ( .A1(n908), .A2(n801), .ZN(n802) );
  NOR2_X1 U903 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U904 ( .A1(n916), .A2(n804), .ZN(n805) );
  XNOR2_X1 U905 ( .A(KEYINPUT39), .B(n805), .ZN(n806) );
  XNOR2_X1 U906 ( .A(n806), .B(KEYINPUT102), .ZN(n808) );
  NAND2_X1 U907 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U908 ( .A1(n922), .A2(n809), .ZN(n811) );
  NAND2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n815) );
  XOR2_X1 U911 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n814) );
  XNOR2_X1 U912 ( .A(n815), .B(n814), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U915 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n818) );
  XOR2_X1 U917 ( .A(KEYINPUT105), .B(n818), .Z(n819) );
  NAND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(G188) );
  XOR2_X1 U919 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G108), .ZN(G238) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n822), .A2(n821), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U926 ( .A(n969), .B(n823), .ZN(n824) );
  NOR2_X1 U927 ( .A1(n824), .A2(G860), .ZN(n826) );
  XNOR2_X1 U928 ( .A(n826), .B(n825), .ZN(G145) );
  XOR2_X1 U929 ( .A(KEYINPUT42), .B(G2090), .Z(n828) );
  XNOR2_X1 U930 ( .A(G2067), .B(G2084), .ZN(n827) );
  XNOR2_X1 U931 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U932 ( .A(n829), .B(G2096), .Z(n831) );
  XNOR2_X1 U933 ( .A(G2072), .B(G2078), .ZN(n830) );
  XNOR2_X1 U934 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U935 ( .A(G2100), .B(KEYINPUT43), .Z(n833) );
  XNOR2_X1 U936 ( .A(G2678), .B(KEYINPUT107), .ZN(n832) );
  XNOR2_X1 U937 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U938 ( .A(n835), .B(n834), .Z(G227) );
  XOR2_X1 U939 ( .A(G1981), .B(G1966), .Z(n837) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U941 ( .A(n837), .B(n836), .ZN(n847) );
  XOR2_X1 U942 ( .A(KEYINPUT110), .B(G2474), .Z(n839) );
  XNOR2_X1 U943 ( .A(G1956), .B(KEYINPUT108), .ZN(n838) );
  XNOR2_X1 U944 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U945 ( .A(G1976), .B(G1971), .Z(n841) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1961), .ZN(n840) );
  XNOR2_X1 U947 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U948 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U949 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n844) );
  XNOR2_X1 U950 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U951 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U952 ( .A1(G136), .A2(n875), .ZN(n848) );
  XNOR2_X1 U953 ( .A(n848), .B(KEYINPUT112), .ZN(n852) );
  XOR2_X1 U954 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n850) );
  NAND2_X1 U955 ( .A1(G124), .A2(n879), .ZN(n849) );
  XNOR2_X1 U956 ( .A(n850), .B(n849), .ZN(n851) );
  NAND2_X1 U957 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n881), .A2(G112), .ZN(n854) );
  NAND2_X1 U959 ( .A1(G100), .A2(n876), .ZN(n853) );
  NAND2_X1 U960 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U961 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U962 ( .A1(G130), .A2(n879), .ZN(n858) );
  NAND2_X1 U963 ( .A1(G118), .A2(n881), .ZN(n857) );
  NAND2_X1 U964 ( .A1(n858), .A2(n857), .ZN(n865) );
  XNOR2_X1 U965 ( .A(KEYINPUT114), .B(KEYINPUT45), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n875), .A2(G142), .ZN(n861) );
  NAND2_X1 U967 ( .A1(G106), .A2(n876), .ZN(n859) );
  XOR2_X1 U968 ( .A(KEYINPUT113), .B(n859), .Z(n860) );
  NAND2_X1 U969 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U970 ( .A(n863), .B(n862), .Z(n864) );
  NOR2_X1 U971 ( .A1(n865), .A2(n864), .ZN(n893) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n866) );
  XNOR2_X1 U973 ( .A(n909), .B(n866), .ZN(n867) );
  XOR2_X1 U974 ( .A(n867), .B(KEYINPUT118), .Z(n869) );
  XNOR2_X1 U975 ( .A(G164), .B(KEYINPUT117), .ZN(n868) );
  XNOR2_X1 U976 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U977 ( .A(G162), .B(n870), .ZN(n874) );
  XOR2_X1 U978 ( .A(n872), .B(n871), .Z(n873) );
  XNOR2_X1 U979 ( .A(n874), .B(n873), .ZN(n888) );
  NAND2_X1 U980 ( .A1(G139), .A2(n875), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G103), .A2(n876), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n887) );
  NAND2_X1 U983 ( .A1(n879), .A2(G127), .ZN(n880) );
  XNOR2_X1 U984 ( .A(KEYINPUT115), .B(n880), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n881), .A2(G115), .ZN(n882) );
  XOR2_X1 U986 ( .A(KEYINPUT116), .B(n882), .Z(n883) );
  NOR2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n885), .B(KEYINPUT47), .ZN(n886) );
  NOR2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n911) );
  XOR2_X1 U990 ( .A(n888), .B(n911), .Z(n891) );
  XNOR2_X1 U991 ( .A(G160), .B(n889), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U993 ( .A(n893), .B(n892), .Z(n894) );
  NOR2_X1 U994 ( .A1(G37), .A2(n894), .ZN(G395) );
  XOR2_X1 U995 ( .A(n960), .B(G286), .Z(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U997 ( .A(G301), .B(n897), .Z(n898) );
  NOR2_X1 U998 ( .A1(G37), .A2(n898), .ZN(n899) );
  XOR2_X1 U999 ( .A(KEYINPUT119), .B(n899), .Z(G397) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n900), .ZN(n901) );
  NOR2_X1 U1002 ( .A1(G401), .A2(n901), .ZN(n902) );
  AND2_X1 U1003 ( .A1(n902), .A2(G319), .ZN(n904) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n903) );
  NAND2_X1 U1005 ( .A1(n904), .A2(n903), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1007 ( .A(KEYINPUT52), .B(KEYINPUT120), .ZN(n927) );
  XNOR2_X1 U1008 ( .A(G160), .B(G2084), .ZN(n906) );
  NAND2_X1 U1009 ( .A1(n906), .A2(n905), .ZN(n907) );
  NOR2_X1 U1010 ( .A1(n908), .A2(n907), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(n921) );
  XOR2_X1 U1012 ( .A(G2072), .B(n911), .Z(n913) );
  XOR2_X1 U1013 ( .A(G164), .B(G2078), .Z(n912) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(KEYINPUT50), .B(n914), .ZN(n919) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n915) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1018 ( .A(KEYINPUT51), .B(n917), .Z(n918) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n927), .B(n926), .ZN(n929) );
  INV_X1 U1024 ( .A(KEYINPUT55), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n930), .A2(G29), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT121), .B(n931), .Z(n1009) );
  XNOR2_X1 U1028 ( .A(G29), .B(KEYINPUT123), .ZN(n953) );
  XNOR2_X1 U1029 ( .A(G32), .B(n932), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(G28), .ZN(n943) );
  XNOR2_X1 U1031 ( .A(G2067), .B(G26), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(G33), .B(G2072), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n941) );
  XOR2_X1 U1034 ( .A(n936), .B(G25), .Z(n939) );
  XNOR2_X1 U1035 ( .A(G27), .B(n937), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1039 ( .A(KEYINPUT53), .B(n944), .Z(n947) );
  XOR2_X1 U1040 ( .A(KEYINPUT54), .B(G34), .Z(n945) );
  XNOR2_X1 U1041 ( .A(G2084), .B(n945), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(KEYINPUT122), .B(G2090), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G35), .B(n948), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT55), .B(n951), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(G11), .A2(n954), .ZN(n1007) );
  XNOR2_X1 U1049 ( .A(G16), .B(KEYINPUT56), .ZN(n977) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G168), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(n957), .B(KEYINPUT57), .ZN(n975) );
  XNOR2_X1 U1053 ( .A(G171), .B(G1961), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n973) );
  XNOR2_X1 U1055 ( .A(n960), .B(G1348), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(G1971), .A2(G303), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(G1956), .B(G299), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n971) );
  XOR2_X1 U1062 ( .A(G1341), .B(n969), .Z(n970) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n1005) );
  INV_X1 U1067 ( .A(G16), .ZN(n1003) );
  XOR2_X1 U1068 ( .A(G1348), .B(KEYINPUT59), .Z(n978) );
  XNOR2_X1 U1069 ( .A(G4), .B(n978), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(G20), .B(G1956), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G1341), .B(G19), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G1981), .B(G6), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(n985), .B(KEYINPUT60), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(KEYINPUT125), .B(n986), .ZN(n997) );
  XNOR2_X1 U1078 ( .A(G1961), .B(KEYINPUT124), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(n987), .B(G5), .ZN(n995) );
  XNOR2_X1 U1080 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n993) );
  XOR2_X1 U1081 ( .A(G1986), .B(G24), .Z(n991) );
  XNOR2_X1 U1082 ( .A(G1971), .B(G22), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(G23), .B(G1976), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1086 ( .A(n993), .B(n992), .Z(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(KEYINPUT126), .B(G1966), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(G21), .B(n998), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(KEYINPUT61), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(KEYINPUT62), .B(n1010), .Z(G311) );
  INV_X1 U1098 ( .A(G311), .ZN(G150) );
endmodule

