//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n453), .B(new_n454), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n455), .A2(new_n460), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n468), .A2(new_n469), .A3(G137), .A4(new_n470), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n465), .A2(new_n467), .A3(G137), .A4(new_n470), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT69), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n471), .A2(new_n473), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n465), .A2(new_n467), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n479), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n475), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT70), .ZN(G160));
  NOR2_X1   g060(.A1(new_n477), .A2(new_n470), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n477), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n465), .A2(new_n467), .A3(G126), .A4(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n468), .A2(new_n498), .A3(G138), .A4(new_n470), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n470), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(G50), .A2(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT71), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n508), .A2(new_n520), .A3(G62), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n511), .B1(new_n522), .B2(G651), .ZN(G166));
  NOR2_X1   g098(.A1(new_n505), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT72), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n504), .A2(new_n506), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n526), .A2(G543), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT73), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n526), .A2(new_n531), .A3(G543), .A4(new_n528), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n530), .A2(G51), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT6), .B(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n516), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n533), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n533), .A2(KEYINPUT74), .A3(new_n536), .A4(new_n538), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G168));
  NAND3_X1  g118(.A1(new_n530), .A2(G52), .A3(new_n532), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n503), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n516), .A2(new_n507), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND3_X1  g125(.A1(new_n530), .A2(G43), .A3(new_n532), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(G81), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT75), .B1(new_n553), .B2(new_n503), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n516), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n557), .A2(new_n558), .A3(G651), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n551), .A2(new_n552), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n551), .A2(KEYINPUT76), .A3(new_n560), .A4(new_n552), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  AND2_X1   g146(.A1(new_n526), .A2(new_n528), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  XOR2_X1   g149(.A(KEYINPUT77), .B(G65), .Z(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n516), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(new_n547), .B2(G91), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n529), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n573), .A2(new_n577), .A3(new_n580), .ZN(G299));
  INV_X1    g156(.A(G168), .ZN(G286));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n583));
  AOI211_X1 g158(.A(new_n583), .B(new_n511), .C1(G651), .C2(new_n522), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n522), .A2(G651), .ZN(new_n585));
  INV_X1    g160(.A(new_n511), .ZN(new_n586));
  AOI21_X1  g161(.A(KEYINPUT78), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n584), .A2(new_n587), .ZN(G303));
  NAND3_X1  g163(.A1(new_n572), .A2(G49), .A3(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n547), .A2(G87), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n516), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G48), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n516), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(G651), .A2(new_n595), .B1(new_n598), .B2(new_n534), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G305));
  NAND3_X1  g175(.A1(new_n530), .A2(G47), .A3(new_n532), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n503), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n547), .A2(G85), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(G290));
  NAND3_X1  g180(.A1(new_n530), .A2(G54), .A3(new_n532), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT80), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n513), .A2(new_n515), .A3(G66), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n503), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n508), .A2(new_n534), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n611), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n615), .A2(G92), .A3(new_n508), .A4(new_n534), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n610), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n606), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G171), .B2(new_n619), .ZN(G284));
  OAI21_X1  g196(.A(new_n620), .B1(G171), .B2(new_n619), .ZN(G321));
  NAND2_X1  g197(.A1(G299), .A2(new_n619), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G168), .B2(new_n619), .ZN(G297));
  XOR2_X1   g199(.A(G297), .B(KEYINPUT81), .Z(G280));
  INV_X1    g200(.A(new_n618), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  NOR2_X1   g203(.A1(new_n618), .A2(G559), .ZN(new_n629));
  MUX2_X1   g204(.A(new_n629), .B(new_n565), .S(new_n619), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT82), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n468), .A2(new_n474), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  AOI22_X1  g212(.A1(G123), .A2(new_n486), .B1(new_n488), .B2(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n641), .B(new_n642), .C1(G111), .C2(new_n470), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n637), .A2(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT15), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2435), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(G2435), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2443), .B(G2446), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(KEYINPUT85), .B2(KEYINPUT17), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n667), .B(new_n668), .C1(KEYINPUT85), .C2(KEYINPUT17), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(G2072), .A2(G2078), .ZN(new_n672));
  OAI22_X1  g247(.A1(new_n666), .A2(new_n670), .B1(new_n444), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(G227));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n687), .B(new_n688), .C1(new_n686), .C2(new_n685), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  INV_X1    g267(.A(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n691), .B(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G16), .A2(G23), .ZN(new_n697));
  INV_X1    g272(.A(G288), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT33), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G1971), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G6), .A2(G16), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n599), .B2(G16), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n701), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  NOR2_X1   g287(.A1(G16), .A2(G24), .ZN(new_n713));
  INV_X1    g288(.A(G290), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G16), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT87), .B(G1986), .Z(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n716), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(KEYINPUT88), .B1(new_n711), .B2(KEYINPUT34), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n718), .B(new_n719), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n486), .A2(G119), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n488), .A2(G131), .ZN(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n470), .A2(G107), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n725), .B(new_n726), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G25), .B(new_n729), .S(G29), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT35), .B(G1991), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT86), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  OR3_X1    g308(.A1(new_n724), .A2(KEYINPUT36), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT36), .B1(new_n724), .B2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G34), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(KEYINPUT91), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(KEYINPUT91), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n740), .B(new_n741), .C1(new_n738), .C2(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G160), .B2(G29), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G2084), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT97), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n702), .A2(G5), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G171), .B2(new_n702), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT96), .Z(new_n748));
  INV_X1    g323(.A(G1961), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n486), .A2(G129), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n474), .A2(G105), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT26), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n488), .A2(G141), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n752), .A2(new_n753), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G32), .B(new_n757), .S(G29), .Z(new_n758));
  XOR2_X1   g333(.A(KEYINPUT27), .B(G1996), .Z(new_n759));
  AOI22_X1  g334(.A1(new_n748), .A2(new_n749), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n745), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT98), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT28), .ZN(new_n764));
  INV_X1    g339(.A(G26), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G29), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(G29), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n486), .A2(G128), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n488), .A2(G140), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n470), .A2(G116), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n769), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n767), .B1(new_n772), .B2(G29), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n766), .B1(new_n773), .B2(new_n764), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G2067), .ZN(new_n775));
  NOR2_X1   g350(.A1(G27), .A2(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G164), .B2(G29), .ZN(new_n777));
  OAI221_X1 g352(.A(new_n775), .B1(G2078), .B2(new_n777), .C1(new_n758), .C2(new_n759), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G29), .B2(G33), .ZN(new_n780));
  OR3_X1    g355(.A1(new_n779), .A2(G29), .A3(G33), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n474), .A2(G103), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT25), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n488), .A2(G139), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n783), .B(new_n784), .C1(new_n470), .C2(new_n785), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n780), .B(new_n781), .C1(new_n786), .C2(new_n737), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(new_n442), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT90), .Z(new_n789));
  NOR2_X1   g364(.A1(new_n778), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G11), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n737), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n737), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT29), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G2090), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n702), .A2(G21), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G168), .B2(new_n702), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n790), .B(new_n798), .C1(G1966), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n702), .A2(G19), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n565), .B2(new_n702), .ZN(new_n803));
  OAI22_X1  g378(.A1(new_n748), .A2(new_n749), .B1(new_n803), .B2(G1341), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n800), .A2(G1966), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n743), .A2(G2084), .ZN(new_n807));
  INV_X1    g382(.A(G28), .ZN(new_n808));
  AOI21_X1  g383(.A(G29), .B1(new_n808), .B2(KEYINPUT30), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(KEYINPUT30), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT95), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n777), .A2(G2078), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n702), .A2(G4), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n626), .B2(new_n702), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G1348), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n807), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n702), .A2(KEYINPUT23), .A3(G20), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT23), .ZN(new_n818));
  INV_X1    g393(.A(G20), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(G16), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n573), .A2(new_n577), .A3(new_n580), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n817), .B(new_n820), .C1(new_n821), .C2(new_n702), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1956), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G2090), .B2(new_n795), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT99), .ZN(new_n825));
  AOI211_X1 g400(.A(new_n806), .B(new_n816), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n814), .A2(G1348), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n824), .A2(new_n825), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G1341), .B2(new_n803), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n805), .A2(new_n826), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n763), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n638), .A2(G29), .A3(new_n643), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n787), .A2(new_n442), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT92), .Z(new_n834));
  NAND4_X1  g409(.A1(new_n736), .A2(new_n831), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n774), .A2(G2067), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n837), .ZN(G311));
  INV_X1    g413(.A(G311), .ZN(G150));
  NAND3_X1  g414(.A1(new_n530), .A2(G55), .A3(new_n532), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(new_n503), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n547), .A2(G93), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  INV_X1    g421(.A(new_n844), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n563), .B2(new_n564), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n847), .A2(new_n561), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n626), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n846), .B1(new_n854), .B2(G860), .ZN(G145));
  XOR2_X1   g430(.A(new_n757), .B(new_n786), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n772), .B(G164), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n856), .B(new_n857), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n635), .B(new_n729), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n486), .A2(G130), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n488), .A2(G142), .ZN(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(G2104), .C1(G118), .C2(new_n470), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n859), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT100), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT101), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n858), .A2(new_n866), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G160), .B(new_n644), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n492), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(G37), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n858), .A2(new_n866), .ZN(new_n874));
  INV_X1    g449(.A(new_n865), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n874), .B(new_n871), .C1(new_n858), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n847), .B2(G868), .ZN(new_n880));
  INV_X1    g455(.A(new_n629), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n850), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n848), .A2(new_n849), .A3(new_n629), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT102), .B1(new_n606), .B2(new_n617), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n606), .A2(KEYINPUT102), .A3(new_n617), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(G299), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n626), .A2(new_n821), .A3(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT103), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n606), .A2(KEYINPUT102), .A3(new_n617), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n892), .A2(new_n885), .A3(new_n821), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n618), .A2(G299), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT41), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n888), .A2(new_n897), .A3(new_n889), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n884), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n901));
  INV_X1    g476(.A(new_n890), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n901), .B(new_n902), .C1(new_n882), .C2(new_n883), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n891), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n891), .A2(new_n906), .A3(new_n900), .A4(new_n903), .ZN(new_n907));
  XNOR2_X1  g482(.A(G305), .B(G166), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n714), .A2(G288), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n698), .A2(G290), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n911), .B1(new_n909), .B2(new_n910), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n913), .A2(new_n908), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n905), .A2(new_n907), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n905), .B2(new_n907), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n880), .B1(new_n920), .B2(G868), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n918), .A2(new_n919), .A3(new_n619), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(KEYINPUT105), .B2(new_n922), .ZN(G295));
  AOI21_X1  g498(.A(new_n921), .B1(KEYINPUT105), .B2(new_n922), .ZN(G331));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n565), .A2(new_n844), .ZN(new_n926));
  NAND2_X1  g501(.A1(G168), .A2(G171), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n847), .A2(new_n561), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n541), .A2(new_n542), .A3(G301), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n926), .A2(new_n927), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n541), .A2(new_n542), .A3(G301), .ZN(new_n931));
  AOI21_X1  g506(.A(G301), .B1(new_n541), .B2(new_n542), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n931), .A2(new_n932), .B1(new_n848), .B2(new_n849), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n899), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n890), .B1(new_n930), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n936), .B2(new_n916), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n933), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n902), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n896), .A2(KEYINPUT106), .A3(new_n898), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n890), .A2(new_n941), .A3(KEYINPUT41), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n940), .A2(new_n930), .A3(new_n933), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n916), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT107), .B1(new_n937), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n899), .A2(new_n930), .A3(new_n933), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n939), .A2(new_n916), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G37), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n950), .A2(new_n951), .A3(new_n944), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n917), .B1(new_n934), .B2(new_n935), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n954), .A2(new_n949), .A3(new_n948), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n925), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n937), .A2(new_n956), .A3(new_n945), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n925), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT108), .B1(new_n958), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n965));
  INV_X1    g540(.A(new_n957), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n937), .A2(KEYINPUT107), .A3(new_n945), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n951), .B1(new_n950), .B2(new_n944), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n969), .B2(KEYINPUT43), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n965), .B(new_n962), .C1(new_n970), .C2(new_n925), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n964), .A2(new_n971), .ZN(G397));
  XNOR2_X1  g547(.A(KEYINPUT109), .B(G1384), .ZN(new_n973));
  NOR2_X1   g548(.A1(G164), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n475), .A2(new_n482), .A3(G40), .A4(new_n483), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G2067), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n772), .B(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT111), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n979), .B1(new_n983), .B2(new_n757), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n985), .B1(new_n979), .B2(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n978), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT47), .Z(new_n990));
  NAND3_X1  g565(.A1(new_n979), .A2(G1996), .A3(new_n757), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT110), .Z(new_n992));
  OAI21_X1  g567(.A(new_n982), .B1(G1996), .B2(new_n757), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n979), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n729), .A2(new_n732), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n729), .A2(new_n732), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n979), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n978), .A2(G1986), .A3(G290), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT48), .Z(new_n1000));
  AND2_X1   g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n994), .A2(new_n996), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(G2067), .B2(new_n772), .ZN(new_n1003));
  AOI211_X1 g578(.A(new_n990), .B(new_n1001), .C1(new_n979), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT123), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n821), .B1(new_n1005), .B2(KEYINPUT57), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(KEYINPUT57), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT124), .ZN(new_n1009));
  OR2_X1    g584(.A1(G164), .A2(G1384), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n1014));
  NOR4_X1   g589(.A1(G164), .A2(KEYINPUT112), .A3(new_n1011), .A4(new_n973), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n977), .B(new_n1012), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT56), .B(G2072), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(G164), .A2(G1384), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1022), .A2(new_n976), .A3(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1024), .A2(G1956), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1019), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1010), .A2(KEYINPUT50), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1023), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n977), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1348), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1010), .A2(new_n976), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1029), .A2(new_n1030), .B1(new_n980), .B2(new_n1031), .ZN(new_n1032));
  OAI22_X1  g607(.A1(new_n1009), .A2(new_n1026), .B1(new_n618), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1026), .A2(new_n1008), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n483), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT68), .B1(new_n479), .B2(G2105), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1038), .A2(new_n1020), .A3(G40), .A4(new_n475), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n1024), .A2(G1348), .B1(G2067), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT60), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT125), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT125), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1032), .A2(new_n1043), .A3(KEYINPUT60), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1044), .A3(new_n626), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT125), .B(new_n618), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1045), .B(new_n1046), .C1(KEYINPUT60), .C2(new_n1032), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT58), .B(G1341), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1016), .A2(G1996), .B1(new_n1031), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1049), .A2(new_n565), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1050), .A2(KEYINPUT59), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(KEYINPUT59), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1047), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1008), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1034), .B1(new_n1054), .B2(KEYINPUT61), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1026), .A2(new_n1056), .A3(new_n1008), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1035), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1016), .A2(new_n705), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1024), .A2(new_n797), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n584), .B2(new_n587), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT55), .B(G8), .C1(new_n584), .C2(new_n587), .ZN(new_n1067));
  NAND2_X1  g642(.A1(KEYINPUT117), .A2(G8), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1063), .A2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1016), .A2(new_n705), .B1(new_n1024), .B2(new_n797), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1072), .A2(new_n1069), .A3(new_n1060), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n698), .A2(G1976), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT113), .B(G8), .C1(new_n1010), .C2(new_n976), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT113), .B1(new_n1039), .B2(G8), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1075), .B(new_n1077), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n595), .A2(G651), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n598), .A2(new_n534), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n693), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT114), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n599), .A2(new_n1086), .A3(new_n693), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT49), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n599), .A2(new_n693), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1089), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1079), .A2(new_n1080), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1031), .B2(new_n1060), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1097), .A2(new_n1078), .B1(G1976), .B2(new_n698), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1081), .B(new_n1095), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1074), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1016), .B2(G2078), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1029), .A2(new_n749), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1020), .B2(KEYINPUT45), .ZN(new_n1107));
  NOR4_X1   g682(.A1(G164), .A2(KEYINPUT118), .A3(new_n1011), .A4(G1384), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n977), .B(new_n1012), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1103), .B(new_n1104), .C1(new_n1105), .C2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(G301), .B(KEYINPUT54), .Z(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n541), .A2(G8), .A3(new_n542), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT51), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G1966), .ZN(new_n1117));
  INV_X1    g692(.A(G2084), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1109), .A2(new_n1117), .B1(new_n1024), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(G8), .B(new_n1116), .C1(new_n1120), .C2(G286), .ZN(new_n1121));
  OAI221_X1 g696(.A(new_n1114), .B1(new_n1115), .B2(KEYINPUT51), .C1(new_n1119), .C2(new_n1060), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(G8), .A3(G286), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n973), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n499), .A2(new_n501), .ZN(new_n1126));
  OAI211_X1 g701(.A(KEYINPUT45), .B(new_n1125), .C1(new_n1126), .C2(new_n497), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT112), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n974), .A2(new_n1013), .A3(KEYINPUT45), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1130), .A2(G40), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n975), .A2(new_n1105), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n475), .A4(new_n480), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(new_n1103), .A3(new_n1104), .A4(new_n1111), .ZN(new_n1134));
  AND4_X1   g709(.A1(new_n1101), .A2(new_n1113), .A3(new_n1124), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1059), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1063), .A2(new_n1070), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1069), .B1(new_n1072), .B2(new_n1060), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1100), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n1110), .A4(G171), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1124), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT62), .A4(new_n1123), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g722(.A(KEYINPUT127), .B(new_n1141), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1136), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1109), .A2(new_n1117), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1029), .A2(G2084), .ZN(new_n1152));
  OAI211_X1 g727(.A(G8), .B(G168), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1100), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n976), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1156));
  AOI21_X1  g731(.A(G1971), .B1(new_n1130), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1029), .A2(G2090), .ZN(new_n1158));
  OAI211_X1 g733(.A(G8), .B(new_n1155), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1159), .A2(KEYINPUT63), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1155), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1072), .B2(new_n1060), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1154), .A2(KEYINPUT121), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1119), .A2(new_n1060), .A3(G286), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1075), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1097), .A2(new_n1078), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT49), .B1(new_n1168), .B2(new_n1090), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1092), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1166), .A2(KEYINPUT52), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1165), .A2(new_n1171), .A3(new_n1081), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1162), .A2(KEYINPUT63), .A3(new_n1159), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1164), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1163), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT119), .B1(new_n1074), .B2(new_n1172), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1154), .A2(new_n1177), .A3(new_n1139), .ZN(new_n1178));
  XNOR2_X1  g753(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(G288), .A2(G1976), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT116), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1168), .B1(new_n1095), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1167), .B(KEYINPUT115), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1187), .B1(new_n1100), .B2(new_n1159), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1150), .B1(new_n1181), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g765(.A(KEYINPUT122), .B(new_n1188), .C1(new_n1175), .C2(new_n1180), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1149), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  XOR2_X1   g767(.A(G290), .B(G1986), .Z(new_n1193));
  OAI21_X1  g768(.A(new_n998), .B1(new_n978), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1004), .B1(new_n1192), .B2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g770(.A(G227), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n661), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n1198), .B1(new_n873), .B2(new_n876), .ZN(new_n1199));
  INV_X1    g773(.A(G229), .ZN(new_n1200));
  NAND4_X1  g774(.A1(new_n1199), .A2(G319), .A3(new_n1200), .A4(new_n961), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


