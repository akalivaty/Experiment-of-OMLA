

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U557 ( .A1(n535), .A2(n534), .ZN(G164) );
  NOR2_X1 U558 ( .A1(n544), .A2(n543), .ZN(G160) );
  NOR2_X1 U559 ( .A1(n531), .A2(G2104), .ZN(n624) );
  NOR2_X2 U560 ( .A1(n798), .A2(n797), .ZN(n799) );
  BUF_X1 U561 ( .A(n624), .Z(n522) );
  NOR2_X1 U562 ( .A1(n724), .A2(n1016), .ZN(n733) );
  INV_X1 U563 ( .A(n1003), .ZN(n792) );
  NOR2_X2 U564 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  AND2_X1 U565 ( .A1(n805), .A2(n526), .ZN(n523) );
  AND2_X1 U566 ( .A1(n530), .A2(n529), .ZN(n524) );
  OR2_X1 U567 ( .A1(n803), .A2(n802), .ZN(n525) );
  AND2_X1 U568 ( .A1(n804), .A2(n525), .ZN(n526) );
  NAND2_X1 U569 ( .A1(n786), .A2(n785), .ZN(n527) );
  AND2_X1 U570 ( .A1(n720), .A2(n721), .ZN(n726) );
  INV_X1 U571 ( .A(KEYINPUT31), .ZN(n760) );
  OR2_X1 U572 ( .A1(n750), .A2(n749), .ZN(n763) );
  INV_X1 U573 ( .A(KEYINPUT95), .ZN(n764) );
  INV_X1 U574 ( .A(n1007), .ZN(n787) );
  NAND2_X1 U575 ( .A1(n721), .A2(n720), .ZN(n766) );
  NOR2_X1 U576 ( .A1(n793), .A2(n792), .ZN(n794) );
  INV_X1 U577 ( .A(G2105), .ZN(n531) );
  INV_X1 U578 ( .A(n532), .ZN(n891) );
  XOR2_X1 U579 ( .A(KEYINPUT72), .B(n602), .Z(n1011) );
  XOR2_X2 U580 ( .A(KEYINPUT17), .B(n528), .Z(n893) );
  NAND2_X1 U581 ( .A1(n893), .A2(G138), .ZN(n535) );
  NAND2_X1 U582 ( .A1(G126), .A2(n624), .ZN(n530) );
  AND2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U584 ( .A1(G114), .A2(n886), .ZN(n529) );
  AND2_X1 U585 ( .A1(n531), .A2(G2104), .ZN(n537) );
  INV_X1 U586 ( .A(n537), .ZN(n532) );
  NAND2_X1 U587 ( .A1(G102), .A2(n891), .ZN(n533) );
  AND2_X1 U588 ( .A1(n524), .A2(n533), .ZN(n534) );
  NAND2_X1 U589 ( .A1(G125), .A2(n624), .ZN(n536) );
  XNOR2_X1 U590 ( .A(n536), .B(KEYINPUT64), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G101), .A2(n537), .ZN(n538) );
  XOR2_X1 U592 ( .A(KEYINPUT23), .B(n538), .Z(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U594 ( .A1(G137), .A2(n893), .ZN(n542) );
  NAND2_X1 U595 ( .A1(G113), .A2(n886), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n542), .A2(n541), .ZN(n543) );
  INV_X1 U597 ( .A(G651), .ZN(n550) );
  NOR2_X1 U598 ( .A1(G543), .A2(n550), .ZN(n545) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n545), .Z(n591) );
  BUF_X1 U600 ( .A(n591), .Z(n661) );
  NAND2_X1 U601 ( .A1(G63), .A2(n661), .ZN(n547) );
  XOR2_X1 U602 ( .A(G543), .B(KEYINPUT0), .Z(n662) );
  NOR2_X1 U603 ( .A1(G651), .A2(n662), .ZN(n595) );
  BUF_X1 U604 ( .A(n595), .Z(n656) );
  NAND2_X1 U605 ( .A1(G51), .A2(n656), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U607 ( .A(KEYINPUT6), .B(n548), .ZN(n556) );
  NOR2_X2 U608 ( .A1(G543), .A2(G651), .ZN(n648) );
  NAND2_X1 U609 ( .A1(n648), .A2(G89), .ZN(n549) );
  XNOR2_X1 U610 ( .A(n549), .B(KEYINPUT4), .ZN(n552) );
  NOR2_X1 U611 ( .A1(n662), .A2(n550), .ZN(n592) );
  BUF_X1 U612 ( .A(n592), .Z(n645) );
  NAND2_X1 U613 ( .A1(G76), .A2(n645), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U615 ( .A(KEYINPUT5), .B(n553), .ZN(n554) );
  XNOR2_X1 U616 ( .A(KEYINPUT73), .B(n554), .ZN(n555) );
  NOR2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U618 ( .A(KEYINPUT7), .B(n557), .Z(G168) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U620 ( .A1(G60), .A2(n661), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G47), .A2(n656), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G72), .A2(n645), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G85), .A2(n648), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U626 ( .A1(n563), .A2(n562), .ZN(G290) );
  AND2_X1 U627 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  NAND2_X1 U631 ( .A1(G64), .A2(n661), .ZN(n565) );
  NAND2_X1 U632 ( .A1(G52), .A2(n656), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G77), .A2(n645), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G90), .A2(n648), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U637 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U638 ( .A1(n570), .A2(n569), .ZN(G171) );
  NAND2_X1 U639 ( .A1(G75), .A2(n645), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G88), .A2(n648), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G62), .A2(n661), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G50), .A2(n656), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U645 ( .A1(n576), .A2(n575), .ZN(G166) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n577) );
  XNOR2_X1 U647 ( .A(n577), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U648 ( .A(G223), .ZN(n826) );
  NAND2_X1 U649 ( .A1(n826), .A2(G567), .ZN(n578) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n578), .Z(G234) );
  NAND2_X1 U651 ( .A1(n656), .A2(G43), .ZN(n579) );
  XNOR2_X1 U652 ( .A(KEYINPUT70), .B(n579), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G56), .A2(n661), .ZN(n580) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n580), .Z(n588) );
  NAND2_X1 U655 ( .A1(n648), .A2(G81), .ZN(n581) );
  XNOR2_X1 U656 ( .A(KEYINPUT12), .B(n581), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n592), .A2(G68), .ZN(n582) );
  XNOR2_X1 U658 ( .A(n582), .B(KEYINPUT68), .ZN(n583) );
  AND2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U660 ( .A(KEYINPUT13), .B(n585), .Z(n586) );
  XNOR2_X1 U661 ( .A(n586), .B(KEYINPUT69), .ZN(n587) );
  NOR2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n1016) );
  INV_X1 U664 ( .A(G860), .ZN(n617) );
  OR2_X1 U665 ( .A1(n1016), .A2(n617), .ZN(G153) );
  INV_X1 U666 ( .A(G171), .ZN(G301) );
  NAND2_X1 U667 ( .A1(G92), .A2(n648), .ZN(n600) );
  NAND2_X1 U668 ( .A1(G66), .A2(n591), .ZN(n594) );
  NAND2_X1 U669 ( .A1(G79), .A2(n592), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U671 ( .A1(G54), .A2(n595), .ZN(n596) );
  XNOR2_X1 U672 ( .A(KEYINPUT71), .B(n596), .ZN(n597) );
  NOR2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT15), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n1011), .A2(G868), .ZN(n604) );
  INV_X1 U677 ( .A(G868), .ZN(n614) );
  NOR2_X1 U678 ( .A1(n614), .A2(G301), .ZN(n603) );
  NOR2_X1 U679 ( .A1(n604), .A2(n603), .ZN(G284) );
  NAND2_X1 U680 ( .A1(G65), .A2(n661), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT66), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G78), .A2(n645), .ZN(n606) );
  XOR2_X1 U683 ( .A(KEYINPUT65), .B(n606), .Z(n607) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G53), .A2(n656), .ZN(n609) );
  XNOR2_X1 U686 ( .A(KEYINPUT67), .B(n609), .ZN(n610) );
  NOR2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n648), .A2(G91), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G299) );
  NOR2_X1 U690 ( .A1(G286), .A2(n614), .ZN(n616) );
  NOR2_X1 U691 ( .A1(G868), .A2(G299), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n616), .A2(n615), .ZN(G297) );
  NAND2_X1 U693 ( .A1(n617), .A2(G559), .ZN(n618) );
  INV_X1 U694 ( .A(n1011), .ZN(n732) );
  NAND2_X1 U695 ( .A1(n618), .A2(n732), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n619), .B(KEYINPUT74), .ZN(n620) );
  XNOR2_X1 U697 ( .A(KEYINPUT16), .B(n620), .ZN(G148) );
  NOR2_X1 U698 ( .A1(G868), .A2(n1016), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n732), .A2(G868), .ZN(n621) );
  NOR2_X1 U700 ( .A1(G559), .A2(n621), .ZN(n622) );
  NOR2_X1 U701 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U702 ( .A1(n522), .A2(G123), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT18), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G135), .A2(n893), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT75), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G99), .A2(n891), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n886), .A2(G111), .ZN(n631) );
  XOR2_X1 U710 ( .A(KEYINPUT76), .B(n631), .Z(n632) );
  NOR2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n953) );
  XNOR2_X1 U712 ( .A(G2096), .B(n953), .ZN(n635) );
  INV_X1 U713 ( .A(G2100), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(G156) );
  NAND2_X1 U715 ( .A1(G67), .A2(n661), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G55), .A2(n656), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G80), .A2(n645), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G93), .A2(n648), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U721 ( .A1(n641), .A2(n640), .ZN(n673) );
  NAND2_X1 U722 ( .A1(n732), .A2(G559), .ZN(n642) );
  XOR2_X1 U723 ( .A(n1016), .B(n642), .Z(n671) );
  XNOR2_X1 U724 ( .A(KEYINPUT77), .B(n671), .ZN(n643) );
  NOR2_X1 U725 ( .A1(G860), .A2(n643), .ZN(n644) );
  XNOR2_X1 U726 ( .A(n673), .B(n644), .ZN(G145) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(KEYINPUT79), .Z(n647) );
  NAND2_X1 U728 ( .A1(G73), .A2(n645), .ZN(n646) );
  XNOR2_X1 U729 ( .A(n647), .B(n646), .ZN(n655) );
  NAND2_X1 U730 ( .A1(G61), .A2(n661), .ZN(n650) );
  NAND2_X1 U731 ( .A1(G86), .A2(n648), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n656), .A2(G48), .ZN(n651) );
  XOR2_X1 U734 ( .A(KEYINPUT80), .B(n651), .Z(n652) );
  NOR2_X1 U735 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n655), .A2(n654), .ZN(G305) );
  NAND2_X1 U737 ( .A1(G49), .A2(n656), .ZN(n658) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n657) );
  NAND2_X1 U739 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U740 ( .A(KEYINPUT78), .B(n659), .ZN(n660) );
  NOR2_X1 U741 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n662), .A2(G87), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n664), .A2(n663), .ZN(G288) );
  INV_X1 U744 ( .A(G299), .ZN(n1006) );
  XNOR2_X1 U745 ( .A(n1006), .B(G305), .ZN(n665) );
  XNOR2_X1 U746 ( .A(n665), .B(G288), .ZN(n668) );
  XOR2_X1 U747 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n666) );
  XNOR2_X1 U748 ( .A(G290), .B(n666), .ZN(n667) );
  XOR2_X1 U749 ( .A(n668), .B(n667), .Z(n670) );
  XNOR2_X1 U750 ( .A(G166), .B(n673), .ZN(n669) );
  XNOR2_X1 U751 ( .A(n670), .B(n669), .ZN(n852) );
  XNOR2_X1 U752 ( .A(n671), .B(n852), .ZN(n672) );
  NAND2_X1 U753 ( .A1(n672), .A2(G868), .ZN(n675) );
  OR2_X1 U754 ( .A1(G868), .A2(n673), .ZN(n674) );
  NAND2_X1 U755 ( .A1(n675), .A2(n674), .ZN(G295) );
  XOR2_X1 U756 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n677) );
  NAND2_X1 U757 ( .A1(G2084), .A2(G2078), .ZN(n676) );
  XNOR2_X1 U758 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U761 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n681) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n681), .Z(n682) );
  NOR2_X1 U765 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U766 ( .A1(G96), .A2(n683), .ZN(n831) );
  NAND2_X1 U767 ( .A1(G2106), .A2(n831), .ZN(n687) );
  NAND2_X1 U768 ( .A1(G69), .A2(G120), .ZN(n684) );
  NOR2_X1 U769 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G108), .A2(n685), .ZN(n830) );
  NAND2_X1 U771 ( .A1(G567), .A2(n830), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n687), .A2(n686), .ZN(n833) );
  NAND2_X1 U773 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U774 ( .A1(n833), .A2(n688), .ZN(n829) );
  NAND2_X1 U775 ( .A1(n829), .A2(G36), .ZN(G176) );
  INV_X1 U776 ( .A(G166), .ZN(G303) );
  NOR2_X2 U777 ( .A1(G164), .A2(G1384), .ZN(n720) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n718) );
  NOR2_X1 U779 ( .A1(n720), .A2(n718), .ZN(n820) );
  NAND2_X1 U780 ( .A1(n893), .A2(G140), .ZN(n689) );
  XNOR2_X1 U781 ( .A(n689), .B(KEYINPUT84), .ZN(n691) );
  NAND2_X1 U782 ( .A1(G104), .A2(n891), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U784 ( .A(KEYINPUT34), .B(n692), .ZN(n697) );
  NAND2_X1 U785 ( .A1(G128), .A2(n522), .ZN(n694) );
  NAND2_X1 U786 ( .A1(G116), .A2(n886), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U788 ( .A(KEYINPUT35), .B(n695), .Z(n696) );
  NOR2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U790 ( .A(KEYINPUT36), .B(n698), .ZN(n903) );
  XNOR2_X1 U791 ( .A(G2067), .B(KEYINPUT37), .ZN(n818) );
  NOR2_X1 U792 ( .A1(n903), .A2(n818), .ZN(n970) );
  NAND2_X1 U793 ( .A1(n820), .A2(n970), .ZN(n816) );
  XOR2_X1 U794 ( .A(KEYINPUT86), .B(G1991), .Z(n923) );
  NAND2_X1 U795 ( .A1(n522), .A2(G119), .ZN(n701) );
  NAND2_X1 U796 ( .A1(G95), .A2(n891), .ZN(n699) );
  XOR2_X1 U797 ( .A(KEYINPUT85), .B(n699), .Z(n700) );
  NAND2_X1 U798 ( .A1(n701), .A2(n700), .ZN(n705) );
  NAND2_X1 U799 ( .A1(G131), .A2(n893), .ZN(n703) );
  NAND2_X1 U800 ( .A1(G107), .A2(n886), .ZN(n702) );
  NAND2_X1 U801 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n877) );
  NOR2_X1 U803 ( .A1(n923), .A2(n877), .ZN(n715) );
  NAND2_X1 U804 ( .A1(G105), .A2(n891), .ZN(n706) );
  XNOR2_X1 U805 ( .A(n706), .B(KEYINPUT38), .ZN(n713) );
  NAND2_X1 U806 ( .A1(G141), .A2(n893), .ZN(n708) );
  NAND2_X1 U807 ( .A1(G129), .A2(n522), .ZN(n707) );
  NAND2_X1 U808 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U809 ( .A1(G117), .A2(n886), .ZN(n709) );
  XNOR2_X1 U810 ( .A(KEYINPUT87), .B(n709), .ZN(n710) );
  NOR2_X1 U811 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U812 ( .A1(n713), .A2(n712), .ZN(n880) );
  AND2_X1 U813 ( .A1(n880), .A2(G1996), .ZN(n714) );
  NOR2_X1 U814 ( .A1(n715), .A2(n714), .ZN(n956) );
  INV_X1 U815 ( .A(n820), .ZN(n716) );
  NOR2_X1 U816 ( .A1(n956), .A2(n716), .ZN(n813) );
  INV_X1 U817 ( .A(n813), .ZN(n717) );
  NAND2_X1 U818 ( .A1(n816), .A2(n717), .ZN(n807) );
  NOR2_X1 U819 ( .A1(G1976), .A2(G288), .ZN(n1013) );
  INV_X1 U820 ( .A(n718), .ZN(n721) );
  AND2_X1 U821 ( .A1(n726), .A2(G1996), .ZN(n719) );
  XOR2_X1 U822 ( .A(n719), .B(KEYINPUT26), .Z(n723) );
  NAND2_X1 U823 ( .A1(n766), .A2(G1341), .ZN(n722) );
  NAND2_X1 U824 ( .A1(n723), .A2(n722), .ZN(n724) );
  OR2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n731) );
  NAND2_X1 U826 ( .A1(G1348), .A2(n766), .ZN(n725) );
  XNOR2_X1 U827 ( .A(KEYINPUT91), .B(n725), .ZN(n729) );
  NAND2_X1 U828 ( .A1(G2067), .A2(n726), .ZN(n727) );
  XOR2_X1 U829 ( .A(KEYINPUT92), .B(n727), .Z(n728) );
  NOR2_X1 U830 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U831 ( .A1(n731), .A2(n730), .ZN(n740) );
  NAND2_X1 U832 ( .A1(n733), .A2(n732), .ZN(n738) );
  NAND2_X1 U833 ( .A1(n726), .A2(G2072), .ZN(n734) );
  XNOR2_X1 U834 ( .A(n734), .B(KEYINPUT27), .ZN(n736) );
  INV_X1 U835 ( .A(G1956), .ZN(n982) );
  NOR2_X1 U836 ( .A1(n982), .A2(n726), .ZN(n735) );
  NOR2_X1 U837 ( .A1(n736), .A2(n735), .ZN(n741) );
  NAND2_X1 U838 ( .A1(n741), .A2(n1006), .ZN(n737) );
  AND2_X1 U839 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U840 ( .A1(n740), .A2(n739), .ZN(n745) );
  NOR2_X1 U841 ( .A1(n741), .A2(n1006), .ZN(n743) );
  XOR2_X1 U842 ( .A(KEYINPUT90), .B(KEYINPUT28), .Z(n742) );
  XNOR2_X1 U843 ( .A(n743), .B(n742), .ZN(n744) );
  NAND2_X1 U844 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U845 ( .A(n746), .B(KEYINPUT29), .ZN(n750) );
  XOR2_X1 U846 ( .A(G2078), .B(KEYINPUT25), .Z(n924) );
  NOR2_X1 U847 ( .A1(n924), .A2(n766), .ZN(n748) );
  NOR2_X1 U848 ( .A1(n726), .A2(G1961), .ZN(n747) );
  NOR2_X1 U849 ( .A1(n748), .A2(n747), .ZN(n757) );
  NOR2_X1 U850 ( .A1(G301), .A2(n757), .ZN(n749) );
  NAND2_X1 U851 ( .A1(G8), .A2(n766), .ZN(n803) );
  NOR2_X1 U852 ( .A1(G1966), .A2(n803), .ZN(n776) );
  NOR2_X1 U853 ( .A1(n766), .A2(G2084), .ZN(n751) );
  XNOR2_X1 U854 ( .A(n751), .B(KEYINPUT88), .ZN(n778) );
  NOR2_X1 U855 ( .A1(n776), .A2(n778), .ZN(n753) );
  INV_X1 U856 ( .A(KEYINPUT93), .ZN(n752) );
  XNOR2_X1 U857 ( .A(n753), .B(n752), .ZN(n754) );
  NAND2_X1 U858 ( .A1(n754), .A2(G8), .ZN(n755) );
  XNOR2_X1 U859 ( .A(n755), .B(KEYINPUT30), .ZN(n756) );
  NOR2_X1 U860 ( .A1(n756), .A2(G168), .ZN(n759) );
  AND2_X1 U861 ( .A1(G301), .A2(n757), .ZN(n758) );
  NOR2_X1 U862 ( .A1(n759), .A2(n758), .ZN(n761) );
  XNOR2_X1 U863 ( .A(n761), .B(n760), .ZN(n762) );
  NAND2_X1 U864 ( .A1(n763), .A2(n762), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n774), .A2(G286), .ZN(n765) );
  XNOR2_X1 U866 ( .A(n765), .B(n764), .ZN(n771) );
  NOR2_X1 U867 ( .A1(G1971), .A2(n803), .ZN(n768) );
  NOR2_X1 U868 ( .A1(G2090), .A2(n766), .ZN(n767) );
  NOR2_X1 U869 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U870 ( .A1(G303), .A2(n769), .ZN(n770) );
  NAND2_X1 U871 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U872 ( .A1(n772), .A2(G8), .ZN(n773) );
  XNOR2_X1 U873 ( .A(n773), .B(KEYINPUT32), .ZN(n783) );
  INV_X1 U874 ( .A(n774), .ZN(n775) );
  NOR2_X1 U875 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U876 ( .A(KEYINPUT94), .B(n777), .Z(n781) );
  NAND2_X1 U877 ( .A1(G8), .A2(n778), .ZN(n779) );
  XNOR2_X1 U878 ( .A(KEYINPUT89), .B(n779), .ZN(n780) );
  OR2_X1 U879 ( .A1(n781), .A2(n780), .ZN(n782) );
  AND2_X2 U880 ( .A1(n783), .A2(n782), .ZN(n798) );
  NOR2_X1 U881 ( .A1(n1013), .A2(n798), .ZN(n786) );
  NOR2_X1 U882 ( .A1(G1971), .A2(G303), .ZN(n784) );
  XOR2_X1 U883 ( .A(n784), .B(KEYINPUT96), .Z(n785) );
  NAND2_X1 U884 ( .A1(G1976), .A2(G288), .ZN(n1007) );
  NOR2_X1 U885 ( .A1(n803), .A2(n787), .ZN(n788) );
  NAND2_X1 U886 ( .A1(n527), .A2(n788), .ZN(n790) );
  INV_X1 U887 ( .A(KEYINPUT33), .ZN(n789) );
  NAND2_X1 U888 ( .A1(n790), .A2(n789), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n1013), .A2(KEYINPUT33), .ZN(n791) );
  NOR2_X1 U890 ( .A1(n791), .A2(n803), .ZN(n793) );
  XOR2_X1 U891 ( .A(G1981), .B(G305), .Z(n1003) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G166), .A2(G8), .ZN(n796) );
  NOR2_X1 U894 ( .A1(G2090), .A2(n796), .ZN(n797) );
  XNOR2_X1 U895 ( .A(n799), .B(KEYINPUT97), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n800), .A2(n803), .ZN(n804) );
  NOR2_X1 U897 ( .A1(G1981), .A2(G305), .ZN(n801) );
  XOR2_X1 U898 ( .A(n801), .B(KEYINPUT24), .Z(n802) );
  XNOR2_X1 U899 ( .A(KEYINPUT98), .B(n523), .ZN(n806) );
  NOR2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n810) );
  XOR2_X1 U901 ( .A(G1986), .B(KEYINPUT83), .Z(n808) );
  XNOR2_X1 U902 ( .A(G290), .B(n808), .ZN(n1010) );
  NAND2_X1 U903 ( .A1(n1010), .A2(n820), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n823) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n880), .ZN(n963) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n811) );
  AND2_X1 U907 ( .A1(n923), .A2(n877), .ZN(n952) );
  NOR2_X1 U908 ( .A1(n811), .A2(n952), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n963), .A2(n814), .ZN(n815) );
  XNOR2_X1 U911 ( .A(n815), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n903), .A2(n818), .ZN(n967) );
  NAND2_X1 U914 ( .A1(n819), .A2(n967), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n825) );
  XOR2_X1 U917 ( .A(KEYINPUT40), .B(KEYINPUT99), .Z(n824) );
  XNOR2_X1 U918 ( .A(n825), .B(n824), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U921 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  NOR2_X1 U928 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n832), .B(KEYINPUT101), .ZN(G261) );
  INV_X1 U930 ( .A(G261), .ZN(G325) );
  XOR2_X1 U931 ( .A(KEYINPUT102), .B(n833), .Z(G319) );
  XOR2_X1 U932 ( .A(KEYINPUT42), .B(G2072), .Z(n835) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2078), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U935 ( .A(n836), .B(G2096), .Z(n838) );
  XNOR2_X1 U936 ( .A(G2084), .B(G2090), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U938 ( .A(KEYINPUT43), .B(KEYINPUT103), .Z(n840) );
  XNOR2_X1 U939 ( .A(G2678), .B(G2100), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n842), .B(n841), .Z(G227) );
  XOR2_X1 U942 ( .A(G1976), .B(G1981), .Z(n844) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1961), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U945 ( .A(n845), .B(G2474), .Z(n847) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1971), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U948 ( .A(KEYINPUT41), .B(G1956), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G229) );
  XNOR2_X1 U952 ( .A(n1016), .B(n852), .ZN(n854) );
  XNOR2_X1 U953 ( .A(G171), .B(n1011), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U955 ( .A(G286), .B(n855), .Z(n856) );
  NOR2_X1 U956 ( .A1(G37), .A2(n856), .ZN(n857) );
  XOR2_X1 U957 ( .A(KEYINPUT115), .B(n857), .Z(G397) );
  NAND2_X1 U958 ( .A1(G100), .A2(n891), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G112), .A2(n886), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U961 ( .A(KEYINPUT106), .B(n860), .ZN(n867) );
  NAND2_X1 U962 ( .A1(n522), .A2(G124), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT44), .B(n861), .Z(n864) );
  NAND2_X1 U964 ( .A1(n893), .A2(G136), .ZN(n862) );
  XOR2_X1 U965 ( .A(KEYINPUT104), .B(n862), .Z(n863) );
  NOR2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n865), .B(KEYINPUT105), .ZN(n866) );
  NOR2_X1 U968 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U969 ( .A1(G139), .A2(n893), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G103), .A2(n891), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G127), .A2(n522), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G115), .A2(n886), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  XNOR2_X1 U976 ( .A(KEYINPUT110), .B(n873), .ZN(n874) );
  NOR2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U978 ( .A(KEYINPUT111), .B(n876), .Z(n946) );
  XNOR2_X1 U979 ( .A(n877), .B(n946), .ZN(n885) );
  XOR2_X1 U980 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n879) );
  XNOR2_X1 U981 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n878) );
  XNOR2_X1 U982 ( .A(n879), .B(n878), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n881), .B(n880), .ZN(n883) );
  XNOR2_X1 U984 ( .A(G164), .B(G160), .ZN(n882) );
  XNOR2_X1 U985 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n900) );
  NAND2_X1 U987 ( .A1(G118), .A2(n886), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n887), .B(KEYINPUT108), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G130), .A2(n522), .ZN(n888) );
  XOR2_X1 U990 ( .A(KEYINPUT107), .B(n888), .Z(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n898) );
  NAND2_X1 U992 ( .A1(n891), .A2(G106), .ZN(n892) );
  XOR2_X1 U993 ( .A(KEYINPUT109), .B(n892), .Z(n895) );
  NAND2_X1 U994 ( .A1(n893), .A2(G142), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U996 ( .A(KEYINPUT45), .B(n896), .Z(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U999 ( .A(G162), .B(n953), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n905), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(KEYINPUT114), .B(n906), .ZN(G395) );
  XOR2_X1 U1004 ( .A(G2443), .B(G2451), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G2446), .B(G2454), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1007 ( .A(n909), .B(G2427), .Z(n911) );
  XNOR2_X1 U1008 ( .A(G1348), .B(G1341), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1010 ( .A(G2435), .B(KEYINPUT100), .Z(n913) );
  XNOR2_X1 U1011 ( .A(G2430), .B(G2438), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1013 ( .A(n915), .B(n914), .Z(n916) );
  NAND2_X1 U1014 ( .A1(G14), .A2(n916), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(n922), .A2(G319), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(G397), .A2(G395), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  INV_X1 U1023 ( .A(n922), .ZN(G401) );
  XOR2_X1 U1024 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n936) );
  XOR2_X1 U1025 ( .A(n923), .B(G25), .Z(n926) );
  XNOR2_X1 U1026 ( .A(G27), .B(n924), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(G1996), .B(G32), .ZN(n928) );
  XNOR2_X1 U1029 ( .A(G33), .B(G2072), .ZN(n927) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1031 ( .A1(G28), .A2(n929), .ZN(n932) );
  XOR2_X1 U1032 ( .A(KEYINPUT121), .B(G2067), .Z(n930) );
  XNOR2_X1 U1033 ( .A(G26), .B(n930), .ZN(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(n936), .B(n935), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(G2090), .B(KEYINPUT120), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(G35), .B(n937), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n942) );
  XOR2_X1 U1040 ( .A(G2084), .B(G34), .Z(n940) );
  XNOR2_X1 U1041 ( .A(KEYINPUT54), .B(n940), .ZN(n941) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(G29), .A2(KEYINPUT55), .ZN(n943) );
  NAND2_X1 U1044 ( .A1(n945), .A2(n943), .ZN(n944) );
  NAND2_X1 U1045 ( .A1(G11), .A2(n944), .ZN(n978) );
  INV_X1 U1046 ( .A(KEYINPUT55), .ZN(n972) );
  OR2_X1 U1047 ( .A1(n972), .A2(n945), .ZN(n976) );
  XNOR2_X1 U1048 ( .A(G2072), .B(n946), .ZN(n949) );
  XNOR2_X1 U1049 ( .A(G164), .B(G2078), .ZN(n947) );
  XNOR2_X1 U1050 ( .A(n947), .B(KEYINPUT118), .ZN(n948) );
  NAND2_X1 U1051 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1052 ( .A(n950), .B(KEYINPUT50), .ZN(n951) );
  XNOR2_X1 U1053 ( .A(KEYINPUT119), .B(n951), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1055 ( .A(KEYINPUT117), .B(n954), .Z(n955) );
  NAND2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1057 ( .A(G2084), .B(G160), .Z(n957) );
  XNOR2_X1 U1058 ( .A(KEYINPUT116), .B(n957), .ZN(n958) );
  NOR2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n966) );
  XOR2_X1 U1061 ( .A(G2090), .B(G162), .Z(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1063 ( .A(n964), .B(KEYINPUT51), .ZN(n965) );
  NOR2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(KEYINPUT52), .B(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(G29), .A2(n974), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n1033) );
  XNOR2_X1 U1072 ( .A(G1341), .B(G19), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G1981), .B(G6), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(KEYINPUT126), .B(n981), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(n982), .B(G20), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1078 ( .A(KEYINPUT59), .B(G1348), .Z(n985) );
  XNOR2_X1 U1079 ( .A(G4), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(KEYINPUT60), .B(n988), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(G1966), .B(G21), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(G5), .B(G1961), .ZN(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G1971), .B(G22), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(G23), .B(G1976), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n996) );
  XOR2_X1 U1089 ( .A(G1986), .B(G24), .Z(n995) );
  NAND2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1091 ( .A(KEYINPUT58), .B(n997), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1093 ( .A(KEYINPUT61), .B(n1000), .Z(n1001) );
  NOR2_X1 U1094 ( .A1(G16), .A2(n1001), .ZN(n1030) );
  XNOR2_X1 U1095 ( .A(G16), .B(KEYINPUT123), .ZN(n1002) );
  XNOR2_X1 U1096 ( .A(n1002), .B(KEYINPUT56), .ZN(n1028) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G168), .ZN(n1004) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1099 ( .A(KEYINPUT57), .B(n1005), .Z(n1025) );
  XNOR2_X1 U1100 ( .A(n1006), .B(G1956), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1022) );
  XNOR2_X1 U1102 ( .A(G1961), .B(G301), .ZN(n1009) );
  NOR2_X1 U1103 ( .A1(n1010), .A2(n1009), .ZN(n1020) );
  XNOR2_X1 U1104 ( .A(G166), .B(G1971), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1011), .B(G1348), .ZN(n1012) );
  NOR2_X1 U1106 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(G1341), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1112 ( .A(KEYINPUT124), .B(n1023), .Z(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1114 ( .A(KEYINPUT125), .B(n1026), .Z(n1027) );
  NOR2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1117 ( .A(KEYINPUT127), .B(n1031), .Z(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1034), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

