//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT28), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n208), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT28), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n202), .A2(new_n210), .A3(new_n203), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n205), .A2(new_n207), .A3(new_n209), .A4(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(new_n203), .ZN(new_n215));
  NAND3_X1  g014(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT23), .B1(new_n208), .B2(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n220), .B(new_n221), .C1(G169gat), .C2(G176gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT25), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n218), .A2(new_n222), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n227), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n215), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n225), .A2(new_n229), .A3(new_n230), .A4(new_n219), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n224), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT70), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n212), .A2(new_n224), .A3(new_n231), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G226gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n237), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT71), .ZN(new_n243));
  XNOR2_X1  g042(.A(G197gat), .B(G204gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT22), .ZN(new_n245));
  NAND2_X1  g044(.A1(G211gat), .A2(G218gat), .ZN(new_n246));
  INV_X1    g045(.A(G211gat), .ZN(new_n247));
  INV_X1    g046(.A(G218gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT22), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n246), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n244), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n256), .A3(new_n237), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n239), .A2(new_n243), .A3(new_n255), .A4(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n232), .A2(new_n237), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n238), .A2(KEYINPUT29), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(new_n236), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n254), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT72), .B(G64gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(G92gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(G8gat), .B(G36gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  NAND4_X1  g065(.A1(new_n258), .A2(new_n262), .A3(KEYINPUT30), .A4(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT73), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n258), .A2(new_n262), .A3(new_n266), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n258), .A2(new_n262), .ZN(new_n273));
  INV_X1    g072(.A(new_n266), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280));
  XOR2_X1   g079(.A(G113gat), .B(G120gat), .Z(new_n281));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G127gat), .B(G134gat), .Z(new_n286));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(KEYINPUT1), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT66), .ZN(new_n289));
  OR2_X1    g088(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n290));
  NAND2_X1  g089(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n285), .A2(new_n289), .B1(new_n280), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G141gat), .B(G148gat), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT74), .ZN(new_n295));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  INV_X1    g095(.A(G155gat), .ZN(new_n297));
  INV_X1    g096(.A(G162gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n296), .B1(new_n299), .B2(KEYINPUT2), .ZN(new_n300));
  XNOR2_X1  g099(.A(G141gat), .B(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n295), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n296), .B(new_n299), .C1(new_n301), .C2(KEYINPUT2), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n293), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT4), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n279), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n280), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n283), .A2(new_n284), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n288), .A2(KEYINPUT66), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n306), .A2(KEYINPUT3), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT3), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n304), .A2(new_n316), .A3(new_n305), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n306), .A2(KEYINPUT75), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n320), .A3(new_n305), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n293), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n310), .B(new_n318), .C1(new_n323), .C2(new_n309), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n314), .A2(new_n306), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n308), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n279), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(KEYINPUT5), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n293), .A2(new_n307), .A3(KEYINPUT4), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n279), .A2(KEYINPUT5), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n304), .A2(new_n316), .A3(new_n305), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n316), .B1(new_n304), .B2(new_n305), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n309), .B1(new_n333), .B2(new_n314), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n314), .B1(new_n319), .B2(new_n321), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n329), .B(new_n330), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT76), .ZN(new_n337));
  INV_X1    g136(.A(new_n329), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n318), .A2(KEYINPUT4), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(new_n323), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n330), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n328), .A2(new_n337), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344));
  INV_X1    g143(.A(G85gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT0), .B(G57gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n346), .B(new_n347), .Z(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT6), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n352));
  INV_X1    g151(.A(new_n348), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n328), .A2(new_n337), .A3(new_n342), .A4(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n349), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n277), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G78gat), .B(G106gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT31), .B(G50gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(G22gat), .ZN(new_n361));
  INV_X1    g160(.A(G22gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(KEYINPUT79), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n254), .B1(new_n331), .B2(KEYINPUT29), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n250), .B(KEYINPUT78), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n253), .B(KEYINPUT77), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT3), .B1(new_n369), .B2(new_n240), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n366), .B1(new_n370), .B2(new_n322), .ZN(new_n371));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n316), .B1(new_n254), .B2(KEYINPUT29), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n306), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n375), .A2(new_n366), .A3(G228gat), .A4(G233gat), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n365), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n373), .A2(new_n376), .A3(new_n365), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n293), .A2(new_n224), .A3(new_n212), .A4(new_n231), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n314), .A2(new_n232), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G227gat), .A2(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT32), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G15gat), .B(G43gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT68), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n381), .A2(new_n384), .A3(new_n382), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT69), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI22_X1  g196(.A1(new_n385), .A2(KEYINPUT69), .B1(KEYINPUT68), .B2(KEYINPUT34), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n397), .A2(KEYINPUT34), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n392), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n386), .B(KEYINPUT32), .C1(new_n388), .C2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n393), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n399), .B1(new_n393), .B2(new_n401), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n380), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT35), .B1(new_n357), .B2(new_n405), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n277), .A2(new_n405), .A3(KEYINPUT35), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n355), .A2(KEYINPUT84), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n349), .A2(new_n409), .A3(new_n352), .A4(new_n354), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n351), .A3(new_n410), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n407), .A2(KEYINPUT87), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT87), .B1(new_n407), .B2(new_n411), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n406), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n408), .A2(new_n351), .A3(new_n410), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT37), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n261), .B2(new_n255), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n239), .A2(new_n243), .A3(new_n257), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n255), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT38), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n422), .B(new_n274), .C1(new_n273), .C2(KEYINPUT37), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT86), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n419), .B(KEYINPUT85), .ZN(new_n425));
  INV_X1    g224(.A(new_n273), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n266), .B1(new_n426), .B2(new_n416), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT86), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n425), .A2(new_n427), .A3(new_n428), .A4(new_n422), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n427), .B1(new_n416), .B2(new_n426), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n431), .A2(KEYINPUT38), .B1(new_n426), .B2(new_n266), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n325), .A2(new_n308), .A3(new_n278), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(KEYINPUT39), .C1(new_n340), .C2(new_n278), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT81), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT39), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n318), .A2(KEYINPUT4), .B1(new_n322), .B2(new_n293), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n438), .B(new_n279), .C1(new_n439), .C2(new_n338), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n437), .B1(new_n440), .B2(new_n353), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n437), .A3(new_n353), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n436), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT82), .B1(new_n444), .B2(KEYINPUT40), .ZN(new_n445));
  INV_X1    g244(.A(new_n443), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n435), .B1(new_n446), .B2(new_n441), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT82), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT40), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(KEYINPUT40), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n350), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n444), .A2(KEYINPUT83), .A3(KEYINPUT40), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n451), .A2(new_n454), .A3(new_n277), .A4(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n433), .A2(new_n380), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n277), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n351), .A2(new_n355), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n380), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n404), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT36), .B1(new_n461), .B2(new_n402), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n403), .A2(new_n404), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT80), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n465), .B(new_n468), .C1(new_n356), .C2(new_n380), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n414), .B1(new_n457), .B2(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(G169gat), .B(G197gat), .Z(new_n472));
  XNOR2_X1  g271(.A(G113gat), .B(G141gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n476), .B(KEYINPUT12), .Z(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT16), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(G1gat), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(G1gat), .B2(new_n478), .ZN(new_n481));
  INV_X1    g280(.A(G8gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G50gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G43gat), .ZN(new_n485));
  INV_X1    g284(.A(G43gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G50gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n487), .A3(KEYINPUT15), .ZN(new_n488));
  INV_X1    g287(.A(G29gat), .ZN(new_n489));
  INV_X1    g288(.A(G36gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n493), .B2(KEYINPUT89), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT14), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(new_n489), .A3(new_n490), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n492), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n488), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G43gat), .B(G50gat), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n501), .A2(KEYINPUT15), .B1(new_n496), .B2(new_n492), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n491), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT90), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT90), .B1(new_n502), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT91), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511));
  OAI22_X1  g310(.A1(new_n501), .A2(KEYINPUT15), .B1(new_n489), .B2(new_n490), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n492), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n488), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n511), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT90), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT91), .A3(new_n500), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n483), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n510), .A2(new_n520), .A3(new_n518), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n508), .A2(KEYINPUT17), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n519), .B1(new_n523), .B2(new_n483), .ZN(new_n524));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT18), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n483), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(new_n521), .B2(new_n522), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n529));
  INV_X1    g328(.A(new_n525), .ZN(new_n530));
  NOR4_X1   g329(.A1(new_n528), .A2(new_n529), .A3(new_n519), .A4(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT91), .B1(new_n517), .B2(new_n500), .ZN(new_n533));
  AOI211_X1 g332(.A(new_n509), .B(new_n499), .C1(new_n515), .C2(new_n516), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n483), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n510), .A2(new_n518), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n527), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n525), .B(KEYINPUT13), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n477), .B1(new_n532), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n522), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n535), .B2(new_n520), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n538), .B(new_n525), .C1(new_n545), .C2(new_n527), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n529), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n524), .A2(KEYINPUT18), .A3(new_n525), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n542), .A4(new_n477), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT92), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(new_n542), .A3(new_n548), .ZN(new_n552));
  INV_X1    g351(.A(new_n477), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n549), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n471), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT99), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(G85gat), .A3(G92gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n563), .B1(new_n345), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n559), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G99gat), .B(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n562), .A2(new_n565), .A3(new_n568), .A4(new_n566), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n570), .A2(KEYINPUT100), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT100), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT17), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(new_n544), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n574), .B1(new_n533), .B2(new_n534), .ZN(new_n578));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT97), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n203), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n574), .B1(new_n521), .B2(new_n522), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n578), .A2(new_n582), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n585), .A2(new_n586), .A3(G190gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n248), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n577), .A2(new_n203), .A3(new_n583), .ZN(new_n589));
  OAI21_X1  g388(.A(G190gat), .B1(new_n585), .B2(new_n586), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(new_n590), .A3(G218gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(KEYINPUT98), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G134gat), .B(G162gat), .Z(new_n595));
  INV_X1    g394(.A(new_n593), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n588), .A2(KEYINPUT98), .A3(new_n596), .A4(new_n591), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n595), .B1(new_n594), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT93), .ZN(new_n601));
  XNOR2_X1  g400(.A(G57gat), .B(G64gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT9), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G71gat), .B(G78gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(KEYINPUT94), .ZN(new_n607));
  INV_X1    g406(.A(G71gat), .ZN(new_n608));
  INV_X1    g407(.A(G78gat), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n603), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(G64gat), .ZN(new_n611));
  OR3_X1    g410(.A1(new_n611), .A2(KEYINPUT94), .A3(G57gat), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n607), .A2(new_n605), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n605), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n614), .B(KEYINPUT93), .C1(new_n603), .C2(new_n602), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n606), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(KEYINPUT21), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT20), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(new_n247), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n483), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(G183gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n214), .A3(new_n483), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n623), .B2(new_n625), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n628), .B1(new_n632), .B2(new_n626), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n620), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n629), .B1(new_n627), .B2(new_n630), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n632), .A2(new_n628), .A3(new_n626), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n639), .A3(new_n619), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n634), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n637), .B1(new_n634), .B2(new_n640), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n606), .A2(new_n613), .A3(new_n615), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n570), .A2(new_n571), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n574), .A2(KEYINPUT10), .A3(new_n616), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n645), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n655), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n600), .A2(new_n643), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n558), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n459), .B(KEYINPUT102), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g467(.A1(new_n558), .A2(new_n277), .A3(new_n663), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  AND3_X1   g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n670), .B2(new_n672), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n670), .A2(KEYINPUT103), .A3(new_n482), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n669), .B2(G8gat), .ZN(new_n677));
  OAI22_X1  g476(.A1(new_n673), .A2(new_n674), .B1(new_n675), .B2(new_n677), .ZN(G1325gat));
  INV_X1    g477(.A(G15gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n461), .A2(new_n402), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n664), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT104), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT104), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n466), .A2(G15gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT105), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n683), .A2(new_n684), .B1(new_n665), .B2(new_n686), .ZN(G1326gat));
  NOR2_X1   g486(.A1(new_n664), .A2(new_n380), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT43), .B(G22gat), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NOR3_X1   g489(.A1(new_n600), .A2(new_n643), .A3(new_n660), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n558), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n489), .A3(new_n666), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT45), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n693), .A2(new_n696), .A3(new_n489), .A4(new_n666), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT87), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT35), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n458), .A2(new_n701), .A3(new_n680), .A4(new_n380), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n702), .B2(new_n415), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n407), .A2(KEYINPUT87), .A3(new_n411), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n433), .A2(new_n380), .A3(new_n456), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n460), .A2(new_n466), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n406), .A2(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n699), .B1(new_n708), .B2(new_n600), .ZN(new_n709));
  INV_X1    g508(.A(new_n600), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n471), .A2(KEYINPUT44), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n554), .A2(new_n549), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n643), .A2(new_n660), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n709), .A2(new_n711), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715));
  INV_X1    g514(.A(new_n666), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n714), .B2(new_n716), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(G29gat), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n698), .A2(new_n719), .ZN(G1328gat));
  NAND4_X1  g519(.A1(new_n558), .A2(new_n490), .A3(new_n277), .A4(new_n691), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n721), .A2(KEYINPUT107), .A3(KEYINPUT46), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT107), .B1(new_n721), .B2(KEYINPUT46), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n721), .A2(KEYINPUT46), .ZN(new_n725));
  OAI21_X1  g524(.A(G36gat), .B1(new_n714), .B2(new_n458), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(G1329gat));
  OAI21_X1  g526(.A(G43gat), .B1(new_n714), .B2(new_n465), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n558), .A2(new_n486), .A3(new_n680), .A4(new_n691), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT47), .B1(new_n729), .B2(KEYINPUT108), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n728), .B(new_n729), .C1(KEYINPUT108), .C2(KEYINPUT47), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1330gat));
  OR3_X1    g533(.A1(new_n714), .A2(new_n484), .A3(new_n380), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n484), .B1(new_n692), .B2(new_n380), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n737), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n714), .A2(new_n484), .A3(new_n380), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT48), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(G1331gat));
  NAND2_X1  g541(.A1(new_n706), .A2(new_n707), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n414), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n641), .A2(new_n642), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n745), .A2(new_n598), .A3(new_n599), .ZN(new_n746));
  INV_X1    g545(.A(new_n712), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n746), .A2(KEYINPUT109), .A3(new_n747), .A4(new_n660), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n594), .A2(new_n597), .ZN(new_n750));
  INV_X1    g549(.A(new_n595), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n752), .A2(new_n747), .A3(new_n643), .A4(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n749), .B1(new_n754), .B2(new_n661), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n748), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n744), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n666), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g559(.A(new_n458), .B(new_n757), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1333gat));
  NAND3_X1  g562(.A1(new_n758), .A2(KEYINPUT111), .A3(new_n680), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n757), .B2(new_n681), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n766), .A3(new_n608), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n744), .A2(G71gat), .A3(new_n756), .A4(new_n466), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT110), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n767), .A2(new_n769), .A3(new_n771), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1334gat));
  NOR2_X1   g574(.A1(new_n757), .A2(new_n380), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n609), .ZN(G1335gat));
  NAND2_X1  g576(.A1(new_n709), .A2(new_n711), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n643), .A2(new_n712), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n660), .ZN(new_n780));
  NOR4_X1   g579(.A1(new_n778), .A2(new_n345), .A3(new_n716), .A4(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n744), .A2(new_n710), .A3(new_n779), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT51), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n744), .A2(new_n784), .A3(new_n710), .A4(new_n779), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n783), .A2(new_n660), .A3(new_n666), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n781), .B1(new_n345), .B2(new_n786), .ZN(G1336gat));
  INV_X1    g586(.A(new_n780), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n709), .A2(new_n711), .A3(new_n277), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G92gat), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n458), .A2(G92gat), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n783), .A2(new_n660), .A3(new_n785), .A4(new_n791), .ZN(new_n792));
  AOI211_X1 g591(.A(KEYINPUT113), .B(KEYINPUT52), .C1(new_n790), .C2(new_n792), .ZN(new_n793));
  OR2_X1    g592(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n794));
  NAND2_X1  g593(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n795));
  AND4_X1   g594(.A1(new_n794), .A2(new_n790), .A3(new_n795), .A4(new_n792), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n793), .A2(new_n796), .ZN(G1337gat));
  NOR3_X1   g596(.A1(new_n778), .A2(new_n465), .A3(new_n780), .ZN(new_n798));
  INV_X1    g597(.A(G99gat), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n783), .A2(new_n799), .A3(new_n660), .A4(new_n785), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n798), .A2(new_n799), .B1(new_n800), .B2(new_n681), .ZN(G1338gat));
  INV_X1    g600(.A(new_n380), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n783), .A2(new_n802), .A3(new_n660), .A4(new_n785), .ZN(new_n803));
  INV_X1    g602(.A(G106gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n380), .A2(new_n804), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n709), .A2(new_n711), .A3(new_n788), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n805), .A2(new_n807), .A3(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(G1339gat));
  OAI21_X1  g611(.A(new_n538), .B1(new_n545), .B2(new_n527), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n536), .A2(new_n538), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n813), .A2(new_n530), .B1(new_n814), .B2(new_n540), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT115), .B1(new_n815), .B2(new_n476), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817));
  INV_X1    g616(.A(new_n476), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n524), .A2(new_n525), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n539), .A2(new_n541), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n816), .A2(new_n549), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n651), .A2(new_n652), .A3(new_n645), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT54), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n653), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n651), .A2(new_n652), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n644), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(KEYINPUT114), .A3(KEYINPUT54), .A4(new_n823), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n830), .A3(new_n658), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n655), .B2(new_n659), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n827), .A2(new_n830), .A3(new_n832), .A4(new_n658), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n822), .A2(new_n660), .B1(new_n712), .B2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(new_n598), .A3(new_n599), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n836), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n752), .B2(new_n753), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n745), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n746), .A2(new_n747), .A3(new_n661), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n716), .A2(new_n405), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n458), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n557), .ZN(new_n846));
  OAI21_X1  g645(.A(G113gat), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n844), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n843), .A2(KEYINPUT116), .A3(new_n844), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n458), .A3(new_n851), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(G113gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n847), .B1(new_n853), .B2(new_n747), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n845), .B2(new_n661), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n852), .A2(G120gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n661), .ZN(G1341gat));
  INV_X1    g656(.A(G127gat), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n845), .A2(new_n858), .A3(new_n745), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n852), .A2(new_n745), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(new_n858), .ZN(G1342gat));
  OR2_X1    g660(.A1(new_n852), .A2(G134gat), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT56), .B1(new_n862), .B2(new_n600), .ZN(new_n863));
  OR4_X1    g662(.A1(KEYINPUT56), .A2(new_n852), .A3(G134gat), .A4(new_n600), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n845), .B2(new_n600), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G1343gat));
  NAND3_X1  g665(.A1(new_n666), .A2(new_n458), .A3(new_n465), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT117), .Z(new_n868));
  NAND2_X1  g667(.A1(new_n802), .A2(KEYINPUT57), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n551), .A2(new_n556), .A3(new_n836), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n816), .A2(new_n549), .A3(new_n660), .A4(new_n821), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n600), .ZN(new_n873));
  AND4_X1   g672(.A1(new_n549), .A2(new_n836), .A3(new_n816), .A4(new_n821), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n598), .B2(new_n599), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(KEYINPUT118), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n872), .A2(new_n877), .A3(new_n600), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n745), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n869), .B1(new_n879), .B2(new_n842), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n843), .B2(new_n802), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n557), .B(new_n868), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n754), .A2(new_n660), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n878), .A2(new_n745), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n876), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n712), .A2(new_n836), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n871), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n752), .A3(new_n753), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n643), .B1(new_n890), .B2(new_n875), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n802), .B1(new_n891), .B2(new_n885), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n887), .A2(new_n869), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n894), .A2(KEYINPUT119), .A3(new_n557), .A4(new_n868), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n884), .A2(G141gat), .A3(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n892), .A2(new_n867), .ZN(new_n897));
  OR3_X1    g696(.A1(new_n897), .A2(G141gat), .A3(new_n846), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n712), .B(new_n868), .C1(new_n880), .C2(new_n881), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G141gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n898), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT58), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n901), .A2(new_n905), .ZN(G1344gat));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  INV_X1    g706(.A(G148gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n840), .B1(new_n600), .B2(new_n872), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n909), .A2(new_n643), .B1(new_n557), .B2(new_n662), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n380), .A2(KEYINPUT57), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n910), .A2(new_n911), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n660), .A3(new_n868), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n912), .A2(KEYINPUT120), .A3(new_n660), .A4(new_n868), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n907), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n894), .A2(new_n660), .A3(new_n868), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(new_n907), .A3(G148gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n660), .A2(new_n908), .ZN(new_n920));
  OAI22_X1  g719(.A1(new_n917), .A2(new_n919), .B1(new_n897), .B2(new_n920), .ZN(G1345gat));
  NAND4_X1  g720(.A1(new_n894), .A2(G155gat), .A3(new_n643), .A4(new_n868), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n297), .B1(new_n897), .B2(new_n745), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  NAND4_X1  g723(.A1(new_n894), .A2(G162gat), .A3(new_n710), .A4(new_n868), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n298), .B1(new_n897), .B2(new_n600), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n666), .A2(new_n458), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT122), .B1(new_n928), .B2(new_n680), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n802), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(KEYINPUT122), .A3(new_n680), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n843), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n846), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n405), .B1(new_n841), .B2(new_n842), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n928), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n935), .A2(KEYINPUT121), .ZN(new_n936));
  INV_X1    g735(.A(G169gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(KEYINPUT121), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n933), .B1(new_n939), .B2(new_n747), .ZN(G1348gat));
  INV_X1    g739(.A(G176gat), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n932), .A2(new_n941), .A3(new_n661), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n936), .A2(new_n660), .A3(new_n938), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n941), .ZN(G1349gat));
  OAI21_X1  g743(.A(G183gat), .B1(new_n932), .B2(new_n745), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n934), .A2(new_n202), .A3(new_n928), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n745), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g747(.A1(new_n930), .A2(new_n710), .A3(new_n843), .A4(new_n931), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(new_n950), .A3(G190gat), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n950), .B1(new_n949), .B2(G190gat), .ZN(new_n954));
  OR3_X1    g753(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n936), .A2(new_n203), .A3(new_n710), .A4(new_n938), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n952), .B2(new_n954), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(G1351gat));
  NOR3_X1   g757(.A1(new_n666), .A2(new_n458), .A3(new_n466), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n912), .A2(new_n557), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G197gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n843), .A2(new_n802), .A3(new_n959), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n962), .A2(G197gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n961), .B1(new_n747), .B2(new_n963), .ZN(G1352gat));
  NOR3_X1   g763(.A1(new_n962), .A2(G204gat), .A3(new_n661), .ZN(new_n965));
  XOR2_X1   g764(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n966));
  OR2_X1    g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n912), .A2(new_n660), .A3(new_n959), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G204gat), .ZN(new_n969));
  NAND2_X1  g768(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n967), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n967), .A2(new_n969), .A3(KEYINPUT125), .A4(new_n971), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1353gat));
  NAND4_X1  g775(.A1(new_n912), .A2(KEYINPUT126), .A3(new_n643), .A4(new_n959), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n892), .A2(KEYINPUT57), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n643), .B1(new_n873), .B2(new_n875), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n662), .A2(new_n557), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n911), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n978), .A2(new_n981), .A3(new_n643), .A4(new_n959), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n977), .A2(new_n984), .A3(G211gat), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT63), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n977), .A2(new_n984), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n893), .A2(new_n247), .A3(new_n643), .A4(new_n959), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1354gat));
  NAND4_X1  g790(.A1(new_n912), .A2(G218gat), .A3(new_n710), .A4(new_n959), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n248), .B1(new_n962), .B2(new_n600), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g793(.A(new_n994), .B(KEYINPUT127), .Z(G1355gat));
endmodule


