//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT18), .ZN(new_n203));
  INV_X1    g002(.A(G29gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT14), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n206), .B(new_n208), .C1(new_n204), .C2(new_n205), .ZN(new_n209));
  INV_X1    g008(.A(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G43gat), .ZN(new_n211));
  INV_X1    g010(.A(G43gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G50gat), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT15), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n217), .B(new_n218), .C1(new_n216), .C2(new_n213), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT85), .B1(new_n209), .B2(new_n214), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n209), .A2(new_n214), .A3(KEYINPUT85), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(G1gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G1gat), .B2(new_n226), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(KEYINPUT87), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT87), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n220), .B(new_n234), .C1(new_n221), .C2(new_n222), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n224), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT88), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n233), .A2(new_n238), .A3(new_n224), .A4(new_n235), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n232), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT89), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n233), .A2(new_n235), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(new_n231), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n203), .B1(new_n245), .B2(KEYINPUT90), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT90), .ZN(new_n247));
  NOR4_X1   g046(.A1(new_n240), .A2(new_n247), .A3(new_n242), .A4(new_n244), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n202), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n237), .A2(new_n239), .ZN(new_n250));
  INV_X1    g049(.A(new_n232), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n244), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n242), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n247), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(KEYINPUT90), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n255), .A2(KEYINPUT91), .A3(new_n256), .A4(new_n203), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(KEYINPUT18), .A3(new_n253), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n243), .B(new_n231), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n242), .B(KEYINPUT13), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n249), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G113gat), .B(G141gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(G197gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT11), .B(G169gat), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n265), .B(new_n266), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT12), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT90), .B1(new_n252), .B2(new_n253), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n270), .A2(new_n248), .A3(KEYINPUT18), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n258), .A2(new_n261), .A3(new_n268), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT92), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n203), .A3(new_n256), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n258), .A2(new_n261), .A3(new_n268), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT92), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n263), .A2(new_n269), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT27), .B(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT68), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n281), .B(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT26), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n289), .B(new_n290), .C1(new_n287), .C2(new_n286), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n288), .B1(new_n285), .B2(KEYINPUT23), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n296), .A2(G169gat), .A3(G176gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G169gat), .ZN(new_n299));
  INV_X1    g098(.A(G176gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT23), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n296), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT65), .A4(new_n288), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n290), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT64), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n306), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT64), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(new_n303), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n301), .A2(new_n302), .A3(new_n288), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n305), .A2(new_n308), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n314), .A2(KEYINPUT66), .A3(new_n315), .A4(KEYINPUT25), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT66), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT25), .A4(new_n288), .ZN(new_n318));
  AND2_X1   g117(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n290), .A2(new_n304), .B1(new_n319), .B2(G190gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n313), .A2(new_n322), .A3(KEYINPUT67), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT67), .B1(new_n313), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n293), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G120gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G113gat), .ZN(new_n327));
  INV_X1    g126(.A(G113gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G120gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G127gat), .B(G134gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n331), .B1(new_n332), .B2(new_n330), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n325), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n293), .B(new_n336), .C1(new_n323), .C2(new_n324), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G227gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G71gat), .B(G99gat), .Z(new_n344));
  XNOR2_X1  g143(.A(G15gat), .B(G43gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n346), .A2(KEYINPUT69), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(KEYINPUT69), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(KEYINPUT33), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n341), .B1(new_n338), .B2(new_n339), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT32), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n346), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n351), .A2(KEYINPUT33), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT34), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n338), .A2(new_n356), .A3(new_n341), .A4(new_n339), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n357), .B(KEYINPUT71), .Z(new_n358));
  NAND3_X1  g157(.A1(new_n338), .A2(new_n341), .A3(new_n339), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n359), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT70), .B1(new_n359), .B2(KEYINPUT34), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n355), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n343), .A2(KEYINPUT32), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT33), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n343), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n366), .A3(new_n346), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n359), .A2(KEYINPUT34), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT70), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n359), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT71), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n367), .A2(new_n372), .A3(new_n373), .A4(new_n350), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT72), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT36), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G197gat), .B(G204gat), .ZN(new_n379));
  INV_X1    g178(.A(G211gat), .ZN(new_n380));
  INV_X1    g179(.A(G218gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n379), .B1(KEYINPUT22), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G211gat), .B(G218gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n313), .A2(new_n322), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n293), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n293), .A2(KEYINPUT74), .A3(new_n386), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n325), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT73), .B(new_n391), .C1(new_n325), .C2(new_n394), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n385), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT75), .ZN(new_n401));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n394), .A3(new_n390), .A4(new_n392), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT67), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n386), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n313), .A2(new_n322), .A3(KEYINPUT67), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n292), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n391), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n385), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n399), .A2(new_n404), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n403), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n399), .A2(KEYINPUT30), .A3(new_n404), .A4(new_n412), .ZN(new_n418));
  XOR2_X1   g217(.A(G1gat), .B(G29gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT0), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT76), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n334), .B2(new_n335), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n330), .A2(new_n332), .ZN(new_n425));
  INV_X1    g224(.A(new_n331), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(KEYINPUT76), .A3(new_n333), .ZN(new_n428));
  XOR2_X1   g227(.A(G141gat), .B(G148gat), .Z(new_n429));
  INV_X1    g228(.A(G155gat), .ZN(new_n430));
  INV_X1    g229(.A(G162gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G155gat), .A2(G162gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(KEYINPUT2), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G141gat), .B(G148gat), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n433), .B(new_n432), .C1(new_n437), .C2(KEYINPUT2), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n428), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n427), .A2(new_n438), .A3(new_n436), .A4(new_n333), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G225gat), .A2(G233gat), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n439), .A2(KEYINPUT3), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT3), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n436), .A2(new_n438), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n446), .A2(new_n424), .A3(new_n428), .A4(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n441), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n439), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT4), .A3(new_n336), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n449), .A2(new_n443), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n445), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n441), .A2(KEYINPUT4), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT79), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n452), .A2(new_n336), .A3(new_n450), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT79), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n441), .A2(new_n461), .A3(KEYINPUT4), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n424), .A2(new_n428), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n436), .A2(new_n438), .A3(new_n447), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n447), .B1(new_n436), .B2(new_n438), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n444), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(new_n468), .A3(new_n455), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n422), .B1(new_n457), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT6), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n457), .A2(new_n469), .A3(new_n422), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n471), .B1(new_n474), .B2(new_n470), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n415), .A2(new_n417), .A3(new_n418), .A4(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n447), .B1(new_n385), .B2(KEYINPUT29), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n439), .ZN(new_n478));
  NAND2_X1  g277(.A1(G228gat), .A2(G233gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n448), .A2(new_n394), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n385), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT80), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n448), .A2(KEYINPUT80), .A3(new_n394), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n385), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n479), .B1(new_n478), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT31), .B(G50gat), .ZN(new_n489));
  OR3_X1    g288(.A1(new_n483), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G78gat), .B(G106gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(G22gat), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n489), .B1(new_n483), .B2(new_n488), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n490), .B2(new_n493), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n476), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n375), .A2(KEYINPUT72), .A3(KEYINPUT36), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n378), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n443), .B1(new_n463), .B2(new_n449), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n422), .B(KEYINPUT81), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT39), .B1(new_n442), .B2(new_n444), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT82), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n502), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n511), .B(new_n502), .C1(new_n507), .C2(new_n509), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n457), .A2(new_n469), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(new_n506), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n496), .ZN(new_n518));
  INV_X1    g317(.A(new_n471), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n506), .B1(new_n457), .B2(new_n469), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n474), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n521), .B2(KEYINPUT83), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT83), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n474), .B2(new_n520), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n413), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT37), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n405), .A2(new_n410), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(new_n385), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n397), .A2(new_n398), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(new_n385), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n530), .B(new_n403), .C1(new_n416), .C2(KEYINPUT37), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT38), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n416), .B2(KEYINPUT37), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n390), .B1(new_n409), .B2(KEYINPUT29), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n395), .A2(new_n396), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(new_n393), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n411), .B1(new_n538), .B2(new_n385), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n404), .B1(new_n539), .B2(new_n526), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n525), .B1(new_n533), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n518), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n500), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n363), .A2(new_n374), .A3(new_n496), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT35), .B1(new_n545), .B2(new_n476), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT84), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT84), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n548), .B(KEYINPUT35), .C1(new_n545), .C2(new_n476), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT35), .B1(new_n522), .B2(new_n524), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n551), .A2(new_n496), .A3(new_n374), .A4(new_n363), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(new_n501), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n278), .B1(new_n544), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n557));
  INV_X1    g356(.A(G64gat), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n558), .A2(G57gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(G57gat), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  OAI22_X1  g362(.A1(new_n557), .A2(KEYINPUT93), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n561), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G127gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n231), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n572), .B1(KEYINPUT21), .B2(new_n565), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n571), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT95), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n430), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n576), .B(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n574), .A2(new_n579), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G99gat), .B(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n586), .A2(KEYINPUT7), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT96), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(KEYINPUT7), .A3(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n593), .B2(KEYINPUT97), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n585), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n593), .A2(KEYINPUT97), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n589), .A2(new_n593), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n601), .A2(new_n584), .A3(new_n602), .A4(new_n598), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n583), .B1(new_n243), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT98), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n250), .A2(new_n225), .A3(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G190gat), .B(G218gat), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n611), .A3(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n610), .A2(new_n616), .A3(new_n612), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n566), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n600), .A2(new_n603), .A3(new_n565), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n626), .A2(new_n625), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n623), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n637), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n582), .A2(new_n621), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n475), .B(KEYINPUT100), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n556), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  INV_X1    g446(.A(new_n501), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  AND3_X1   g449(.A1(new_n649), .A2(new_n556), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n230), .B1(new_n649), .B2(new_n556), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT42), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(KEYINPUT42), .B2(new_n651), .ZN(G1325gat));
  NAND2_X1  g453(.A1(new_n556), .A2(new_n644), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n378), .A2(new_n499), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT101), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(G15gat), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n375), .A2(G15gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n556), .A2(new_n644), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(G1326gat));
  NOR2_X1   g461(.A1(new_n655), .A2(new_n496), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT102), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  INV_X1    g465(.A(new_n582), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n667), .A2(new_n620), .A3(new_n641), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n556), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n204), .A3(new_n645), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT45), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n582), .B(KEYINPUT103), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(new_n278), .A3(new_n641), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n550), .B2(new_n554), .ZN(new_n676));
  AOI211_X1 g475(.A(KEYINPUT104), .B(new_n553), .C1(new_n547), .C2(new_n549), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n544), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n620), .A2(KEYINPUT44), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n500), .A2(new_n543), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n553), .B1(new_n547), .B2(new_n549), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n621), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(KEYINPUT44), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n674), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n645), .ZN(new_n686));
  OAI21_X1  g485(.A(G29gat), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n687), .ZN(G1328gat));
  NOR3_X1   g487(.A1(new_n669), .A2(G36gat), .A3(new_n648), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT46), .ZN(new_n690));
  OAI21_X1  g489(.A(G36gat), .B1(new_n685), .B2(new_n648), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(G1329gat));
  NOR2_X1   g491(.A1(new_n375), .A2(G43gat), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n556), .A2(new_n668), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT106), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT108), .B1(new_n685), .B2(new_n656), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G43gat), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n685), .A2(KEYINPUT108), .A3(new_n656), .ZN(new_n698));
  OAI211_X1 g497(.A(KEYINPUT47), .B(new_n695), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n678), .A2(new_n679), .B1(KEYINPUT44), .B2(new_n683), .ZN(new_n701));
  INV_X1    g500(.A(new_n674), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(new_n658), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n703), .B2(new_n212), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n657), .B(new_n674), .C1(new_n680), .C2(new_n684), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(KEYINPUT105), .A3(G43gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n706), .A3(new_n695), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n699), .B1(new_n710), .B2(new_n711), .ZN(G1330gat));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n685), .A2(new_n496), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n210), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT48), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n670), .A2(new_n210), .A3(new_n497), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n714), .B2(new_n210), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n716), .B(new_n718), .ZN(G1331gat));
  INV_X1    g518(.A(new_n678), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n278), .A2(new_n667), .A3(new_n620), .A4(new_n641), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n645), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT110), .B(G57gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1332gat));
  NAND2_X1  g524(.A1(new_n722), .A2(KEYINPUT111), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n720), .B2(new_n721), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n648), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n730), .A2(KEYINPUT112), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(KEYINPUT112), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(G1333gat));
  AND2_X1   g535(.A1(new_n726), .A2(new_n728), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(G71gat), .A3(new_n657), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n720), .A2(new_n375), .A3(new_n721), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n739), .A2(G71gat), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n738), .A2(KEYINPUT50), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT50), .B1(new_n738), .B2(new_n740), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n737), .A2(new_n497), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  INV_X1    g544(.A(new_n278), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n667), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n641), .B(new_n747), .C1(new_n680), .C2(new_n684), .ZN(new_n748));
  OAI21_X1  g547(.A(G85gat), .B1(new_n748), .B2(new_n686), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n621), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n720), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n678), .A2(KEYINPUT51), .A3(new_n621), .A4(new_n747), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n645), .A2(new_n596), .A3(new_n641), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n749), .B1(new_n755), .B2(new_n756), .ZN(G1336gat));
  INV_X1    g556(.A(new_n641), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n648), .A2(G92gat), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n754), .A2(new_n759), .B1(new_n760), .B2(KEYINPUT52), .ZN(new_n761));
  OAI21_X1  g560(.A(G92gat), .B1(new_n748), .B2(new_n648), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n760), .A2(KEYINPUT52), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n763), .B(new_n764), .Z(G1337gat));
  OAI21_X1  g564(.A(G99gat), .B1(new_n748), .B2(new_n658), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n375), .A2(G99gat), .A3(new_n758), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n755), .B2(new_n767), .ZN(G1338gat));
  OAI21_X1  g567(.A(G106gat), .B1(new_n748), .B2(new_n496), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n758), .A2(new_n496), .A3(G106gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n627), .A2(new_n628), .A3(new_n623), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n775), .A2(new_n629), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n629), .A2(new_n776), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(new_n637), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n778), .A3(new_n637), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n638), .B1(new_n783), .B2(KEYINPUT55), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785));
  INV_X1    g584(.A(new_n782), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n780), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n787), .B2(new_n777), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n263), .A2(new_n269), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n273), .A2(new_n277), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n259), .A2(new_n260), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n242), .B1(new_n240), .B2(new_n244), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(new_n267), .ZN(new_n796));
  AOI211_X1 g595(.A(new_n796), .B(new_n758), .C1(new_n273), .C2(new_n277), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n620), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n784), .A2(new_n618), .A3(new_n788), .A4(new_n619), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n796), .B1(new_n273), .B2(new_n277), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n796), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n791), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT115), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n673), .B1(new_n798), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n642), .A2(new_n278), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n774), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n791), .A2(new_n641), .A3(new_n803), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n278), .B2(new_n789), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n812), .A2(new_n620), .B1(new_n802), .B2(new_n805), .ZN(new_n813));
  OAI211_X1 g612(.A(KEYINPUT116), .B(new_n808), .C1(new_n813), .C2(new_n673), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n545), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n686), .A2(new_n501), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n278), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(new_n328), .ZN(G1340gat));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n758), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(new_n326), .ZN(G1341gat));
  INV_X1    g621(.A(new_n673), .ZN(new_n823));
  OAI21_X1  g622(.A(G127gat), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n582), .A2(G127gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n818), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT117), .Z(G1342gat));
  NOR2_X1   g626(.A1(new_n620), .A2(new_n501), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n686), .A2(G134gat), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n815), .A2(new_n816), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT56), .Z(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n818), .B2(new_n620), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1343gat));
  INV_X1    g632(.A(G141gat), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n656), .A2(new_n817), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n497), .A2(KEYINPUT57), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n789), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n746), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n621), .B1(new_n839), .B2(new_n811), .ZN(new_n840));
  INV_X1    g639(.A(new_n806), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n582), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n836), .B1(new_n842), .B2(new_n808), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n810), .A2(new_n497), .A3(new_n814), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n843), .B1(new_n846), .B2(KEYINPUT118), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(new_n848), .A3(new_n845), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n835), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n834), .B1(new_n850), .B2(new_n746), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n844), .A2(new_n686), .A3(new_n657), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n648), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n746), .A2(new_n834), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT58), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  INV_X1    g656(.A(new_n855), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n278), .B(new_n835), .C1(new_n847), .C2(new_n849), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n834), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n860), .ZN(G1344gat));
  INV_X1    g660(.A(G148gat), .ZN(new_n862));
  AOI211_X1 g661(.A(KEYINPUT59), .B(new_n862), .C1(new_n850), .C2(new_n641), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n842), .B1(new_n643), .B2(new_n746), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n497), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n845), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n815), .A2(KEYINPUT57), .A3(new_n497), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n835), .A2(KEYINPUT122), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n758), .B1(new_n835), .B2(KEYINPUT122), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n864), .B1(new_n872), .B2(G148gat), .ZN(new_n873));
  INV_X1    g672(.A(new_n853), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n758), .A2(G148gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(KEYINPUT120), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(KEYINPUT120), .ZN(new_n878));
  OAI22_X1  g677(.A1(new_n863), .A2(new_n873), .B1(new_n877), .B2(new_n878), .ZN(G1345gat));
  NAND3_X1  g678(.A1(new_n874), .A2(new_n430), .A3(new_n667), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n850), .A2(new_n673), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n430), .ZN(G1346gat));
  NAND3_X1  g681(.A1(new_n852), .A2(new_n431), .A3(new_n828), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n850), .A2(new_n621), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n431), .ZN(G1347gat));
  AND2_X1   g684(.A1(new_n815), .A2(new_n686), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n648), .A2(new_n545), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G169gat), .B1(new_n888), .B2(new_n278), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT124), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n887), .B(KEYINPUT123), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n299), .A3(new_n746), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(new_n894), .ZN(G1348gat));
  OAI21_X1  g694(.A(G176gat), .B1(new_n888), .B2(new_n758), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n641), .A2(new_n300), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n892), .B2(new_n897), .ZN(G1349gat));
  OAI21_X1  g697(.A(G183gat), .B1(new_n888), .B2(new_n823), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n886), .A2(new_n279), .A3(new_n667), .A4(new_n891), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT60), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n899), .A2(new_n900), .A3(new_n904), .A4(new_n901), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n888), .B2(new_n620), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT61), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n280), .A3(new_n621), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1351gat));
  NOR3_X1   g709(.A1(new_n657), .A2(new_n496), .A3(new_n648), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n815), .A2(new_n686), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(G197gat), .B1(new_n913), .B2(new_n746), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n657), .A2(new_n648), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n686), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n916), .B1(new_n867), .B2(new_n868), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n746), .A2(G197gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(G1352gat));
  INV_X1    g718(.A(new_n917), .ZN(new_n920));
  OAI21_X1  g719(.A(G204gat), .B1(new_n920), .B2(new_n758), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n758), .A2(G204gat), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT62), .B1(new_n912), .B2(new_n922), .ZN(new_n923));
  OR3_X1    g722(.A1(new_n912), .A2(KEYINPUT62), .A3(new_n922), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(G1353gat));
  NAND3_X1  g724(.A1(new_n913), .A2(new_n380), .A3(new_n667), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n917), .A2(new_n667), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n927), .B2(G211gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(G1354gat));
  AOI211_X1 g729(.A(new_n381), .B(new_n620), .C1(new_n917), .C2(KEYINPUT127), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n917), .A2(KEYINPUT127), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n381), .B1(new_n912), .B2(new_n620), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  AOI22_X1  g735(.A1(new_n931), .A2(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G1355gat));
endmodule


