//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(G104), .B(G107), .Z(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G101), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT81), .B1(new_n190), .B2(G104), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT81), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(new_n192), .A3(G107), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n190), .A3(G104), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n195), .A4(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n189), .B1(new_n198), .B2(G101), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G116), .B(G119), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT2), .B(G113), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G113), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n209), .A2(G116), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n207), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n205), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n189), .B(KEYINPUT83), .C1(new_n198), .C2(G101), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n201), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n216), .B1(new_n198), .B2(G101), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n193), .A2(new_n197), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n218), .A2(new_n219), .A3(new_n191), .A4(new_n195), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n202), .B(new_n204), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n198), .A2(new_n216), .A3(G101), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G110), .B(G122), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n215), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G953), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G224), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT7), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G143), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G146), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT64), .B(G143), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n232), .A2(KEYINPUT64), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G143), .ZN(new_n243));
  AOI21_X1  g057(.A(G146), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(G143), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n232), .A2(KEYINPUT65), .A3(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n240), .B1(new_n244), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n238), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G125), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  OAI21_X1  g068(.A(G128), .B1(new_n233), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n244), .B2(new_n249), .ZN(new_n256));
  INV_X1    g070(.A(new_n233), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n241), .A2(new_n243), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n257), .B(new_n259), .C1(new_n260), .C2(new_n246), .ZN(new_n261));
  AOI21_X1  g075(.A(G125), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n231), .B1(new_n253), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n262), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(new_n230), .C1(new_n252), .C2(new_n251), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n227), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  XOR2_X1   g080(.A(new_n226), .B(KEYINPUT8), .Z(new_n267));
  INV_X1    g081(.A(new_n199), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n213), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n202), .A2(KEYINPUT5), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n205), .B1(new_n211), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n201), .A2(new_n271), .A3(new_n214), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n267), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n187), .B1(new_n266), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT85), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(KEYINPUT85), .B(new_n187), .C1(new_n266), .C2(new_n273), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n215), .A2(new_n225), .ZN(new_n278));
  INV_X1    g092(.A(new_n226), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT6), .A3(new_n227), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n264), .B1(new_n252), .B2(new_n251), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n282), .B(new_n229), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n278), .A2(new_n284), .A3(new_n279), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n281), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n276), .A2(new_n277), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G210), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n276), .A2(new_n288), .A3(new_n277), .A4(new_n286), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(KEYINPUT86), .A3(new_n291), .ZN(new_n292));
  OR3_X1    g106(.A1(new_n287), .A2(KEYINPUT86), .A3(new_n289), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G214), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  OAI21_X1  g112(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT1), .B1(new_n234), .B2(G146), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n258), .B1(new_n301), .B2(KEYINPUT82), .ZN(new_n302));
  OR3_X1    g116(.A1(new_n244), .A2(KEYINPUT82), .A3(new_n254), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n235), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n261), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n268), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n256), .A2(new_n261), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n201), .A2(KEYINPUT10), .A3(new_n309), .A4(new_n214), .ZN(new_n310));
  OR2_X1    g124(.A1(new_n237), .A2(new_n239), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n247), .A2(new_n248), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n242), .A2(G143), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n232), .A2(KEYINPUT64), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n246), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  AOI211_X1 g130(.A(new_n233), .B(new_n236), .C1(new_n234), .C2(G146), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n221), .A3(new_n224), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT11), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(KEYINPUT67), .ZN(new_n322));
  INV_X1    g136(.A(G134), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G137), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(KEYINPUT67), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT67), .ZN(new_n327));
  INV_X1    g141(.A(G137), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT11), .A4(G134), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(G137), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n326), .A2(new_n331), .A3(G131), .ZN(new_n332));
  INV_X1    g146(.A(G131), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n328), .A2(G134), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n324), .B2(new_n322), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n328), .A2(G134), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n333), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT68), .B1(new_n332), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G131), .B1(new_n326), .B2(new_n331), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n335), .A2(new_n333), .A3(new_n339), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n308), .A2(new_n320), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n201), .A2(new_n214), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n248), .B(new_n247), .C1(new_n234), .C2(G146), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n349), .A2(new_n255), .B1(new_n235), .B2(new_n259), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n306), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n332), .A2(new_n340), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT12), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n343), .B1(new_n342), .B2(new_n344), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT12), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n347), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G140), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT79), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n228), .A2(G227), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n364), .B(KEYINPUT80), .Z(new_n365));
  XNOR2_X1  g179(.A(new_n363), .B(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n347), .A2(new_n366), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n308), .A2(new_n320), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n359), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n361), .A2(new_n367), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G469), .B1(new_n371), .B2(G902), .ZN(new_n372));
  INV_X1    g186(.A(G469), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n352), .A2(new_n359), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n374), .A2(new_n354), .B1(new_n352), .B2(new_n355), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n347), .A2(new_n366), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n366), .B1(new_n370), .B2(new_n347), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n373), .B(new_n187), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n300), .B1(new_n372), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(G234), .A2(G237), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n381), .A2(G952), .A3(new_n228), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(G902), .A3(G953), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(KEYINPUT91), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT21), .B(G898), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n382), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(G475), .A2(G902), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n192), .ZN(new_n390));
  INV_X1    g204(.A(G237), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n228), .A3(G214), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n241), .A3(new_n243), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n391), .A2(new_n228), .A3(G143), .A4(G214), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n333), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n395), .B2(G131), .ZN(new_n399));
  AOI211_X1 g213(.A(KEYINPUT87), .B(new_n333), .C1(new_n393), .C2(new_n394), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT88), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n397), .B(new_n403), .C1(new_n399), .C2(new_n400), .ZN(new_n404));
  XNOR2_X1  g218(.A(G125), .B(G140), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT16), .ZN(new_n406));
  OR3_X1    g220(.A1(new_n252), .A2(KEYINPUT16), .A3(G140), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n406), .A2(G146), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(KEYINPUT89), .A3(KEYINPUT19), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n409), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n408), .B1(new_n246), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n402), .A2(new_n404), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n396), .B1(new_n414), .B2(new_n333), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n405), .B(new_n246), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n395), .A2(G131), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n415), .B(new_n416), .C1(new_n414), .C2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n390), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT17), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n397), .B(new_n420), .C1(new_n399), .C2(new_n400), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n417), .A2(KEYINPUT87), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n395), .A2(new_n398), .A3(G131), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(KEYINPUT17), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(G146), .B1(new_n406), .B2(new_n407), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n408), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n390), .A3(new_n418), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n388), .B1(new_n419), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT20), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n432), .B(new_n388), .C1(new_n419), .C2(new_n429), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n390), .B1(new_n427), .B2(new_n418), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n187), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n431), .A2(new_n433), .B1(G475), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT13), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n234), .A2(new_n437), .A3(G128), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n234), .A2(G128), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n258), .A2(G143), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(G134), .B(new_n438), .C1(new_n441), .C2(new_n437), .ZN(new_n442));
  XNOR2_X1  g256(.A(G116), .B(G122), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(new_n190), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n323), .A3(new_n440), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT90), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n439), .A2(KEYINPUT90), .A3(new_n323), .A4(new_n440), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n442), .A2(new_n444), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G116), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n190), .B1(new_n451), .B2(KEYINPUT14), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n443), .ZN(new_n453));
  INV_X1    g267(.A(new_n445), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n323), .B1(new_n439), .B2(new_n440), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G217), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n298), .A2(new_n458), .A3(G953), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n449), .A2(new_n456), .A3(new_n459), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n187), .ZN(new_n464));
  INV_X1    g278(.A(G478), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(KEYINPUT15), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n464), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n436), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AND4_X1   g284(.A1(new_n297), .A2(new_n380), .A3(new_n387), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n406), .A2(G146), .A3(new_n407), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n405), .A2(new_n246), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n258), .A2(G119), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n209), .A2(G128), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT74), .A4(KEYINPUT23), .ZN(new_n476));
  OR2_X1    g290(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n477));
  NAND2_X1  g291(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n477), .A2(G119), .A3(new_n258), .A4(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(G110), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n474), .A2(new_n475), .ZN(new_n481));
  XOR2_X1   g295(.A(KEYINPUT24), .B(G110), .Z(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n472), .B(new_n473), .C1(new_n480), .C2(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT73), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT73), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  OAI22_X1  g300(.A1(new_n408), .A2(new_n425), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G110), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n476), .A2(new_n479), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT75), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT75), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n476), .A2(new_n479), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n484), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT77), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT76), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT22), .B(G137), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT77), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n500), .B(new_n484), .C1(new_n487), .C2(new_n493), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n499), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n494), .A2(KEYINPUT77), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT25), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n458), .B1(G234), .B2(new_n187), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n505), .B2(new_n506), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n502), .A2(new_n504), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n508), .A2(G902), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT78), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n391), .A2(new_n228), .A3(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT26), .B(G101), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT71), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT28), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT69), .ZN(new_n524));
  OAI21_X1  g338(.A(G131), .B1(new_n324), .B2(new_n334), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n344), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n524), .B1(new_n350), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n309), .A2(KEYINPUT69), .A3(new_n344), .A4(new_n525), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n341), .A2(new_n318), .A3(new_n345), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n222), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT66), .B1(new_n316), .B2(new_n317), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT66), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n238), .A2(new_n533), .A3(new_n250), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n353), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n350), .A2(new_n526), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n223), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n523), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n536), .A2(new_n223), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT28), .B1(new_n539), .B2(new_n530), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n522), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n520), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n359), .A2(new_n318), .B1(new_n527), .B2(new_n528), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n222), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n529), .A2(KEYINPUT30), .A3(new_n530), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n535), .B2(new_n536), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n547), .A3(new_n223), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT31), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n544), .A2(new_n548), .A3(KEYINPUT70), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT70), .B1(new_n544), .B2(new_n548), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n551), .B1(new_n554), .B2(KEYINPUT31), .ZN(new_n555));
  NOR2_X1   g369(.A1(G472), .A2(G902), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT32), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n551), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT70), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n545), .A2(new_n547), .A3(new_n223), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n531), .A2(new_n520), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n544), .A2(new_n548), .A3(KEYINPUT70), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT31), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT32), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n556), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n558), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n529), .A2(new_n530), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n223), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n523), .B1(new_n571), .B2(new_n531), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n540), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n531), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n222), .B1(new_n529), .B2(new_n530), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT28), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT72), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n574), .A2(new_n578), .A3(KEYINPUT29), .A4(new_n520), .ZN(new_n579));
  OR3_X1    g393(.A1(new_n538), .A2(new_n540), .A3(new_n522), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT29), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n548), .A2(new_n531), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n542), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n579), .A2(new_n584), .A3(new_n187), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G472), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n516), .B1(new_n569), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n471), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  INV_X1    g403(.A(new_n347), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n367), .B1(new_n375), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n368), .A2(new_n370), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(G469), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(G469), .A2(G902), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n379), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n299), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n516), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n566), .A2(new_n187), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n598), .A2(G472), .B1(new_n556), .B2(new_n566), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n296), .B1(new_n290), .B2(new_n291), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n463), .A2(new_n465), .A3(new_n187), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n462), .A2(KEYINPUT92), .ZN(new_n603));
  INV_X1    g417(.A(new_n462), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n459), .B1(new_n449), .B2(new_n456), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n603), .B(KEYINPUT33), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n461), .B(new_n462), .C1(KEYINPUT92), .C2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(G902), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n602), .B1(new_n609), .B2(new_n465), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n436), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n601), .A2(new_n611), .A3(new_n387), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n600), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  NAND2_X1  g429(.A1(new_n290), .A2(new_n291), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n295), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n436), .A2(new_n467), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n617), .A2(new_n386), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n600), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT93), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT35), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G107), .ZN(G9));
  NOR2_X1   g437(.A1(new_n499), .A2(KEYINPUT36), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n494), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n514), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n511), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n471), .A2(new_n599), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT37), .B(G110), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT94), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n628), .B(new_n630), .ZN(G12));
  AOI21_X1  g445(.A(new_n567), .B1(new_n566), .B2(new_n556), .ZN(new_n632));
  AOI211_X1 g446(.A(KEYINPUT32), .B(new_n557), .C1(new_n559), .C2(new_n565), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n586), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(G900), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n384), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n382), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n436), .A2(new_n467), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n596), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n601), .A2(new_n627), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n634), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n634), .A2(new_n640), .A3(KEYINPUT95), .A4(new_n642), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  XOR2_X1   g462(.A(KEYINPUT97), .B(KEYINPUT39), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n637), .B(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n596), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT40), .Z(new_n653));
  XOR2_X1   g467(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n294), .B(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n521), .B1(new_n571), .B2(new_n531), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n552), .A2(new_n553), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n657), .B2(G902), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n569), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n627), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n436), .A2(new_n468), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n662), .A3(new_n295), .ZN(new_n663));
  OR4_X1    g477(.A1(new_n653), .A2(new_n655), .A3(new_n660), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n260), .ZN(G45));
  NAND2_X1  g479(.A1(new_n435), .A2(G475), .ZN(new_n666));
  INV_X1    g480(.A(new_n418), .ZN(new_n667));
  INV_X1    g481(.A(new_n411), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n472), .B1(new_n668), .B2(G146), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(KEYINPUT88), .B2(new_n401), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n667), .B1(new_n670), .B2(new_n404), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n428), .B1(new_n671), .B2(new_n390), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n432), .B1(new_n672), .B2(new_n388), .ZN(new_n673));
  INV_X1    g487(.A(new_n433), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n666), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n602), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n606), .A2(new_n608), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n187), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n676), .B1(new_n678), .B2(G478), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n675), .A2(new_n679), .A3(new_n638), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n617), .A2(new_n680), .A3(KEYINPUT98), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT98), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n436), .A2(new_n610), .A3(new_n637), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n682), .B1(new_n683), .B2(new_n601), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n595), .A2(new_n299), .A3(new_n627), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n569), .B2(new_n586), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  OAI21_X1  g503(.A(new_n187), .B1(new_n377), .B2(new_n378), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n691), .A2(new_n299), .A3(new_n379), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n587), .A2(KEYINPUT99), .A3(new_n612), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n516), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n634), .A2(new_n694), .A3(new_n612), .A4(new_n692), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n634), .A2(new_n619), .A3(new_n694), .A4(new_n692), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT100), .B(G116), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G18));
  NAND3_X1  g517(.A1(new_n691), .A2(new_n299), .A3(new_n379), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n386), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n634), .A2(new_n470), .A3(new_n705), .A4(new_n642), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  AND2_X1   g521(.A1(new_n574), .A2(new_n578), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n565), .B(new_n550), .C1(new_n708), .C2(new_n521), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n709), .A2(new_n556), .B1(new_n598), .B2(G472), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n516), .A2(KEYINPUT101), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n511), .A2(new_n712), .A3(new_n515), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n662), .A2(new_n601), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n710), .A2(new_n705), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  NAND2_X1  g531(.A1(new_n598), .A2(G472), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n565), .A2(new_n550), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n521), .B1(new_n574), .B2(new_n578), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n556), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n627), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n611), .A2(KEYINPUT102), .A3(new_n638), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT102), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n680), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n692), .A2(new_n601), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n722), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n252), .ZN(G27));
  INV_X1    g543(.A(new_n726), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n380), .A2(new_n294), .A3(new_n295), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n731), .A3(new_n634), .A4(new_n714), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT42), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n587), .A2(new_n730), .A3(new_n734), .A4(new_n731), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  INV_X1    g551(.A(new_n639), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n587), .A2(new_n738), .A3(new_n731), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  NOR2_X1   g554(.A1(new_n675), .A2(new_n610), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT43), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(KEYINPUT103), .Z(new_n743));
  NOR2_X1   g557(.A1(new_n599), .A2(new_n661), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n294), .A2(new_n295), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n747), .A2(new_n748), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n371), .B(KEYINPUT45), .Z(new_n753));
  OAI21_X1  g567(.A(G469), .B1(new_n753), .B2(G902), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n379), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(KEYINPUT46), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n299), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n651), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n749), .A2(new_n751), .A3(new_n752), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  XNOR2_X1  g575(.A(new_n758), .B(KEYINPUT47), .ZN(new_n762));
  OR4_X1    g576(.A1(new_n694), .A2(new_n634), .A3(new_n680), .A4(new_n750), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  AND3_X1   g579(.A1(new_n511), .A2(new_n626), .A3(new_n638), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n595), .A3(new_n299), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n662), .A2(new_n601), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n685), .A2(new_n687), .B1(new_n659), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n722), .A2(new_n726), .ZN(new_n771));
  INV_X1    g585(.A(new_n727), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n641), .B1(new_n569), .B2(new_n586), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT95), .B1(new_n774), .B2(new_n640), .ZN(new_n775));
  INV_X1    g589(.A(new_n646), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n770), .B(new_n773), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n728), .B1(new_n645), .B2(new_n646), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(KEYINPUT52), .A3(new_n770), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT107), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n695), .B(KEYINPUT99), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n701), .A2(new_n706), .A3(new_n716), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n611), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n618), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n600), .A2(new_n297), .A3(new_n387), .A4(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n628), .A2(new_n789), .A3(new_n588), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n785), .B1(new_n693), .B2(new_n697), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n791), .B2(KEYINPUT107), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n470), .A2(new_n627), .A3(new_n638), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n569), .B2(new_n586), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n731), .B1(new_n771), .B2(new_n794), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n733), .A2(new_n795), .A3(new_n735), .A4(new_n739), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n782), .A2(new_n786), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n785), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n698), .A3(KEYINPUT107), .ZN(new_n801));
  INV_X1    g615(.A(new_n790), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n786), .A2(new_n796), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT108), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n778), .B1(new_n769), .B2(new_n659), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n780), .A2(KEYINPUT109), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n780), .A2(KEYINPUT109), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n688), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n779), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n803), .A2(new_n804), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n805), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n799), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n790), .A2(new_n813), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n791), .A3(new_n796), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n809), .B2(new_n779), .ZN(new_n820));
  AND4_X1   g634(.A1(KEYINPUT52), .A2(new_n647), .A3(new_n773), .A4(new_n770), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(new_n780), .B2(new_n770), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n798), .B1(new_n803), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(KEYINPUT112), .B(new_n798), .C1(new_n803), .C2(new_n823), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n820), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n829));
  AOI22_X1  g643(.A1(new_n817), .A2(KEYINPUT54), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n382), .A2(new_n742), .A3(new_n710), .A4(new_n714), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n296), .A3(new_n655), .A4(new_n692), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT50), .Z(new_n833));
  NOR2_X1   g647(.A1(new_n750), .A2(new_n704), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n660), .A2(new_n694), .A3(new_n382), .A4(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n675), .A3(new_n679), .ZN(new_n836));
  INV_X1    g650(.A(new_n722), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n834), .A2(new_n382), .A3(new_n742), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n831), .A2(new_n751), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n691), .A2(new_n300), .A3(new_n379), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n762), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT51), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT115), .ZN(new_n846));
  MUX2_X1   g660(.A(new_n846), .B(KEYINPUT115), .S(new_n840), .Z(new_n847));
  XOR2_X1   g661(.A(new_n762), .B(KEYINPUT114), .Z(new_n848));
  AOI21_X1  g662(.A(new_n841), .B1(new_n848), .B2(new_n842), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n844), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n228), .A2(G952), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n831), .B2(new_n772), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT48), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n634), .A2(new_n714), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n838), .A2(new_n854), .ZN(new_n855));
  OAI221_X1 g669(.A(new_n852), .B1(new_n853), .B2(new_n855), .C1(new_n787), .C2(new_n835), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n853), .B2(new_n855), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n830), .A2(new_n850), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(G952), .A2(G953), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n714), .A2(new_n295), .A3(new_n299), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n860), .A2(KEYINPUT105), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n741), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(KEYINPUT105), .B2(new_n860), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT106), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n691), .A2(new_n379), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT49), .Z(new_n868));
  NAND4_X1  g682(.A1(new_n866), .A2(new_n655), .A3(new_n660), .A4(new_n868), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n858), .A2(new_n859), .B1(new_n865), .B2(new_n869), .ZN(G75));
  NAND2_X1  g684(.A1(new_n281), .A2(new_n285), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(new_n283), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n828), .A2(new_n187), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(G210), .ZN(new_n875));
  NOR2_X1   g689(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n873), .A3(new_n876), .ZN(new_n879));
  XOR2_X1   g693(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n878), .B2(new_n879), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n228), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  AND3_X1   g699(.A1(new_n874), .A2(G469), .A3(new_n753), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n377), .A2(new_n378), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT119), .B1(new_n828), .B2(new_n829), .ZN(new_n888));
  INV_X1    g702(.A(new_n820), .ZN(new_n889));
  INV_X1    g703(.A(new_n827), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT112), .B1(new_n797), .B2(new_n798), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  INV_X1    g707(.A(new_n829), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n889), .B(new_n829), .C1(new_n890), .C2(new_n891), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT118), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n828), .A2(new_n899), .A3(new_n829), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n594), .B(KEYINPUT57), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n887), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n886), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n896), .B2(new_n901), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT120), .B1(new_n908), .B2(new_n887), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n884), .B1(new_n907), .B2(new_n909), .ZN(G54));
  NAND3_X1  g724(.A1(new_n874), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  INV_X1    g725(.A(new_n672), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n884), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n913), .A2(new_n918), .A3(new_n914), .A4(new_n915), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(G60));
  INV_X1    g734(.A(new_n902), .ZN(new_n921));
  INV_X1    g735(.A(new_n677), .ZN(new_n922));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT59), .Z(new_n924));
  OR2_X1    g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n914), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n830), .A2(new_n924), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n922), .ZN(G63));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n930));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n828), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n512), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT123), .B1(new_n934), .B2(new_n884), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n625), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n934), .A2(KEYINPUT123), .A3(new_n884), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n929), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n884), .A2(new_n929), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n936), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n939), .B1(new_n940), .B2(new_n943), .ZN(G66));
  NAND2_X1  g758(.A1(new_n792), .A2(new_n786), .ZN(new_n945));
  NAND2_X1  g759(.A1(G224), .A2(G953), .ZN(new_n946));
  OAI22_X1  g760(.A1(new_n945), .A2(G953), .B1(new_n385), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT125), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n871), .B1(G898), .B2(new_n228), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT126), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  AOI21_X1  g765(.A(new_n228), .B1(G227), .B2(G900), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n545), .A2(new_n547), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n411), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n807), .A2(new_n808), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n664), .A3(new_n688), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n587), .A2(new_n652), .A3(new_n751), .A4(new_n788), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n764), .A2(new_n760), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n955), .B1(new_n961), .B2(G953), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n764), .A2(new_n760), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n956), .A2(new_n688), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n759), .A2(new_n715), .A3(new_n854), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n965), .A2(new_n736), .A3(new_n739), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n228), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n955), .B1(G900), .B2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n953), .B1(new_n962), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n971), .B(new_n972), .Z(G72));
  NOR2_X1   g787(.A1(new_n582), .A2(new_n520), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n542), .B1(new_n548), .B2(new_n531), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT63), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n884), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n961), .A2(new_n975), .B1(new_n967), .B2(new_n974), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n979), .B1(new_n980), .B2(new_n945), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n978), .B1(new_n554), .B2(new_n583), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n817), .B2(new_n982), .ZN(G57));
endmodule


