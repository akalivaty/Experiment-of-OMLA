

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729;

  AND2_X1 U367 ( .A1(n715), .A2(n410), .ZN(n365) );
  NOR2_X1 U368 ( .A1(G902), .A2(n691), .ZN(n467) );
  INV_X1 U369 ( .A(G953), .ZN(n707) );
  NOR2_X2 U370 ( .A1(n537), .A2(n432), .ZN(n554) );
  NOR2_X2 U371 ( .A1(n670), .A2(n671), .ZN(n542) );
  XNOR2_X2 U372 ( .A(n584), .B(n583), .ZN(n726) );
  XNOR2_X2 U373 ( .A(n563), .B(n351), .ZN(n541) );
  XNOR2_X2 U374 ( .A(n472), .B(G134), .ZN(n505) );
  XNOR2_X2 U375 ( .A(n360), .B(G128), .ZN(n472) );
  XNOR2_X2 U376 ( .A(n536), .B(KEYINPUT107), .ZN(n537) );
  AND2_X2 U377 ( .A1(n586), .A2(n429), .ZN(n536) );
  AND2_X2 U378 ( .A1(n606), .A2(n605), .ZN(n693) );
  NAND2_X1 U379 ( .A1(n409), .A2(n354), .ZN(n606) );
  AND2_X1 U380 ( .A1(n373), .A2(n372), .ZN(n371) );
  NAND2_X1 U381 ( .A1(n436), .A2(n591), .ZN(n435) );
  XNOR2_X1 U382 ( .A(n431), .B(n430), .ZN(n556) );
  OR2_X1 U383 ( .A1(n589), .A2(n656), .ZN(n573) );
  NAND2_X1 U384 ( .A1(n585), .A2(n586), .ZN(n661) );
  XNOR2_X1 U385 ( .A(n427), .B(KEYINPUT102), .ZN(n642) );
  NOR2_X1 U386 ( .A1(n592), .A2(n579), .ZN(n586) );
  XNOR2_X1 U387 ( .A(n531), .B(n453), .ZN(n592) );
  BUF_X1 U388 ( .A(n470), .Z(n468) );
  XNOR2_X1 U389 ( .A(n505), .B(n463), .ZN(n713) );
  XNOR2_X1 U390 ( .A(G902), .B(KEYINPUT15), .ZN(n601) );
  NOR2_X1 U391 ( .A1(n537), .A2(n432), .ZN(n345) );
  XOR2_X1 U392 ( .A(G146), .B(G125), .Z(n469) );
  XNOR2_X1 U393 ( .A(n469), .B(n433), .ZN(n524) );
  INV_X1 U394 ( .A(KEYINPUT10), .ZN(n433) );
  AND2_X1 U395 ( .A1(n424), .A2(n451), .ZN(n604) );
  XNOR2_X1 U396 ( .A(n485), .B(n416), .ZN(n614) );
  XNOR2_X1 U397 ( .A(n491), .B(n484), .ZN(n416) );
  XNOR2_X1 U398 ( .A(n713), .B(G146), .ZN(n485) );
  NOR2_X1 U399 ( .A1(G953), .A2(G237), .ZN(n486) );
  XNOR2_X1 U400 ( .A(n389), .B(KEYINPUT71), .ZN(n388) );
  XOR2_X1 U401 ( .A(KEYINPUT18), .B(KEYINPUT73), .Z(n471) );
  XNOR2_X1 U402 ( .A(n450), .B(n471), .ZN(n449) );
  XNOR2_X1 U403 ( .A(n423), .B(G110), .ZN(n527) );
  INV_X1 U404 ( .A(G119), .ZN(n423) );
  XNOR2_X1 U405 ( .A(n525), .B(KEYINPUT85), .ZN(n380) );
  XNOR2_X1 U406 ( .A(n524), .B(n347), .ZN(n714) );
  INV_X1 U407 ( .A(G143), .ZN(n360) );
  OR2_X1 U408 ( .A1(G237), .A2(G902), .ZN(n481) );
  NOR2_X1 U409 ( .A1(n661), .A2(n587), .ZN(n588) );
  INV_X1 U410 ( .A(n579), .ZN(n443) );
  XNOR2_X1 U411 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n570) );
  INV_X1 U412 ( .A(KEYINPUT77), .ZN(n566) );
  XNOR2_X1 U413 ( .A(n393), .B(n391), .ZN(n458) );
  XNOR2_X1 U414 ( .A(n415), .B(KEYINPUT79), .ZN(n411) );
  NAND2_X1 U415 ( .A1(n604), .A2(KEYINPUT2), .ZN(n415) );
  INV_X1 U416 ( .A(n367), .ZN(n563) );
  INV_X1 U417 ( .A(G472), .ZN(n438) );
  NOR2_X1 U418 ( .A1(n362), .A2(n574), .ZN(n549) );
  XNOR2_X1 U419 ( .A(n383), .B(KEYINPUT28), .ZN(n362) );
  NAND2_X1 U420 ( .A1(n384), .A2(n662), .ZN(n383) );
  INV_X1 U421 ( .A(n544), .ZN(n384) );
  XNOR2_X1 U422 ( .A(n506), .B(n428), .ZN(n552) );
  XNOR2_X1 U423 ( .A(KEYINPUT100), .B(G478), .ZN(n428) );
  NAND2_X1 U424 ( .A1(n400), .A2(n399), .ZN(n398) );
  NOR2_X1 U425 ( .A1(n574), .A2(KEYINPUT90), .ZN(n399) );
  INV_X1 U426 ( .A(n573), .ZN(n400) );
  XNOR2_X1 U427 ( .A(n662), .B(n437), .ZN(n596) );
  INV_X1 U428 ( .A(KEYINPUT6), .ZN(n437) );
  XNOR2_X1 U429 ( .A(n440), .B(n485), .ZN(n691) );
  XNOR2_X1 U430 ( .A(n468), .B(n466), .ZN(n440) );
  INV_X1 U431 ( .A(n374), .ZN(n370) );
  INV_X1 U432 ( .A(KEYINPUT48), .ZN(n425) );
  XNOR2_X1 U433 ( .A(KEYINPUT20), .B(KEYINPUT88), .ZN(n520) );
  XOR2_X1 U434 ( .A(KEYINPUT91), .B(G137), .Z(n488) );
  XOR2_X1 U435 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n483) );
  XNOR2_X1 U436 ( .A(G119), .B(G101), .ZN(n482) );
  XNOR2_X1 U437 ( .A(n419), .B(KEYINPUT3), .ZN(n489) );
  XNOR2_X1 U438 ( .A(G116), .B(G113), .ZN(n419) );
  XOR2_X1 U439 ( .A(KEYINPUT12), .B(G104), .Z(n455) );
  XNOR2_X1 U440 ( .A(G113), .B(G131), .ZN(n454) );
  XNOR2_X1 U441 ( .A(n394), .B(G140), .ZN(n393) );
  NAND2_X1 U442 ( .A1(n486), .A2(G214), .ZN(n394) );
  XNOR2_X1 U443 ( .A(n457), .B(n392), .ZN(n391) );
  XNOR2_X1 U444 ( .A(G143), .B(G122), .ZN(n457) );
  XNOR2_X1 U445 ( .A(KEYINPUT94), .B(KEYINPUT11), .ZN(n392) );
  XNOR2_X1 U446 ( .A(G131), .B(KEYINPUT4), .ZN(n463) );
  XNOR2_X1 U447 ( .A(n450), .B(n471), .ZN(n448) );
  INV_X1 U448 ( .A(n574), .ZN(n429) );
  XNOR2_X1 U449 ( .A(n538), .B(n361), .ZN(n539) );
  INV_X1 U450 ( .A(KEYINPUT30), .ZN(n361) );
  NAND2_X1 U451 ( .A1(n592), .A2(n385), .ZN(n544) );
  AND2_X1 U452 ( .A1(n653), .A2(n535), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n420), .B(n489), .ZN(n700) );
  XNOR2_X1 U454 ( .A(n527), .B(n421), .ZN(n420) );
  XNOR2_X1 U455 ( .A(n422), .B(G122), .ZN(n421) );
  INV_X1 U456 ( .A(KEYINPUT16), .ZN(n422) );
  XNOR2_X1 U457 ( .A(n378), .B(n377), .ZN(n618) );
  XNOR2_X1 U458 ( .A(n382), .B(n379), .ZN(n378) );
  XNOR2_X1 U459 ( .A(n381), .B(n380), .ZN(n379) );
  XNOR2_X1 U460 ( .A(KEYINPUT9), .B(KEYINPUT98), .ZN(n495) );
  XNOR2_X1 U461 ( .A(G116), .B(G122), .ZN(n493) );
  INV_X1 U462 ( .A(KEYINPUT2), .ZN(n375) );
  INV_X1 U463 ( .A(KEYINPUT39), .ZN(n430) );
  INV_X1 U464 ( .A(n596), .ZN(n587) );
  NAND2_X1 U465 ( .A1(n580), .A2(n443), .ZN(n442) );
  XNOR2_X1 U466 ( .A(n615), .B(n352), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n618), .B(KEYINPUT122), .ZN(n619) );
  XNOR2_X1 U468 ( .A(n545), .B(n366), .ZN(n724) );
  XNOR2_X1 U469 ( .A(KEYINPUT42), .B(KEYINPUT109), .ZN(n366) );
  NAND2_X1 U470 ( .A1(n387), .A2(n585), .ZN(n386) );
  XNOR2_X1 U471 ( .A(n533), .B(KEYINPUT36), .ZN(n387) );
  INV_X1 U472 ( .A(KEYINPUT35), .ZN(n434) );
  XNOR2_X1 U473 ( .A(n572), .B(n571), .ZN(n641) );
  NOR2_X1 U474 ( .A1(n573), .A2(n445), .ZN(n572) );
  NAND2_X1 U475 ( .A1(n585), .A2(n662), .ZN(n445) );
  NOR2_X1 U476 ( .A1(n547), .A2(n552), .ZN(n427) );
  NOR2_X2 U477 ( .A1(n396), .A2(n395), .ZN(n626) );
  NAND2_X1 U478 ( .A1(n398), .A2(n350), .ZN(n396) );
  XNOR2_X1 U479 ( .A(n694), .B(n404), .ZN(n697) );
  XNOR2_X1 U480 ( .A(n696), .B(n695), .ZN(n404) );
  XNOR2_X1 U481 ( .A(n607), .B(n353), .ZN(n403) );
  XNOR2_X1 U482 ( .A(n689), .B(n405), .ZN(n692) );
  XNOR2_X1 U483 ( .A(n691), .B(n690), .ZN(n405) );
  NAND2_X1 U484 ( .A1(n407), .A2(n406), .ZN(n401) );
  XNOR2_X1 U485 ( .A(n479), .B(n480), .ZN(n346) );
  XNOR2_X1 U486 ( .A(G137), .B(G140), .ZN(n347) );
  AND2_X1 U487 ( .A1(n388), .A2(n386), .ZN(n348) );
  NAND2_X1 U488 ( .A1(n593), .A2(n575), .ZN(n349) );
  AND2_X1 U489 ( .A1(n397), .A2(n575), .ZN(n350) );
  XOR2_X1 U490 ( .A(n534), .B(KEYINPUT38), .Z(n351) );
  XOR2_X1 U491 ( .A(n614), .B(KEYINPUT62), .Z(n352) );
  XNOR2_X1 U492 ( .A(n507), .B(KEYINPUT59), .ZN(n353) );
  XOR2_X1 U493 ( .A(n603), .B(KEYINPUT65), .Z(n354) );
  XNOR2_X1 U494 ( .A(n611), .B(n610), .ZN(n355) );
  XNOR2_X1 U495 ( .A(KEYINPUT78), .B(KEYINPUT45), .ZN(n356) );
  NOR2_X1 U496 ( .A1(G952), .A2(n707), .ZN(n698) );
  INV_X1 U497 ( .A(n698), .ZN(n406) );
  XOR2_X1 U498 ( .A(n613), .B(KEYINPUT56), .Z(n357) );
  XOR2_X1 U499 ( .A(KEYINPUT60), .B(KEYINPUT66), .Z(n358) );
  XOR2_X1 U500 ( .A(n617), .B(n616), .Z(n359) );
  NAND2_X1 U501 ( .A1(n708), .A2(n411), .ZN(n605) );
  XNOR2_X2 U502 ( .A(n600), .B(n356), .ZN(n708) );
  XNOR2_X1 U503 ( .A(n612), .B(n355), .ZN(n407) );
  NAND2_X1 U504 ( .A1(n390), .A2(n729), .ZN(n389) );
  XNOR2_X1 U505 ( .A(n363), .B(n359), .ZN(G57) );
  NAND2_X1 U506 ( .A1(n402), .A2(n406), .ZN(n363) );
  XNOR2_X1 U507 ( .A(n364), .B(n358), .ZN(G60) );
  NAND2_X1 U508 ( .A1(n403), .A2(n406), .ZN(n364) );
  NAND2_X1 U509 ( .A1(n693), .A2(G217), .ZN(n620) );
  NAND2_X1 U510 ( .A1(n365), .A2(n708), .ZN(n409) );
  NAND2_X1 U511 ( .A1(n414), .A2(n348), .ZN(n426) );
  NAND2_X1 U512 ( .A1(n367), .A2(n668), .ZN(n444) );
  XNOR2_X2 U513 ( .A(n418), .B(n346), .ZN(n367) );
  AND2_X1 U514 ( .A1(n591), .A2(n367), .ZN(n553) );
  NAND2_X1 U515 ( .A1(n371), .A2(n368), .ZN(n594) );
  NAND2_X1 U516 ( .A1(n370), .A2(n369), .ZN(n368) );
  NOR2_X1 U517 ( .A1(n726), .A2(KEYINPUT44), .ZN(n369) );
  NAND2_X1 U518 ( .A1(n726), .A2(KEYINPUT44), .ZN(n372) );
  NAND2_X1 U519 ( .A1(n374), .A2(KEYINPUT44), .ZN(n373) );
  NAND2_X1 U520 ( .A1(n725), .A2(n630), .ZN(n374) );
  NAND2_X1 U521 ( .A1(n715), .A2(n708), .ZN(n376) );
  AND2_X1 U522 ( .A1(n376), .A2(n375), .ZN(n650) );
  INV_X1 U523 ( .A(n714), .ZN(n377) );
  XNOR2_X1 U524 ( .A(n527), .B(n526), .ZN(n381) );
  NAND2_X1 U525 ( .A1(n523), .A2(G221), .ZN(n382) );
  XNOR2_X1 U526 ( .A(n500), .B(n501), .ZN(n523) );
  INV_X1 U527 ( .A(n662), .ZN(n575) );
  XNOR2_X2 U528 ( .A(n492), .B(n438), .ZN(n662) );
  INV_X1 U529 ( .A(n386), .ZN(n644) );
  XNOR2_X1 U530 ( .A(n550), .B(KEYINPUT47), .ZN(n390) );
  AND2_X1 U531 ( .A1(n573), .A2(KEYINPUT90), .ZN(n395) );
  NAND2_X1 U532 ( .A1(n574), .A2(KEYINPUT90), .ZN(n397) );
  XNOR2_X1 U533 ( .A(n401), .B(n357), .ZN(G51) );
  XNOR2_X1 U534 ( .A(n548), .B(KEYINPUT19), .ZN(n569) );
  XNOR2_X1 U535 ( .A(n408), .B(n622), .ZN(G66) );
  NOR2_X2 U536 ( .A1(n621), .A2(n698), .ZN(n408) );
  INV_X1 U537 ( .A(n601), .ZN(n410) );
  INV_X1 U538 ( .A(n605), .ZN(n651) );
  XNOR2_X1 U539 ( .A(n412), .B(KEYINPUT104), .ZN(n413) );
  NOR2_X1 U540 ( .A1(n576), .A2(n672), .ZN(n412) );
  NOR2_X1 U541 ( .A1(n626), .A2(n641), .ZN(n576) );
  XNOR2_X2 U542 ( .A(n444), .B(KEYINPUT80), .ZN(n548) );
  NOR2_X1 U543 ( .A1(n594), .A2(n413), .ZN(n599) );
  NAND2_X1 U544 ( .A1(n611), .A2(n601), .ZN(n418) );
  XNOR2_X1 U545 ( .A(n478), .B(n477), .ZN(n611) );
  XNOR2_X1 U546 ( .A(n426), .B(n425), .ZN(n424) );
  XNOR2_X1 U547 ( .A(n546), .B(KEYINPUT46), .ZN(n414) );
  NAND2_X1 U548 ( .A1(n554), .A2(n541), .ZN(n431) );
  NOR2_X1 U549 ( .A1(n724), .A2(n727), .ZN(n546) );
  XNOR2_X2 U550 ( .A(n417), .B(n570), .ZN(n589) );
  AND2_X2 U551 ( .A1(n569), .A2(n568), .ZN(n417) );
  INV_X1 U552 ( .A(n586), .ZN(n656) );
  NAND2_X1 U553 ( .A1(n539), .A2(n535), .ZN(n432) );
  XNOR2_X2 U554 ( .A(n435), .B(n434), .ZN(n725) );
  XNOR2_X1 U555 ( .A(n590), .B(KEYINPUT34), .ZN(n436) );
  XNOR2_X2 U556 ( .A(n574), .B(n439), .ZN(n585) );
  INV_X1 U557 ( .A(KEYINPUT1), .ZN(n439) );
  XNOR2_X2 U558 ( .A(n467), .B(G469), .ZN(n574) );
  NOR2_X2 U559 ( .A1(n595), .A2(n582), .ZN(n584) );
  XNOR2_X2 U560 ( .A(n441), .B(n581), .ZN(n595) );
  OR2_X2 U561 ( .A1(n589), .A2(n442), .ZN(n441) );
  NAND2_X1 U562 ( .A1(n447), .A2(n446), .ZN(n476) );
  NAND2_X1 U563 ( .A1(n470), .A2(n448), .ZN(n446) );
  OR2_X2 U564 ( .A1(n470), .A2(n449), .ZN(n447) );
  INV_X1 U565 ( .A(n469), .ZN(n450) );
  BUF_X1 U566 ( .A(n699), .Z(n701) );
  AND2_X1 U567 ( .A1(n565), .A2(n647), .ZN(n451) );
  AND2_X1 U568 ( .A1(G953), .A2(G898), .ZN(n452) );
  XOR2_X1 U569 ( .A(n530), .B(n529), .Z(n453) );
  INV_X1 U570 ( .A(n728), .ZN(n565) );
  NOR2_X1 U571 ( .A1(n567), .A2(n452), .ZN(n568) );
  XNOR2_X1 U572 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U573 ( .A(KEYINPUT22), .B(KEYINPUT64), .ZN(n581) );
  XNOR2_X1 U574 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U575 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U576 ( .A(n524), .B(n456), .ZN(n459) );
  XNOR2_X1 U577 ( .A(n459), .B(n458), .ZN(n507) );
  XNOR2_X2 U578 ( .A(G104), .B(KEYINPUT83), .ZN(n460) );
  INV_X1 U579 ( .A(n460), .ZN(n462) );
  XNOR2_X1 U580 ( .A(G101), .B(G107), .ZN(n461) );
  XNOR2_X1 U581 ( .A(n462), .B(n461), .ZN(n699) );
  XNOR2_X1 U582 ( .A(n699), .B(KEYINPUT70), .ZN(n470) );
  XNOR2_X1 U583 ( .A(G110), .B(n347), .ZN(n465) );
  NAND2_X1 U584 ( .A1(G227), .A2(n707), .ZN(n464) );
  XNOR2_X1 U585 ( .A(n465), .B(n464), .ZN(n466) );
  INV_X1 U586 ( .A(n585), .ZN(n655) );
  XOR2_X1 U587 ( .A(n472), .B(KEYINPUT17), .Z(n474) );
  NAND2_X1 U588 ( .A1(G224), .A2(n707), .ZN(n473) );
  XNOR2_X1 U589 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U590 ( .A(n476), .B(n475), .ZN(n478) );
  XOR2_X1 U591 ( .A(KEYINPUT4), .B(n700), .Z(n477) );
  NAND2_X1 U592 ( .A1(G210), .A2(n481), .ZN(n479) );
  INV_X1 U593 ( .A(KEYINPUT84), .ZN(n480) );
  NAND2_X1 U594 ( .A1(G214), .A2(n481), .ZN(n668) );
  XNOR2_X1 U595 ( .A(n483), .B(n482), .ZN(n484) );
  NAND2_X1 U596 ( .A1(n486), .A2(G210), .ZN(n487) );
  XNOR2_X1 U597 ( .A(n488), .B(n487), .ZN(n490) );
  NOR2_X1 U598 ( .A1(n614), .A2(G902), .ZN(n492) );
  XOR2_X1 U599 ( .A(KEYINPUT97), .B(G107), .Z(n494) );
  XNOR2_X1 U600 ( .A(n494), .B(n493), .ZN(n498) );
  XOR2_X1 U601 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n496) );
  XNOR2_X1 U602 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U603 ( .A(n498), .B(n497), .Z(n503) );
  NAND2_X1 U604 ( .A1(n707), .A2(G234), .ZN(n501) );
  XNOR2_X1 U605 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n499) );
  XNOR2_X1 U606 ( .A(n499), .B(KEYINPUT68), .ZN(n500) );
  NAND2_X1 U607 ( .A1(n523), .A2(G217), .ZN(n502) );
  XNOR2_X1 U608 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U609 ( .A(n505), .B(n504), .ZN(n696) );
  NOR2_X1 U610 ( .A1(G902), .A2(n696), .ZN(n506) );
  NOR2_X1 U611 ( .A1(n507), .A2(G902), .ZN(n511) );
  XOR2_X1 U612 ( .A(KEYINPUT96), .B(KEYINPUT13), .Z(n509) );
  XNOR2_X1 U613 ( .A(KEYINPUT95), .B(G475), .ZN(n508) );
  XNOR2_X1 U614 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U615 ( .A(n511), .B(n510), .Z(n551) );
  INV_X1 U616 ( .A(n551), .ZN(n547) );
  NAND2_X1 U617 ( .A1(n552), .A2(n547), .ZN(n512) );
  XOR2_X1 U618 ( .A(KEYINPUT101), .B(n512), .Z(n636) );
  NAND2_X1 U619 ( .A1(G234), .A2(G237), .ZN(n513) );
  XNOR2_X1 U620 ( .A(n513), .B(KEYINPUT14), .ZN(n680) );
  NOR2_X1 U621 ( .A1(G902), .A2(n707), .ZN(n515) );
  NOR2_X1 U622 ( .A1(G953), .A2(G952), .ZN(n514) );
  NOR2_X1 U623 ( .A1(n515), .A2(n514), .ZN(n516) );
  NAND2_X1 U624 ( .A1(n680), .A2(n516), .ZN(n567) );
  INV_X1 U625 ( .A(n567), .ZN(n518) );
  NAND2_X1 U626 ( .A1(G953), .A2(G900), .ZN(n517) );
  NAND2_X1 U627 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U628 ( .A(KEYINPUT75), .B(n519), .ZN(n535) );
  NAND2_X1 U629 ( .A1(n601), .A2(G234), .ZN(n521) );
  XNOR2_X1 U630 ( .A(n521), .B(n520), .ZN(n528) );
  NAND2_X1 U631 ( .A1(n528), .A2(G221), .ZN(n522) );
  XOR2_X1 U632 ( .A(KEYINPUT21), .B(n522), .Z(n653) );
  XOR2_X1 U633 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n526) );
  XNOR2_X1 U634 ( .A(G128), .B(KEYINPUT24), .ZN(n525) );
  NOR2_X1 U635 ( .A1(n618), .A2(G902), .ZN(n531) );
  XOR2_X1 U636 ( .A(KEYINPUT87), .B(KEYINPUT25), .Z(n530) );
  NAND2_X1 U637 ( .A1(G217), .A2(n528), .ZN(n529) );
  NOR2_X1 U638 ( .A1(n636), .A2(n544), .ZN(n532) );
  NAND2_X1 U639 ( .A1(n596), .A2(n532), .ZN(n559) );
  NOR2_X1 U640 ( .A1(n548), .A2(n559), .ZN(n533) );
  INV_X1 U641 ( .A(KEYINPUT72), .ZN(n534) );
  XNOR2_X1 U642 ( .A(KEYINPUT89), .B(n653), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n668), .A2(n662), .ZN(n538) );
  NOR2_X1 U644 ( .A1(n556), .A2(n636), .ZN(n540) );
  XNOR2_X1 U645 ( .A(n540), .B(KEYINPUT40), .ZN(n727) );
  NAND2_X1 U646 ( .A1(n552), .A2(n551), .ZN(n670) );
  NAND2_X1 U647 ( .A1(n541), .A2(n668), .ZN(n671) );
  XNOR2_X1 U648 ( .A(KEYINPUT41), .B(n542), .ZN(n543) );
  INV_X1 U649 ( .A(n543), .ZN(n666) );
  NAND2_X1 U650 ( .A1(n666), .A2(n549), .ZN(n545) );
  XNOR2_X1 U651 ( .A(KEYINPUT103), .B(n642), .ZN(n557) );
  AND2_X1 U652 ( .A1(n636), .A2(n557), .ZN(n672) );
  NAND2_X1 U653 ( .A1(n549), .A2(n569), .ZN(n635) );
  NOR2_X1 U654 ( .A1(n672), .A2(n635), .ZN(n550) );
  NOR2_X1 U655 ( .A1(n552), .A2(n551), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n345), .A2(n553), .ZN(n555) );
  XNOR2_X1 U657 ( .A(KEYINPUT108), .B(n555), .ZN(n729) );
  NOR2_X1 U658 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U659 ( .A(n558), .B(KEYINPUT110), .ZN(n728) );
  NOR2_X1 U660 ( .A1(n585), .A2(n559), .ZN(n560) );
  NAND2_X1 U661 ( .A1(n668), .A2(n560), .ZN(n561) );
  XNOR2_X1 U662 ( .A(n561), .B(KEYINPUT106), .ZN(n562) );
  XNOR2_X1 U663 ( .A(KEYINPUT43), .B(n562), .ZN(n564) );
  NAND2_X1 U664 ( .A1(n564), .A2(n563), .ZN(n647) );
  XNOR2_X2 U665 ( .A(n604), .B(n566), .ZN(n715) );
  XNOR2_X1 U666 ( .A(KEYINPUT93), .B(KEYINPUT31), .ZN(n571) );
  XNOR2_X1 U667 ( .A(KEYINPUT105), .B(n592), .ZN(n652) );
  INV_X1 U668 ( .A(n652), .ZN(n577) );
  AND2_X1 U669 ( .A1(n585), .A2(n577), .ZN(n578) );
  NAND2_X1 U670 ( .A1(n587), .A2(n578), .ZN(n582) );
  INV_X1 U671 ( .A(n670), .ZN(n580) );
  XNOR2_X1 U672 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n583) );
  XNOR2_X1 U673 ( .A(n588), .B(KEYINPUT33), .ZN(n648) );
  NOR2_X1 U674 ( .A1(n589), .A2(n648), .ZN(n590) );
  AND2_X1 U675 ( .A1(n592), .A2(n655), .ZN(n593) );
  OR2_X1 U676 ( .A1(n595), .A2(n349), .ZN(n630) );
  NOR2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n598) );
  AND2_X1 U678 ( .A1(n652), .A2(n655), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n623) );
  NAND2_X1 U680 ( .A1(n599), .A2(n623), .ZN(n600) );
  XOR2_X1 U681 ( .A(n601), .B(KEYINPUT76), .Z(n602) );
  NAND2_X1 U682 ( .A1(n602), .A2(KEYINPUT2), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n693), .A2(G475), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n693), .A2(G210), .ZN(n612) );
  XOR2_X1 U685 ( .A(KEYINPUT82), .B(KEYINPUT55), .Z(n609) );
  XNOR2_X1 U686 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n608) );
  XNOR2_X1 U687 ( .A(n609), .B(n608), .ZN(n610) );
  INV_X1 U688 ( .A(KEYINPUT119), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n693), .A2(G472), .ZN(n615) );
  XNOR2_X1 U690 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n617) );
  INV_X1 U691 ( .A(KEYINPUT81), .ZN(n616) );
  INV_X1 U692 ( .A(KEYINPUT123), .ZN(n622) );
  XNOR2_X1 U693 ( .A(G101), .B(KEYINPUT112), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n624), .B(n623), .ZN(G3) );
  INV_X1 U695 ( .A(n636), .ZN(n638) );
  NAND2_X1 U696 ( .A1(n626), .A2(n638), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n625), .B(G104), .ZN(G6) );
  XOR2_X1 U698 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n628) );
  NAND2_X1 U699 ( .A1(n626), .A2(n642), .ZN(n627) );
  XNOR2_X1 U700 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U701 ( .A(G107), .B(n629), .ZN(G9) );
  XNOR2_X1 U702 ( .A(G110), .B(n630), .ZN(G12) );
  INV_X1 U703 ( .A(n642), .ZN(n631) );
  NOR2_X1 U704 ( .A1(n631), .A2(n635), .ZN(n633) );
  XNOR2_X1 U705 ( .A(KEYINPUT113), .B(KEYINPUT29), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(n634) );
  XOR2_X1 U707 ( .A(G128), .B(n634), .Z(G30) );
  NOR2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U709 ( .A(G146), .B(n637), .Z(G48) );
  NAND2_X1 U710 ( .A1(n641), .A2(n638), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n639), .B(KEYINPUT114), .ZN(n640) );
  XNOR2_X1 U712 ( .A(G113), .B(n640), .ZN(G15) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n643), .B(G116), .ZN(G18) );
  XNOR2_X1 U715 ( .A(G125), .B(n644), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U717 ( .A(G140), .B(KEYINPUT115), .Z(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(G42) );
  NOR2_X1 U719 ( .A1(n648), .A2(n543), .ZN(n649) );
  NOR2_X1 U720 ( .A1(G953), .A2(n649), .ZN(n686) );
  NOR2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n684) );
  NOR2_X1 U722 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U723 ( .A(KEYINPUT49), .B(n654), .ZN(n659) );
  NAND2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(KEYINPUT50), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n575), .A2(n660), .ZN(n664) );
  NAND2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U730 ( .A(KEYINPUT51), .B(n665), .ZN(n667) );
  NAND2_X1 U731 ( .A1(n667), .A2(n666), .ZN(n678) );
  NOR2_X1 U732 ( .A1(n541), .A2(n668), .ZN(n669) );
  NOR2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U734 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U735 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n675), .A2(n648), .ZN(n676) );
  XOR2_X1 U737 ( .A(KEYINPUT116), .B(n676), .Z(n677) );
  NAND2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U739 ( .A(KEYINPUT52), .B(n679), .Z(n682) );
  NAND2_X1 U740 ( .A1(n680), .A2(G952), .ZN(n681) );
  NOR2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U743 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U744 ( .A(n687), .B(KEYINPUT53), .ZN(n688) );
  XNOR2_X1 U745 ( .A(KEYINPUT117), .B(n688), .ZN(G75) );
  XOR2_X1 U746 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n690) );
  NAND2_X1 U747 ( .A1(n693), .A2(G469), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n698), .A2(n692), .ZN(G54) );
  XOR2_X1 U749 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n695) );
  NAND2_X1 U750 ( .A1(n693), .A2(G478), .ZN(n694) );
  NOR2_X1 U751 ( .A1(n698), .A2(n697), .ZN(G63) );
  XNOR2_X1 U752 ( .A(n701), .B(n700), .ZN(n703) );
  NOR2_X1 U753 ( .A1(n707), .A2(G898), .ZN(n702) );
  NOR2_X1 U754 ( .A1(n703), .A2(n702), .ZN(n712) );
  NAND2_X1 U755 ( .A1(G953), .A2(G224), .ZN(n704) );
  XNOR2_X1 U756 ( .A(KEYINPUT61), .B(n704), .ZN(n705) );
  NAND2_X1 U757 ( .A1(n705), .A2(G898), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n706), .B(KEYINPUT124), .ZN(n710) );
  NAND2_X1 U759 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U760 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U761 ( .A(n712), .B(n711), .ZN(G69) );
  XNOR2_X1 U762 ( .A(n714), .B(n713), .ZN(n718) );
  XNOR2_X1 U763 ( .A(n718), .B(n715), .ZN(n716) );
  NOR2_X1 U764 ( .A1(G953), .A2(n716), .ZN(n717) );
  XNOR2_X1 U765 ( .A(n717), .B(KEYINPUT125), .ZN(n722) );
  XNOR2_X1 U766 ( .A(G227), .B(n718), .ZN(n719) );
  NAND2_X1 U767 ( .A1(n719), .A2(G900), .ZN(n720) );
  NAND2_X1 U768 ( .A1(n720), .A2(G953), .ZN(n721) );
  NAND2_X1 U769 ( .A1(n722), .A2(n721), .ZN(G72) );
  XOR2_X1 U770 ( .A(G137), .B(KEYINPUT126), .Z(n723) );
  XNOR2_X1 U771 ( .A(n724), .B(n723), .ZN(G39) );
  XNOR2_X1 U772 ( .A(G122), .B(n725), .ZN(G24) );
  XOR2_X1 U773 ( .A(n726), .B(G119), .Z(G21) );
  XOR2_X1 U774 ( .A(n727), .B(G131), .Z(G33) );
  XOR2_X1 U775 ( .A(G134), .B(n728), .Z(G36) );
  XNOR2_X1 U776 ( .A(G143), .B(n729), .ZN(G45) );
endmodule

