//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT24), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT23), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT65), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT23), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n208), .A2(new_n212), .A3(KEYINPUT64), .A4(new_n209), .ZN(new_n224));
  INV_X1    g023(.A(new_n220), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n215), .A2(new_n223), .A3(new_n224), .A4(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n206), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n207), .A3(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n211), .A3(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n235), .A2(new_n209), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n228), .A2(KEYINPUT25), .A3(new_n218), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n240), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n238), .A3(new_n209), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n231), .A2(new_n241), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G120gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G113gat), .ZN(new_n248));
  INV_X1    g047(.A(G113gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G120gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n252));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G134gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G127gat), .ZN(new_n257));
  INV_X1    g056(.A(G127gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G134gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n252), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G120gat), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(KEYINPUT1), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n255), .A2(new_n263), .A3(KEYINPUT73), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT73), .B1(new_n255), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT70), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n226), .B1(new_n267), .B2(KEYINPUT70), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT71), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n267), .A2(KEYINPUT70), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n268), .A4(new_n226), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n271), .B(new_n274), .C1(KEYINPUT26), .C2(new_n225), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT27), .B(G183gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(KEYINPUT28), .A3(new_n211), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n236), .A2(KEYINPUT27), .A3(new_n237), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n210), .B2(KEYINPUT27), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT27), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n211), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n277), .B1(new_n284), .B2(KEYINPUT28), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n275), .A2(new_n285), .A3(new_n206), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n246), .A2(new_n266), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n266), .B1(new_n246), .B2(new_n286), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n205), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT34), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n287), .A2(new_n288), .A3(new_n205), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n246), .A2(new_n286), .ZN(new_n296));
  INV_X1    g095(.A(new_n266), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n246), .A2(new_n286), .A3(new_n266), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n204), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(KEYINPUT74), .A3(KEYINPUT32), .ZN(new_n301));
  XNOR2_X1  g100(.A(G15gat), .B(G43gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G71gat), .B(G99gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT33), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n295), .A2(new_n301), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT75), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n295), .A2(new_n306), .A3(new_n309), .A4(new_n301), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n300), .A2(KEYINPUT32), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n304), .A2(new_n305), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n291), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  AOI211_X1 g115(.A(new_n314), .B(new_n290), .C1(new_n308), .C2(new_n310), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT5), .ZN(new_n319));
  NOR2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT2), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n326));
  INV_X1    g125(.A(G141gat), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(G148gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n324), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n323), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(new_n320), .ZN(new_n333));
  XNOR2_X1  g132(.A(G141gat), .B(G148gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(KEYINPUT2), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n255), .A2(new_n263), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n331), .A2(new_n335), .A3(new_n255), .A4(new_n263), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n319), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n339), .A2(KEYINPUT4), .ZN(new_n344));
  OR2_X1    g143(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(G141gat), .A3(new_n346), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n347), .A2(new_n329), .B1(new_n323), .B2(new_n322), .ZN(new_n348));
  XNOR2_X1  g147(.A(G155gat), .B(G162gat), .ZN(new_n349));
  INV_X1    g148(.A(G148gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n329), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n349), .B1(new_n321), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n264), .B2(new_n265), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n344), .B1(new_n355), .B2(KEYINPUT4), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT3), .B1(new_n348), .B2(new_n353), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n325), .A2(new_n326), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n330), .B1(new_n359), .B2(G141gat), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n332), .B1(new_n321), .B2(new_n320), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n335), .B(new_n358), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(new_n362), .A3(new_n337), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n341), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n343), .B1(new_n356), .B2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G1gat), .B(G29gat), .Z(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n339), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(new_n355), .B2(new_n371), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n363), .A2(new_n319), .A3(new_n341), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n365), .A2(KEYINPUT82), .A3(new_n370), .A4(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT6), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n370), .ZN(new_n379));
  INV_X1    g178(.A(new_n365), .ZN(new_n380));
  INV_X1    g179(.A(new_n375), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n355), .A2(KEYINPUT4), .ZN(new_n383));
  INV_X1    g182(.A(new_n344), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n364), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n343), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n370), .B(new_n375), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n378), .A2(new_n382), .A3(new_n389), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n382), .A2(new_n377), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT78), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n296), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G226gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(new_n203), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n246), .A2(new_n286), .A3(KEYINPUT78), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n400), .A2(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n296), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT76), .B(G197gat), .ZN(new_n406));
  INV_X1    g205(.A(G204gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G211gat), .B(G218gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT77), .B(G211gat), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT22), .B1(new_n411), .B2(G218gat), .ZN(new_n412));
  OR3_X1    g211(.A1(new_n408), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n410), .B1(new_n408), .B2(new_n412), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n405), .A2(new_n416), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n246), .A2(KEYINPUT78), .A3(new_n286), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT78), .B1(new_n246), .B2(new_n286), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n403), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n296), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n400), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n415), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n396), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT79), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n417), .A2(new_n423), .A3(new_n396), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT30), .B1(new_n424), .B2(KEYINPUT79), .ZN(new_n430));
  AND4_X1   g229(.A1(new_n392), .A2(new_n428), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G78gat), .B(G106gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(G22gat), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G228gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(new_n203), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n362), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n413), .B(new_n414), .C1(KEYINPUT29), .C2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n414), .A2(KEYINPUT83), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(KEYINPUT29), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n413), .A2(KEYINPUT83), .A3(new_n414), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT3), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n437), .B(new_n439), .C1(new_n443), .C2(new_n354), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT29), .B1(new_n413), .B2(new_n414), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n336), .B1(new_n445), .B2(KEYINPUT3), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n439), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n436), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT31), .B(G50gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n444), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n444), .B2(new_n448), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n434), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n444), .A2(new_n448), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n449), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n433), .A3(new_n451), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n318), .A2(new_n431), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n365), .A2(KEYINPUT86), .A3(new_n375), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT86), .B1(new_n365), .B2(new_n375), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n463), .A2(new_n464), .A3(new_n370), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n389), .A2(new_n377), .A3(new_n376), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT87), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n464), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(new_n379), .A3(new_n462), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n389), .A4(new_n378), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n467), .A2(new_n391), .A3(new_n471), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n461), .A2(new_n472), .A3(KEYINPUT35), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n316), .A2(new_n317), .A3(new_n458), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n460), .A2(KEYINPUT35), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT40), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n341), .B1(new_n373), .B2(new_n363), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n338), .A2(new_n341), .A3(new_n339), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n478), .A2(KEYINPUT85), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT39), .ZN(new_n480));
  AOI211_X1 g279(.A(new_n477), .B(new_n480), .C1(KEYINPUT85), .C2(new_n478), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n370), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n476), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n469), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n481), .A2(new_n476), .A3(new_n484), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n458), .B1(new_n461), .B2(new_n488), .ZN(new_n489));
  AND4_X1   g288(.A1(new_n391), .A2(new_n467), .A3(new_n425), .A4(new_n471), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT91), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n492));
  INV_X1    g291(.A(new_n400), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n418), .A2(new_n419), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n404), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n415), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT89), .A4(new_n416), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n420), .A2(new_n422), .A3(new_n416), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT89), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n405), .A2(KEYINPUT88), .A3(new_n415), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n498), .A2(new_n499), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n492), .B1(new_n504), .B2(KEYINPUT37), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n492), .A3(KEYINPUT37), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n396), .A2(KEYINPUT37), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT38), .B1(new_n429), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n490), .B(new_n491), .C1(new_n505), .C2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT38), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n429), .A2(new_n507), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n417), .A2(KEYINPUT37), .A3(new_n423), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT92), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n505), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n506), .A3(new_n508), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n491), .B1(new_n518), .B2(new_n490), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n489), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n311), .A2(new_n315), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n290), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n311), .A2(new_n315), .A3(new_n291), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT36), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n316), .A2(new_n317), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT84), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n452), .A2(new_n434), .A3(new_n453), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n433), .B1(new_n456), .B2(new_n451), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n454), .A2(KEYINPUT84), .A3(new_n457), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OAI22_X1  g332(.A1(new_n524), .A2(new_n526), .B1(new_n533), .B2(new_n431), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n475), .B1(new_n520), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(G43gat), .A2(G50gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(G43gat), .A2(G50gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT95), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT95), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n540), .A2(KEYINPUT15), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G29gat), .ZN(new_n544));
  INV_X1    g343(.A(G36gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT14), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(G29gat), .B2(G36gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G29gat), .A2(G36gat), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n550), .B(new_n551), .C1(KEYINPUT15), .C2(new_n539), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n543), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(KEYINPUT96), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT96), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n546), .A2(new_n548), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n556), .A3(new_n551), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n543), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT97), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT97), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n553), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G15gat), .B(G22gat), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n563), .A2(G1gat), .ZN(new_n564));
  INV_X1    g363(.A(G8gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT16), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n563), .B1(new_n566), .B2(G1gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n565), .B1(new_n564), .B2(new_n567), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n543), .A2(new_n560), .A3(new_n557), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n560), .B1(new_n543), .B2(new_n557), .ZN(new_n574));
  OAI22_X1  g373(.A1(new_n573), .A2(new_n574), .B1(new_n543), .B2(new_n552), .ZN(new_n575));
  INV_X1    g374(.A(new_n571), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT13), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT99), .B1(new_n569), .B2(new_n570), .ZN(new_n582));
  INV_X1    g381(.A(new_n570), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n568), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(KEYINPUT17), .B2(new_n562), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n562), .A2(new_n588), .A3(KEYINPUT17), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT98), .B1(new_n575), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n587), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n592), .A2(new_n579), .A3(new_n577), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT18), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n581), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n588), .B1(new_n562), .B2(KEYINPUT17), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n575), .A2(KEYINPUT98), .A3(new_n590), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n598), .A2(new_n587), .B1(new_n575), .B2(new_n576), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT18), .B1(new_n599), .B2(new_n579), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT94), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G113gat), .B(G141gat), .Z(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G169gat), .B(G197gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g408(.A(KEYINPUT94), .B(new_n607), .C1(new_n595), .C2(new_n600), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n536), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(G71gat), .A2(G78gat), .ZN(new_n614));
  XOR2_X1   g413(.A(G57gat), .B(G64gat), .Z(new_n615));
  AOI211_X1 g414(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(KEYINPUT9), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n613), .B1(KEYINPUT9), .B2(new_n614), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT100), .B(G57gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(G64gat), .ZN(new_n619));
  INV_X1    g418(.A(G64gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(G57gat), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n617), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n576), .B1(KEYINPUT21), .B2(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT102), .Z(new_n625));
  NOR2_X1   g424(.A1(new_n623), .A2(KEYINPUT21), .ZN(new_n626));
  XOR2_X1   g425(.A(G127gat), .B(G155gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n625), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT101), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G183gat), .B(G211gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n629), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT7), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(KEYINPUT105), .A2(KEYINPUT7), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G85gat), .A2(G92gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n637), .A2(new_n638), .B1(G85gat), .B2(G92gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(KEYINPUT106), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n642), .B1(new_n639), .B2(new_n640), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n648), .B1(new_n649), .B2(new_n645), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(G99gat), .A2(G106gat), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT8), .ZN(new_n653));
  OAI22_X1  g452(.A1(new_n652), .A2(new_n653), .B1(G85gat), .B2(G92gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(G99gat), .A2(G106gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n651), .A2(new_n660), .A3(new_n655), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n623), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(new_n651), .B2(new_n655), .ZN(new_n663));
  AOI211_X1 g462(.A(new_n658), .B(new_n654), .C1(new_n647), .C2(new_n650), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n663), .A2(new_n664), .B1(new_n622), .B2(new_n616), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT10), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n662), .A2(new_n665), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n659), .A2(KEYINPUT10), .A3(new_n623), .A4(new_n661), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n674), .A3(new_n667), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n674), .B1(new_n673), .B2(new_n667), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n669), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n673), .A2(new_n667), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT107), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n673), .A2(new_n686), .A3(new_n667), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n682), .B1(new_n666), .B2(new_n668), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n659), .A2(new_n661), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n598), .B(new_n692), .C1(new_n590), .C2(new_n575), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n562), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g493(.A1(G232gat), .A2(G233gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT103), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n694), .B1(KEYINPUT41), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(G190gat), .B(G218gat), .Z(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n697), .A2(KEYINPUT41), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT104), .ZN(new_n703));
  XOR2_X1   g502(.A(G134gat), .B(G162gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n700), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n693), .A2(new_n707), .A3(new_n698), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n701), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n693), .A2(new_n707), .A3(new_n698), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n707), .B1(new_n693), .B2(new_n698), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n705), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n636), .A2(new_n691), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n612), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n392), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(G1gat), .Z(G1324gat));
  NAND3_X1  g515(.A1(new_n612), .A2(new_n461), .A3(new_n713), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT110), .B(KEYINPUT16), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G8gat), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT109), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n717), .A2(G8gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(KEYINPUT42), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(G1325gat));
  NOR2_X1   g524(.A1(new_n524), .A2(new_n526), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G15gat), .B1(new_n714), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(G15gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n318), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n714), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT111), .ZN(G1326gat));
  NOR2_X1   g531(.A1(new_n714), .A2(new_n533), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT43), .B(G22gat), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1327gat));
  NAND2_X1  g534(.A1(new_n712), .A2(new_n709), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n636), .A2(new_n737), .A3(new_n690), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n612), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n390), .A2(new_n391), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n544), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n739), .A2(KEYINPUT112), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT112), .B1(new_n739), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n536), .B2(new_n737), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n509), .A2(new_n505), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n467), .A2(new_n471), .A3(new_n391), .A4(new_n425), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT91), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(new_n510), .A3(new_n515), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n534), .B1(new_n752), .B2(new_n489), .ZN(new_n753));
  OAI211_X1 g552(.A(KEYINPUT44), .B(new_n736), .C1(new_n753), .C2(new_n475), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n690), .B(KEYINPUT113), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n756), .A2(new_n611), .A3(new_n636), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n740), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G29gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n742), .A2(KEYINPUT45), .A3(new_n743), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n746), .A2(new_n759), .A3(new_n760), .ZN(G1328gat));
  INV_X1    g560(.A(new_n461), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n739), .A2(G36gat), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT46), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n755), .A2(new_n461), .A3(new_n757), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G36gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1329gat));
  NAND4_X1  g566(.A1(new_n748), .A2(new_n726), .A3(new_n754), .A4(new_n757), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G43gat), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT47), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(G43gat), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n612), .A2(new_n772), .A3(new_n318), .A4(new_n738), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n769), .B(new_n773), .C1(new_n770), .C2(KEYINPUT47), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1330gat));
  NAND3_X1  g576(.A1(new_n755), .A2(new_n458), .A3(new_n757), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(G50gat), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n739), .A2(G50gat), .A3(new_n533), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT48), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n755), .A2(new_n532), .A3(new_n757), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n783), .B2(G50gat), .ZN(new_n784));
  OAI22_X1  g583(.A1(new_n779), .A2(new_n782), .B1(new_n784), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g584(.A1(new_n756), .A2(new_n611), .A3(new_n636), .A4(new_n737), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n536), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n740), .B(KEYINPUT115), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(new_n618), .ZN(G1332gat));
  NOR2_X1   g590(.A1(new_n788), .A2(new_n762), .ZN(new_n792));
  NOR2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  AND2_X1   g592(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n792), .B2(new_n793), .ZN(G1333gat));
  NAND2_X1  g595(.A1(new_n787), .A2(new_n726), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n316), .A2(new_n317), .A3(G71gat), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n797), .A2(G71gat), .B1(new_n787), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g599(.A1(new_n787), .A2(new_n532), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  INV_X1    g601(.A(new_n611), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n636), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n736), .B(new_n804), .C1(new_n753), .C2(new_n475), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n475), .ZN(new_n808));
  INV_X1    g607(.A(new_n489), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT92), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n514), .B(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n506), .A2(new_n508), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n750), .B1(new_n812), .B2(new_n517), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n491), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n809), .B1(new_n814), .B2(new_n751), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n808), .B1(new_n815), .B2(new_n534), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n816), .A2(KEYINPUT51), .A3(new_n736), .A4(new_n804), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n807), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(G85gat), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n740), .A4(new_n690), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n803), .A2(new_n636), .A3(new_n691), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n755), .A2(new_n740), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n822), .B2(new_n819), .ZN(G1336gat));
  INV_X1    g622(.A(new_n756), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(G92gat), .A3(new_n762), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n748), .A2(new_n461), .A3(new_n754), .A4(new_n821), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G92gat), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n826), .A2(new_n828), .A3(new_n829), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1337gat));
  INV_X1    g633(.A(G99gat), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n818), .A2(new_n835), .A3(new_n318), .A4(new_n690), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n755), .A2(new_n726), .A3(new_n821), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n835), .ZN(G1338gat));
  NAND4_X1  g637(.A1(new_n748), .A2(new_n532), .A3(new_n754), .A4(new_n821), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(G106gat), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n824), .A2(G106gat), .A3(new_n459), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT117), .Z(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n807), .B2(new_n817), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT53), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n818), .A2(new_n841), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n748), .A2(new_n458), .A3(new_n754), .A4(new_n821), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(G106gat), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n849));
  AND4_X1   g648(.A1(new_n845), .A2(new_n846), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT53), .B1(new_n818), .B2(new_n841), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n845), .B1(new_n851), .B2(new_n848), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n844), .B1(new_n850), .B2(new_n852), .ZN(G1339gat));
  AND4_X1   g652(.A1(new_n611), .A2(new_n636), .A3(new_n737), .A4(new_n691), .ZN(new_n854));
  INV_X1    g653(.A(new_n689), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n671), .A2(new_n668), .A3(new_n672), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n671), .A2(KEYINPUT119), .A3(new_n668), .A4(new_n672), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n860), .A2(new_n685), .A3(KEYINPUT54), .A4(new_n687), .ZN(new_n861));
  INV_X1    g660(.A(new_n677), .ZN(new_n862));
  XOR2_X1   g661(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n675), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n861), .A2(new_n682), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n855), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT55), .A4(new_n682), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n867), .A2(new_n609), .A3(new_n610), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n593), .A2(new_n594), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n599), .A2(KEYINPUT18), .A3(new_n579), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n581), .A4(new_n607), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n599), .A2(new_n579), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n578), .A2(new_n580), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n606), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n736), .B1(new_n877), .B2(new_n690), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n636), .B1(new_n869), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n872), .A2(new_n875), .A3(KEYINPUT121), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n881), .A2(new_n867), .A3(new_n882), .A4(new_n868), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n736), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n854), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n461), .A2(new_n392), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(new_n533), .A3(new_n318), .A4(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(new_n249), .A3(new_n611), .ZN(new_n889));
  INV_X1    g688(.A(new_n474), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n885), .A2(new_n890), .A3(new_n789), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(new_n762), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n803), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n889), .B1(new_n893), .B2(new_n249), .ZN(G1340gat));
  NOR3_X1   g693(.A1(new_n888), .A2(new_n247), .A3(new_n824), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n690), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n247), .ZN(G1341gat));
  NAND3_X1  g696(.A1(new_n892), .A2(new_n258), .A3(new_n636), .ZN(new_n898));
  INV_X1    g697(.A(new_n636), .ZN(new_n899));
  OAI21_X1  g698(.A(G127gat), .B1(new_n888), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1342gat));
  NAND4_X1  g700(.A1(new_n891), .A2(new_n256), .A3(new_n762), .A4(new_n736), .ZN(new_n902));
  XNOR2_X1  g701(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  OAI21_X1  g704(.A(G134gat), .B1(new_n888), .B2(new_n737), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G1343gat));
  INV_X1    g706(.A(new_n789), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n886), .A2(new_n458), .A3(new_n727), .A4(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n461), .ZN(new_n910));
  AOI21_X1  g709(.A(G141gat), .B1(new_n910), .B2(new_n803), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n879), .A2(new_n884), .ZN(new_n912));
  INV_X1    g711(.A(new_n854), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n459), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n726), .A2(new_n392), .A3(new_n461), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT57), .B1(new_n885), .B2(new_n533), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(new_n327), .A3(new_n611), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n911), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g721(.A1(new_n910), .A2(new_n359), .A3(new_n690), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n917), .A2(new_n690), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n915), .B1(new_n885), .B2(new_n533), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n926), .A2(KEYINPUT123), .B1(new_n914), .B2(KEYINPUT57), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n928), .B(new_n915), .C1(new_n885), .C2(new_n533), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n925), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n350), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n926), .A2(KEYINPUT123), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n914), .A2(KEYINPUT57), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n690), .A3(new_n917), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT124), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n924), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n919), .A2(new_n691), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(KEYINPUT59), .A3(new_n359), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n923), .B1(new_n938), .B2(new_n940), .ZN(G1345gat));
  OAI21_X1  g740(.A(G155gat), .B1(new_n919), .B2(new_n899), .ZN(new_n942));
  INV_X1    g741(.A(G155gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n910), .A2(new_n943), .A3(new_n636), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1346gat));
  OAI21_X1  g744(.A(G162gat), .B1(new_n919), .B2(new_n737), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n737), .A2(new_n461), .A3(G162gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n909), .B2(new_n947), .ZN(G1347gat));
  NOR4_X1   g747(.A1(new_n885), .A2(new_n740), .A3(new_n762), .A4(new_n890), .ZN(new_n949));
  AOI21_X1  g748(.A(G169gat), .B1(new_n949), .B2(new_n803), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n789), .A2(new_n461), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT125), .ZN(new_n952));
  AND4_X1   g751(.A1(new_n533), .A2(new_n886), .A3(new_n318), .A4(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n611), .A2(new_n216), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(G1348gat));
  NAND3_X1  g754(.A1(new_n949), .A2(new_n217), .A3(new_n690), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n953), .A2(new_n756), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n217), .ZN(G1349gat));
  NAND3_X1  g757(.A1(new_n949), .A2(new_n276), .A3(new_n636), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n953), .A2(new_n636), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n236), .A2(new_n237), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n211), .A3(new_n736), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n953), .A2(new_n736), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(G190gat), .ZN(new_n968));
  AOI211_X1 g767(.A(KEYINPUT61), .B(new_n211), .C1(new_n953), .C2(new_n736), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g771(.A(KEYINPUT126), .B(new_n965), .C1(new_n968), .C2(new_n969), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1351gat));
  NAND2_X1  g773(.A1(new_n935), .A2(KEYINPUT127), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n927), .A2(new_n976), .A3(new_n929), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n952), .A2(new_n727), .ZN(new_n978));
  INV_X1    g777(.A(G197gat), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n611), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n975), .A2(new_n977), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n885), .A2(new_n740), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n726), .A2(new_n459), .A3(new_n762), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n979), .B1(new_n985), .B2(new_n611), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n981), .A2(new_n986), .ZN(G1352gat));
  NAND3_X1  g786(.A1(new_n984), .A2(new_n407), .A3(new_n690), .ZN(new_n988));
  XOR2_X1   g787(.A(new_n988), .B(KEYINPUT62), .Z(new_n989));
  AND4_X1   g788(.A1(new_n756), .A2(new_n975), .A3(new_n977), .A4(new_n978), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n990), .B2(new_n407), .ZN(G1353gat));
  INV_X1    g790(.A(G211gat), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n978), .A2(new_n636), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n935), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT63), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n899), .A2(new_n411), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n985), .B2(new_n996), .ZN(G1354gat));
  INV_X1    g796(.A(G218gat), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n737), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n975), .A2(new_n977), .A3(new_n978), .A4(new_n999), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n998), .B1(new_n985), .B2(new_n737), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1355gat));
endmodule


