

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765;

  INV_X1 U372 ( .A(G125), .ZN(n422) );
  XNOR2_X1 U373 ( .A(KEYINPUT73), .B(G110), .ZN(n393) );
  NAND2_X1 U374 ( .A1(n536), .A2(n544), .ZN(n625) );
  XNOR2_X1 U375 ( .A(n422), .B(G146), .ZN(n469) );
  XNOR2_X1 U376 ( .A(n394), .B(n393), .ZN(n518) );
  INV_X1 U377 ( .A(G953), .ZN(n705) );
  NOR2_X1 U378 ( .A1(n544), .A2(n543), .ZN(n727) );
  AND2_X2 U379 ( .A1(n401), .A2(n668), .ZN(n399) );
  OR2_X2 U380 ( .A1(n686), .A2(n476), .ZN(n478) );
  NOR2_X2 U381 ( .A1(n552), .A2(n553), .ZN(n559) );
  NAND2_X1 U382 ( .A1(n699), .A2(n386), .ZN(n427) );
  NOR2_X2 U383 ( .A1(n434), .A2(n433), .ZN(n585) );
  INV_X1 U384 ( .A(n759), .ZN(n578) );
  INV_X1 U385 ( .A(n530), .ZN(n623) );
  XNOR2_X1 U386 ( .A(n469), .B(n421), .ZN(n748) );
  AND2_X1 U387 ( .A1(n375), .A2(n673), .ZN(n681) );
  AND2_X1 U388 ( .A1(n396), .A2(n599), .ZN(n395) );
  XNOR2_X1 U389 ( .A(n373), .B(n558), .ZN(n366) );
  NOR2_X2 U390 ( .A1(n758), .A2(n760), .ZN(n535) );
  OR2_X1 U391 ( .A1(n633), .A2(n416), .ZN(n415) );
  XNOR2_X1 U392 ( .A(n376), .B(n565), .ZN(n633) );
  NAND2_X1 U393 ( .A1(n352), .A2(n564), .ZN(n376) );
  AND2_X1 U394 ( .A1(n389), .A2(n388), .ZN(n387) );
  XNOR2_X1 U395 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U396 ( .A(G107), .B(G104), .ZN(n394) );
  XNOR2_X2 U397 ( .A(n521), .B(n520), .ZN(n371) );
  NAND2_X1 U398 ( .A1(G469), .A2(n386), .ZN(n385) );
  INV_X1 U399 ( .A(G146), .ZN(n486) );
  XNOR2_X1 U400 ( .A(n607), .B(KEYINPUT87), .ZN(n583) );
  NOR2_X1 U401 ( .A1(G953), .A2(G237), .ZN(n487) );
  AND2_X1 U402 ( .A1(n606), .A2(n525), .ZN(n638) );
  NOR2_X1 U403 ( .A1(n762), .A2(n424), .ZN(n423) );
  INV_X1 U404 ( .A(n746), .ZN(n424) );
  XNOR2_X1 U405 ( .A(n391), .B(n465), .ZN(n491) );
  XNOR2_X1 U406 ( .A(G116), .B(G113), .ZN(n465) );
  XNOR2_X1 U407 ( .A(n466), .B(n464), .ZN(n391) );
  INV_X1 U408 ( .A(G119), .ZN(n464) );
  XNOR2_X1 U409 ( .A(G128), .B(G137), .ZN(n496) );
  INV_X1 U410 ( .A(KEYINPUT92), .ZN(n497) );
  XNOR2_X1 U411 ( .A(G119), .B(G110), .ZN(n498) );
  XOR2_X1 U412 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n443) );
  XNOR2_X1 U413 ( .A(G140), .B(KEYINPUT10), .ZN(n421) );
  XNOR2_X1 U414 ( .A(G113), .B(G143), .ZN(n454) );
  XNOR2_X1 U415 ( .A(n560), .B(KEYINPUT43), .ZN(n383) );
  XNOR2_X1 U416 ( .A(n721), .B(KEYINPUT103), .ZN(n562) );
  INV_X1 U417 ( .A(KEYINPUT76), .ZN(n582) );
  BUF_X1 U418 ( .A(n561), .Z(n379) );
  INV_X1 U419 ( .A(KEYINPUT0), .ZN(n405) );
  XNOR2_X1 U420 ( .A(n420), .B(n419), .ZN(n606) );
  XNOR2_X1 U421 ( .A(n507), .B(n505), .ZN(n419) );
  OR2_X1 U422 ( .A1(n742), .A2(G902), .ZN(n420) );
  XNOR2_X1 U423 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n505) );
  AND2_X1 U424 ( .A1(n689), .A2(G953), .ZN(n745) );
  NOR2_X1 U425 ( .A1(n562), .A2(n727), .ZN(n627) );
  INV_X1 U426 ( .A(G137), .ZN(n482) );
  XOR2_X1 U427 ( .A(KEYINPUT69), .B(G134), .Z(n484) );
  NAND2_X1 U428 ( .A1(G234), .A2(G237), .ZN(n508) );
  AND2_X1 U429 ( .A1(n414), .A2(n413), .ZN(n412) );
  INV_X1 U430 ( .A(n577), .ZN(n413) );
  INV_X1 U431 ( .A(G237), .ZN(n477) );
  NAND2_X1 U432 ( .A1(n390), .A2(G902), .ZN(n388) );
  XNOR2_X1 U433 ( .A(G101), .B(KEYINPUT3), .ZN(n466) );
  XNOR2_X1 U434 ( .A(KEYINPUT67), .B(KEYINPUT4), .ZN(n472) );
  XNOR2_X1 U435 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n468) );
  OR2_X1 U436 ( .A1(n606), .A2(n425), .ZN(n550) );
  NAND2_X1 U437 ( .A1(n426), .A2(n529), .ZN(n425) );
  INV_X1 U438 ( .A(n635), .ZN(n426) );
  XNOR2_X1 U439 ( .A(n521), .B(n492), .ZN(n699) );
  XNOR2_X1 U440 ( .A(G116), .B(G107), .ZN(n446) );
  XOR2_X1 U441 ( .A(KEYINPUT7), .B(G122), .Z(n447) );
  NAND2_X1 U442 ( .A1(n441), .A2(n439), .ZN(n537) );
  NOR2_X1 U443 ( .A1(n593), .A2(n440), .ZN(n439) );
  INV_X1 U444 ( .A(n529), .ZN(n440) );
  XOR2_X1 U445 ( .A(n699), .B(KEYINPUT62), .Z(n700) );
  XNOR2_X1 U446 ( .A(n677), .B(n749), .ZN(n750) );
  XNOR2_X1 U447 ( .A(n392), .B(n491), .ZN(n711) );
  XNOR2_X1 U448 ( .A(n353), .B(n518), .ZN(n392) );
  XNOR2_X1 U449 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n463) );
  XNOR2_X1 U450 ( .A(n504), .B(n503), .ZN(n742) );
  XNOR2_X1 U451 ( .A(n369), .B(n367), .ZN(n694) );
  XNOR2_X1 U452 ( .A(n456), .B(n368), .ZN(n367) );
  XNOR2_X1 U453 ( .A(n459), .B(n748), .ZN(n369) );
  INV_X1 U454 ( .A(KEYINPUT108), .ZN(n380) );
  NAND2_X1 U455 ( .A1(n383), .A2(n382), .ZN(n381) );
  INV_X1 U456 ( .A(n379), .ZN(n382) );
  XNOR2_X1 U457 ( .A(KEYINPUT40), .B(n534), .ZN(n760) );
  XNOR2_X1 U458 ( .A(n374), .B(KEYINPUT113), .ZN(n763) );
  XNOR2_X1 U459 ( .A(n430), .B(n429), .ZN(n428) );
  INV_X1 U460 ( .A(KEYINPUT36), .ZN(n429) );
  INV_X1 U461 ( .A(KEYINPUT75), .ZN(n584) );
  NOR2_X1 U462 ( .A1(n634), .A2(n404), .ZN(n592) );
  XNOR2_X1 U463 ( .A(n370), .B(KEYINPUT102), .ZN(n721) );
  INV_X1 U464 ( .A(n721), .ZN(n730) );
  INV_X1 U465 ( .A(n593), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n400), .B(KEYINPUT106), .ZN(n668) );
  XNOR2_X1 U467 ( .A(n735), .B(n734), .ZN(n736) );
  AND2_X1 U468 ( .A1(n372), .A2(n410), .ZN(n351) );
  INV_X1 U469 ( .A(n762), .ZN(n436) );
  XNOR2_X1 U470 ( .A(n381), .B(n380), .ZN(n762) );
  AND2_X1 U471 ( .A1(n637), .A2(n638), .ZN(n352) );
  XOR2_X1 U472 ( .A(n463), .B(G122), .Z(n353) );
  INV_X1 U473 ( .A(G902), .ZN(n386) );
  INV_X1 U474 ( .A(n606), .ZN(n435) );
  XOR2_X1 U475 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n354) );
  AND2_X1 U476 ( .A1(n479), .A2(G210), .ZN(n355) );
  XOR2_X1 U477 ( .A(n580), .B(KEYINPUT105), .Z(n356) );
  AND2_X1 U478 ( .A1(n415), .A2(n412), .ZN(n357) );
  INV_X1 U479 ( .A(G469), .ZN(n390) );
  AND2_X1 U480 ( .A1(n436), .A2(n615), .ZN(n358) );
  INV_X1 U481 ( .A(n576), .ZN(n418) );
  NAND2_X1 U482 ( .A1(n357), .A2(n351), .ZN(n409) );
  NOR2_X1 U483 ( .A1(n625), .A2(n626), .ZN(n480) );
  XNOR2_X1 U484 ( .A(n604), .B(n582), .ZN(n433) );
  XOR2_X1 U485 ( .A(n427), .B(n493), .Z(n359) );
  NAND2_X1 U486 ( .A1(n428), .A2(n583), .ZN(n374) );
  NAND2_X1 U487 ( .A1(n583), .A2(n435), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n686), .B(n685), .ZN(n687) );
  AND2_X2 U489 ( .A1(n366), .A2(n423), .ZN(n677) );
  INV_X1 U490 ( .A(n578), .ZN(n360) );
  BUF_X1 U491 ( .A(n633), .Z(n361) );
  NAND2_X1 U492 ( .A1(n431), .A2(n484), .ZN(n364) );
  NAND2_X1 U493 ( .A1(n362), .A2(n363), .ZN(n365) );
  NAND2_X1 U494 ( .A1(n365), .A2(n364), .ZN(n437) );
  INV_X1 U495 ( .A(n431), .ZN(n362) );
  INV_X1 U496 ( .A(n484), .ZN(n363) );
  NAND2_X1 U497 ( .A1(n411), .A2(n409), .ZN(n759) );
  BUF_X1 U498 ( .A(n732), .Z(n741) );
  BUF_X1 U499 ( .A(n675), .Z(n706) );
  NAND2_X1 U500 ( .A1(n633), .A2(n576), .ZN(n372) );
  AND2_X1 U501 ( .A1(n372), .A2(n412), .ZN(n408) );
  NAND2_X1 U502 ( .A1(n366), .A2(n358), .ZN(n616) );
  NOR2_X1 U503 ( .A1(n694), .A2(G902), .ZN(n461) );
  XNOR2_X1 U504 ( .A(n483), .B(KEYINPUT12), .ZN(n368) );
  NAND2_X1 U505 ( .A1(n544), .A2(n543), .ZN(n370) );
  NAND2_X1 U506 ( .A1(n371), .A2(n390), .ZN(n389) );
  OR2_X1 U507 ( .A1(n371), .A2(n385), .ZN(n384) );
  XNOR2_X1 U508 ( .A(n371), .B(n733), .ZN(n734) );
  NAND2_X1 U509 ( .A1(n557), .A2(n378), .ZN(n373) );
  NAND2_X1 U510 ( .A1(n559), .A2(n379), .ZN(n430) );
  NAND2_X1 U511 ( .A1(n408), .A2(n415), .ZN(n407) );
  NAND2_X2 U512 ( .A1(n387), .A2(n384), .ZN(n554) );
  NAND2_X1 U513 ( .A1(n669), .A2(n677), .ZN(n375) );
  NAND2_X1 U514 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X2 U515 ( .A(n377), .B(KEYINPUT65), .ZN(n732) );
  NAND2_X1 U516 ( .A1(n683), .A2(n682), .ZN(n377) );
  NOR2_X1 U517 ( .A1(n537), .A2(n530), .ZN(n438) );
  XNOR2_X1 U518 ( .A(n535), .B(KEYINPUT46), .ZN(n378) );
  NAND2_X1 U519 ( .A1(n617), .A2(n706), .ZN(n682) );
  XNOR2_X1 U520 ( .A(KEYINPUT111), .B(n481), .ZN(n650) );
  XNOR2_X2 U521 ( .A(n554), .B(KEYINPUT1), .ZN(n607) );
  NAND2_X1 U522 ( .A1(n352), .A2(n644), .ZN(n634) );
  NAND2_X1 U523 ( .A1(n561), .A2(n622), .ZN(n541) );
  XNOR2_X1 U524 ( .A(n561), .B(KEYINPUT38), .ZN(n530) );
  XNOR2_X2 U525 ( .A(n478), .B(n355), .ZN(n561) );
  NAND2_X1 U526 ( .A1(n395), .A2(n399), .ZN(n611) );
  NAND2_X1 U527 ( .A1(n398), .A2(n397), .ZN(n396) );
  INV_X1 U528 ( .A(n432), .ZN(n397) );
  NAND2_X1 U529 ( .A1(n406), .A2(KEYINPUT66), .ZN(n398) );
  NAND2_X1 U530 ( .A1(n609), .A2(n608), .ZN(n400) );
  NAND2_X1 U531 ( .A1(n402), .A2(n603), .ZN(n401) );
  NAND2_X1 U532 ( .A1(n601), .A2(n600), .ZN(n402) );
  NAND2_X1 U533 ( .A1(n356), .A2(n417), .ZN(n581) );
  AND2_X1 U534 ( .A1(n417), .A2(n403), .ZN(n594) );
  OR2_X1 U535 ( .A1(n417), .A2(n418), .ZN(n414) );
  INV_X1 U536 ( .A(n417), .ZN(n404) );
  XNOR2_X2 U537 ( .A(n574), .B(n405), .ZN(n417) );
  NAND2_X1 U538 ( .A1(n578), .A2(n602), .ZN(n406) );
  NAND2_X1 U539 ( .A1(n407), .A2(KEYINPUT35), .ZN(n411) );
  INV_X1 U540 ( .A(KEYINPUT35), .ZN(n410) );
  NAND2_X1 U541 ( .A1(n417), .A2(n418), .ZN(n416) );
  NOR2_X1 U542 ( .A1(n604), .A2(n550), .ZN(n551) );
  XNOR2_X2 U543 ( .A(n549), .B(n548), .ZN(n604) );
  XNOR2_X2 U544 ( .A(n427), .B(n493), .ZN(n549) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n431) );
  XNOR2_X2 U546 ( .A(KEYINPUT68), .B(G131), .ZN(n483) );
  NAND2_X1 U547 ( .A1(n432), .A2(KEYINPUT66), .ZN(n601) );
  NAND2_X2 U548 ( .A1(n666), .A2(n665), .ZN(n432) );
  XNOR2_X2 U549 ( .A(n588), .B(KEYINPUT32), .ZN(n666) );
  INV_X1 U550 ( .A(n607), .ZN(n637) );
  INV_X1 U551 ( .A(n604), .ZN(n564) );
  XNOR2_X2 U552 ( .A(n747), .B(n486), .ZN(n521) );
  XNOR2_X2 U553 ( .A(n437), .B(n485), .ZN(n747) );
  XNOR2_X1 U554 ( .A(n438), .B(n533), .ZN(n563) );
  INV_X1 U555 ( .A(n528), .ZN(n441) );
  XNOR2_X2 U556 ( .A(n541), .B(KEYINPUT19), .ZN(n573) );
  INV_X1 U557 ( .A(n549), .ZN(n644) );
  XNOR2_X2 U558 ( .A(G475), .B(n462), .ZN(n544) );
  AND2_X1 U559 ( .A1(n556), .A2(n555), .ZN(n557) );
  INV_X1 U560 ( .A(KEYINPUT48), .ZN(n558) );
  INV_X1 U561 ( .A(n579), .ZN(n525) );
  XNOR2_X1 U562 ( .A(n471), .B(n470), .ZN(n474) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(n499) );
  INV_X1 U564 ( .A(KEYINPUT39), .ZN(n531) );
  XNOR2_X1 U565 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U566 ( .A(n737), .B(KEYINPUT124), .ZN(n738) );
  INV_X1 U567 ( .A(KEYINPUT121), .ZN(n662) );
  XNOR2_X1 U568 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U569 ( .A(n664), .B(n663), .ZN(G75) );
  XNOR2_X1 U570 ( .A(KEYINPUT101), .B(G478), .ZN(n453) );
  XOR2_X1 U571 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n445) );
  NAND2_X1 U572 ( .A1(G234), .A2(n705), .ZN(n442) );
  XNOR2_X1 U573 ( .A(n443), .B(n442), .ZN(n502) );
  NAND2_X1 U574 ( .A1(G217), .A2(n502), .ZN(n444) );
  XNOR2_X1 U575 ( .A(n445), .B(n444), .ZN(n451) );
  XNOR2_X1 U576 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U577 ( .A(G134), .B(n448), .ZN(n449) );
  XNOR2_X1 U578 ( .A(G143), .B(G128), .ZN(n473) );
  XNOR2_X1 U579 ( .A(n449), .B(n473), .ZN(n450) );
  XNOR2_X1 U580 ( .A(n451), .B(n450), .ZN(n737) );
  NOR2_X1 U581 ( .A1(G902), .A2(n737), .ZN(n452) );
  XOR2_X1 U582 ( .A(n453), .B(n452), .Z(n536) );
  XOR2_X1 U583 ( .A(G122), .B(G104), .Z(n455) );
  XNOR2_X1 U584 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U585 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n458) );
  NAND2_X1 U586 ( .A1(G214), .A2(n487), .ZN(n457) );
  XNOR2_X1 U587 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U588 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n460) );
  XNOR2_X1 U589 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U590 ( .A1(n705), .A2(G224), .ZN(n467) );
  XNOR2_X1 U591 ( .A(n467), .B(KEYINPUT89), .ZN(n471) );
  XNOR2_X1 U592 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U593 ( .A(n473), .B(n472), .ZN(n485) );
  XNOR2_X1 U594 ( .A(n474), .B(n485), .ZN(n475) );
  XNOR2_X1 U595 ( .A(n475), .B(n711), .ZN(n686) );
  XNOR2_X1 U596 ( .A(G902), .B(KEYINPUT15), .ZN(n674) );
  INV_X1 U597 ( .A(n674), .ZN(n476) );
  NAND2_X1 U598 ( .A1(n386), .A2(n477), .ZN(n479) );
  NAND2_X1 U599 ( .A1(n479), .A2(G214), .ZN(n622) );
  NAND2_X1 U600 ( .A1(n623), .A2(n622), .ZN(n626) );
  XOR2_X1 U601 ( .A(KEYINPUT41), .B(n480), .Z(n481) );
  XOR2_X1 U602 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n515) );
  XOR2_X1 U603 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n489) );
  NAND2_X1 U604 ( .A1(n487), .A2(G210), .ZN(n488) );
  XNOR2_X1 U605 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U606 ( .A(n491), .B(n490), .ZN(n492) );
  INV_X1 U607 ( .A(G472), .ZN(n493) );
  NAND2_X1 U608 ( .A1(n674), .A2(G234), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n494), .B(KEYINPUT20), .ZN(n506) );
  NAND2_X1 U610 ( .A1(n506), .A2(G221), .ZN(n495) );
  XNOR2_X1 U611 ( .A(KEYINPUT21), .B(n495), .ZN(n635) );
  XNOR2_X1 U612 ( .A(n354), .B(n496), .ZN(n500) );
  XNOR2_X1 U613 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U614 ( .A(n501), .B(n748), .ZN(n504) );
  AND2_X1 U615 ( .A1(n502), .A2(G221), .ZN(n503) );
  NAND2_X1 U616 ( .A1(n506), .A2(G217), .ZN(n507) );
  XNOR2_X1 U617 ( .A(n508), .B(KEYINPUT14), .ZN(n511) );
  NAND2_X1 U618 ( .A1(G952), .A2(n511), .ZN(n656) );
  NOR2_X1 U619 ( .A1(n656), .A2(G953), .ZN(n510) );
  INV_X1 U620 ( .A(KEYINPUT90), .ZN(n509) );
  XNOR2_X1 U621 ( .A(n510), .B(n509), .ZN(n571) );
  NAND2_X1 U622 ( .A1(G902), .A2(n511), .ZN(n566) );
  NOR2_X1 U623 ( .A1(G900), .A2(n566), .ZN(n512) );
  NAND2_X1 U624 ( .A1(G953), .A2(n512), .ZN(n513) );
  NAND2_X1 U625 ( .A1(n571), .A2(n513), .ZN(n529) );
  NOR2_X1 U626 ( .A1(n549), .A2(n550), .ZN(n514) );
  XOR2_X1 U627 ( .A(n515), .B(n514), .Z(n522) );
  XOR2_X1 U628 ( .A(G101), .B(G140), .Z(n517) );
  NAND2_X1 U629 ( .A1(G227), .A2(n705), .ZN(n516) );
  XNOR2_X1 U630 ( .A(n517), .B(n516), .ZN(n519) );
  XNOR2_X1 U631 ( .A(n519), .B(n518), .ZN(n520) );
  INV_X1 U632 ( .A(n554), .ZN(n526) );
  NAND2_X1 U633 ( .A1(n522), .A2(n526), .ZN(n540) );
  NOR2_X1 U634 ( .A1(n650), .A2(n540), .ZN(n524) );
  XNOR2_X1 U635 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n523) );
  XNOR2_X1 U636 ( .A(n524), .B(n523), .ZN(n758) );
  INV_X1 U637 ( .A(n536), .ZN(n543) );
  XNOR2_X1 U638 ( .A(KEYINPUT94), .B(n635), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n526), .A2(n638), .ZN(n593) );
  NAND2_X1 U640 ( .A1(n359), .A2(n622), .ZN(n527) );
  XNOR2_X1 U641 ( .A(KEYINPUT30), .B(n527), .ZN(n528) );
  XNOR2_X1 U642 ( .A(KEYINPUT70), .B(KEYINPUT84), .ZN(n532) );
  AND2_X1 U643 ( .A1(n727), .A2(n563), .ZN(n534) );
  OR2_X1 U644 ( .A1(n536), .A2(n544), .ZN(n577) );
  NOR2_X1 U645 ( .A1(n537), .A2(n577), .ZN(n538) );
  NAND2_X1 U646 ( .A1(n379), .A2(n538), .ZN(n539) );
  XNOR2_X1 U647 ( .A(n539), .B(KEYINPUT109), .ZN(n757) );
  INV_X1 U648 ( .A(n540), .ZN(n542) );
  NAND2_X1 U649 ( .A1(n542), .A2(n573), .ZN(n725) );
  NOR2_X1 U650 ( .A1(n725), .A2(n627), .ZN(n545) );
  XOR2_X1 U651 ( .A(KEYINPUT47), .B(n545), .Z(n546) );
  NOR2_X1 U652 ( .A1(n757), .A2(n546), .ZN(n556) );
  NAND2_X1 U653 ( .A1(n727), .A2(n622), .ZN(n553) );
  INV_X1 U654 ( .A(KEYINPUT104), .ZN(n547) );
  XNOR2_X1 U655 ( .A(n547), .B(KEYINPUT6), .ZN(n548) );
  XNOR2_X1 U656 ( .A(n551), .B(KEYINPUT107), .ZN(n552) );
  INV_X1 U657 ( .A(n763), .ZN(n555) );
  NAND2_X1 U658 ( .A1(n607), .A2(n559), .ZN(n560) );
  NAND2_X1 U659 ( .A1(n563), .A2(n562), .ZN(n746) );
  XOR2_X1 U660 ( .A(KEYINPUT86), .B(KEYINPUT33), .Z(n565) );
  INV_X1 U661 ( .A(n566), .ZN(n567) );
  NOR2_X1 U662 ( .A1(G898), .A2(n705), .ZN(n712) );
  NAND2_X1 U663 ( .A1(n567), .A2(n712), .ZN(n569) );
  INV_X1 U664 ( .A(KEYINPUT91), .ZN(n568) );
  XNOR2_X1 U665 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U666 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U667 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U668 ( .A(KEYINPUT34), .B(KEYINPUT74), .ZN(n575) );
  XOR2_X1 U669 ( .A(n575), .B(KEYINPUT71), .Z(n576) );
  NOR2_X1 U670 ( .A1(n625), .A2(n579), .ZN(n580) );
  XNOR2_X1 U671 ( .A(n581), .B(KEYINPUT22), .ZN(n589) );
  INV_X1 U672 ( .A(n589), .ZN(n587) );
  XNOR2_X1 U673 ( .A(n585), .B(n584), .ZN(n586) );
  AND2_X1 U674 ( .A1(n549), .A2(n435), .ZN(n590) );
  AND2_X1 U675 ( .A1(n607), .A2(n590), .ZN(n591) );
  NAND2_X1 U676 ( .A1(n587), .A2(n591), .ZN(n665) );
  XOR2_X1 U677 ( .A(KEYINPUT31), .B(n592), .Z(n729) );
  XNOR2_X1 U678 ( .A(n594), .B(KEYINPUT95), .ZN(n595) );
  NOR2_X1 U679 ( .A1(n644), .A2(n595), .ZN(n717) );
  NOR2_X1 U680 ( .A1(n729), .A2(n717), .ZN(n596) );
  XNOR2_X1 U681 ( .A(n596), .B(KEYINPUT97), .ZN(n598) );
  INV_X1 U682 ( .A(n627), .ZN(n597) );
  NAND2_X1 U683 ( .A1(n598), .A2(n597), .ZN(n599) );
  INV_X1 U684 ( .A(KEYINPUT44), .ZN(n602) );
  NOR2_X1 U685 ( .A1(n759), .A2(n602), .ZN(n600) );
  NAND2_X1 U686 ( .A1(n602), .A2(KEYINPUT66), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n587), .A2(n604), .ZN(n605) );
  XNOR2_X1 U688 ( .A(n605), .B(KEYINPUT85), .ZN(n609) );
  AND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U690 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n610) );
  XNOR2_X2 U691 ( .A(n611), .B(n610), .ZN(n675) );
  NAND2_X1 U692 ( .A1(n677), .A2(n706), .ZN(n612) );
  INV_X1 U693 ( .A(KEYINPUT2), .ZN(n671) );
  NAND2_X1 U694 ( .A1(n612), .A2(n671), .ZN(n613) );
  XNOR2_X1 U695 ( .A(n613), .B(KEYINPUT78), .ZN(n618) );
  NAND2_X1 U696 ( .A1(KEYINPUT2), .A2(n746), .ZN(n614) );
  XNOR2_X1 U697 ( .A(KEYINPUT77), .B(n614), .ZN(n615) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT83), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n682), .ZN(n620) );
  INV_X1 U700 ( .A(KEYINPUT82), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n620), .B(n619), .ZN(n661) );
  NOR2_X1 U702 ( .A1(n361), .A2(n650), .ZN(n621) );
  NOR2_X1 U703 ( .A1(G953), .A2(n621), .ZN(n659) );
  NOR2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n630) );
  NOR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U707 ( .A(n628), .B(KEYINPUT118), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U709 ( .A(KEYINPUT119), .B(n631), .Z(n632) );
  NOR2_X1 U710 ( .A1(n361), .A2(n632), .ZN(n653) );
  INV_X1 U711 ( .A(n634), .ZN(n646) );
  AND2_X1 U712 ( .A1(n635), .A2(n435), .ZN(n636) );
  XNOR2_X1 U713 ( .A(KEYINPUT49), .B(n636), .ZN(n642) );
  NOR2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n640) );
  XNOR2_X1 U715 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n640), .B(n639), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U720 ( .A(n647), .B(KEYINPUT116), .Z(n648) );
  XNOR2_X1 U721 ( .A(KEYINPUT51), .B(n648), .ZN(n649) );
  NOR2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U723 ( .A(KEYINPUT117), .B(n651), .Z(n652) );
  NOR2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U725 ( .A(KEYINPUT52), .B(n654), .ZN(n655) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U727 ( .A(KEYINPUT120), .B(n657), .Z(n658) );
  NAND2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n662), .B(KEYINPUT53), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n665), .B(G110), .ZN(G12) );
  XOR2_X1 U732 ( .A(G119), .B(KEYINPUT126), .Z(n667) );
  XOR2_X1 U733 ( .A(n667), .B(n666), .Z(G21) );
  XNOR2_X1 U734 ( .A(n668), .B(G101), .ZN(G3) );
  NOR2_X1 U735 ( .A1(n674), .A2(KEYINPUT81), .ZN(n670) );
  AND2_X2 U736 ( .A1(n675), .A2(n670), .ZN(n669) );
  INV_X1 U737 ( .A(n670), .ZN(n672) );
  OR2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U739 ( .A1(n674), .A2(KEYINPUT2), .ZN(n676) );
  AND2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n678) );
  NAND2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U742 ( .A1(n679), .A2(KEYINPUT81), .ZN(n680) );
  NAND2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U744 ( .A1(n732), .A2(G210), .ZN(n688) );
  XNOR2_X1 U745 ( .A(KEYINPUT79), .B(KEYINPUT54), .ZN(n684) );
  XNOR2_X1 U746 ( .A(n684), .B(KEYINPUT55), .ZN(n685) );
  XNOR2_X1 U747 ( .A(n688), .B(n687), .ZN(n690) );
  INV_X1 U748 ( .A(G952), .ZN(n689) );
  NOR2_X2 U749 ( .A1(n690), .A2(n745), .ZN(n692) );
  XNOR2_X1 U750 ( .A(KEYINPUT122), .B(KEYINPUT56), .ZN(n691) );
  XNOR2_X1 U751 ( .A(n692), .B(n691), .ZN(G51) );
  NAND2_X1 U752 ( .A1(n732), .A2(G475), .ZN(n696) );
  XNOR2_X1 U753 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n693) );
  XNOR2_X1 U754 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X2 U755 ( .A1(n697), .A2(n745), .ZN(n698) );
  XNOR2_X1 U756 ( .A(n698), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U757 ( .A1(n732), .A2(G472), .ZN(n701) );
  XNOR2_X1 U758 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X2 U759 ( .A1(n702), .A2(n745), .ZN(n704) );
  XOR2_X1 U760 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n703) );
  XNOR2_X1 U761 ( .A(n704), .B(n703), .ZN(G57) );
  NAND2_X1 U762 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n707) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n707), .ZN(n708) );
  NAND2_X1 U765 ( .A1(n708), .A2(G898), .ZN(n709) );
  NAND2_X1 U766 ( .A1(n710), .A2(n709), .ZN(n715) );
  INV_X1 U767 ( .A(n711), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U769 ( .A(n715), .B(n714), .ZN(G69) );
  NAND2_X1 U770 ( .A1(n717), .A2(n727), .ZN(n716) );
  XNOR2_X1 U771 ( .A(n716), .B(G104), .ZN(G6) );
  XOR2_X1 U772 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n719) );
  NAND2_X1 U773 ( .A1(n717), .A2(n730), .ZN(n718) );
  XNOR2_X1 U774 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U775 ( .A(G107), .B(n720), .ZN(G9) );
  NOR2_X1 U776 ( .A1(n725), .A2(n721), .ZN(n723) );
  XNOR2_X1 U777 ( .A(G128), .B(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n723), .B(n722), .ZN(G30) );
  INV_X1 U779 ( .A(n727), .ZN(n724) );
  NOR2_X1 U780 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U781 ( .A(G146), .B(n726), .Z(G48) );
  NAND2_X1 U782 ( .A1(n729), .A2(n727), .ZN(n728) );
  XNOR2_X1 U783 ( .A(n728), .B(G113), .ZN(G15) );
  NAND2_X1 U784 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U785 ( .A(n731), .B(G116), .ZN(G18) );
  XNOR2_X1 U786 ( .A(G134), .B(n746), .ZN(G36) );
  NAND2_X1 U787 ( .A1(n741), .A2(G469), .ZN(n735) );
  XOR2_X1 U788 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n733) );
  NOR2_X1 U789 ( .A1(n745), .A2(n736), .ZN(G54) );
  NAND2_X1 U790 ( .A1(n741), .A2(G478), .ZN(n739) );
  NOR2_X1 U791 ( .A1(n745), .A2(n740), .ZN(G63) );
  NAND2_X1 U792 ( .A1(n741), .A2(G217), .ZN(n743) );
  XNOR2_X1 U793 ( .A(n743), .B(n742), .ZN(n744) );
  NOR2_X1 U794 ( .A1(n745), .A2(n744), .ZN(G66) );
  XOR2_X1 U795 ( .A(n747), .B(n748), .Z(n752) );
  INV_X1 U796 ( .A(n752), .ZN(n749) );
  NOR2_X1 U797 ( .A1(G953), .A2(n750), .ZN(n751) );
  XNOR2_X1 U798 ( .A(KEYINPUT125), .B(n751), .ZN(n756) );
  XOR2_X1 U799 ( .A(G227), .B(n752), .Z(n753) );
  NAND2_X1 U800 ( .A1(n753), .A2(G900), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n754), .A2(G953), .ZN(n755) );
  NAND2_X1 U802 ( .A1(n756), .A2(n755), .ZN(G72) );
  XOR2_X1 U803 ( .A(G143), .B(n757), .Z(G45) );
  XOR2_X1 U804 ( .A(G137), .B(n758), .Z(G39) );
  XOR2_X1 U805 ( .A(n360), .B(G122), .Z(G24) );
  XNOR2_X1 U806 ( .A(G131), .B(KEYINPUT127), .ZN(n761) );
  XNOR2_X1 U807 ( .A(n761), .B(n760), .ZN(G33) );
  XOR2_X1 U808 ( .A(G140), .B(n762), .Z(G42) );
  XNOR2_X1 U809 ( .A(n763), .B(KEYINPUT114), .ZN(n764) );
  XNOR2_X1 U810 ( .A(n764), .B(KEYINPUT37), .ZN(n765) );
  XNOR2_X1 U811 ( .A(G125), .B(n765), .ZN(G27) );
endmodule

