//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G128), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT24), .B(G110), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT74), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT74), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n196), .B2(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n204));
  INV_X1    g018(.A(new_n195), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n204), .B(new_n193), .C1(new_n205), .C2(KEYINPUT23), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G110), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT75), .A3(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(G125), .ZN(new_n212));
  INV_X1    g026(.A(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(KEYINPUT16), .B(new_n211), .C1(new_n215), .C2(KEYINPUT75), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n209), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n209), .A3(new_n218), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(KEYINPUT76), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT76), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n216), .A2(new_n222), .A3(new_n209), .A4(new_n218), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n208), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n216), .A2(new_n218), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n212), .A2(new_n214), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n209), .ZN(new_n228));
  OAI22_X1  g042(.A1(new_n206), .A2(G110), .B1(new_n197), .B2(new_n199), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n191), .B1(new_n224), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n220), .A2(KEYINPUT76), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n223), .A3(new_n226), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n207), .A3(new_n203), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n230), .A3(new_n190), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n232), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT77), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT77), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n232), .A2(new_n236), .A3(new_n241), .A4(new_n237), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n232), .A2(new_n236), .A3(KEYINPUT25), .A4(new_n237), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT78), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n239), .A2(KEYINPUT78), .A3(new_n240), .A4(new_n242), .ZN(new_n249));
  INV_X1    g063(.A(G217), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G234), .B2(new_n237), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(G902), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n232), .A2(new_n236), .A3(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G110), .B(G122), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT2), .B(G113), .Z(new_n258));
  XNOR2_X1  g072(.A(G116), .B(G119), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT2), .B(G113), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G119), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n192), .A2(G116), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n260), .A2(new_n265), .A3(KEYINPUT65), .ZN(new_n266));
  OR3_X1    g080(.A1(new_n258), .A2(KEYINPUT65), .A3(new_n259), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT79), .ZN(new_n269));
  INV_X1    g083(.A(G107), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(G104), .ZN(new_n271));
  INV_X1    g085(.A(G104), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT79), .A3(G107), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n272), .B2(G107), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n270), .A2(KEYINPUT3), .A3(G104), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G101), .ZN(new_n280));
  INV_X1    g094(.A(G101), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n278), .A2(new_n281), .A3(new_n271), .A4(new_n273), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(KEYINPUT4), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n284), .A3(G101), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n268), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n287));
  INV_X1    g101(.A(G113), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n263), .B2(new_n289), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n287), .A2(new_n290), .B1(new_n258), .B2(new_n259), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n272), .A2(G107), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n270), .A2(G104), .ZN(new_n293));
  OAI21_X1  g107(.A(G101), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n282), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT82), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n282), .A2(new_n294), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT82), .A3(new_n291), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n257), .B1(new_n286), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n268), .A2(new_n283), .A3(new_n285), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n302), .A2(new_n256), .A3(new_n297), .A4(new_n299), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(KEYINPUT6), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G143), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(G146), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n209), .A2(G143), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n194), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n305), .A2(KEYINPUT1), .A3(G146), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n209), .A2(G143), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(G146), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(G128), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n308), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n213), .ZN(new_n316));
  AOI211_X1 g130(.A(KEYINPUT0), .B(new_n194), .C1(new_n311), .C2(new_n312), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n311), .A2(new_n312), .A3(G128), .ZN(new_n318));
  XNOR2_X1  g132(.A(G143), .B(G146), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT0), .A2(G128), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n317), .B1(new_n322), .B2(KEYINPUT0), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n316), .B1(new_n213), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G224), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(G953), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT83), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n324), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT6), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n329), .B(new_n257), .C1(new_n286), .C2(new_n300), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n304), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n256), .B(KEYINPUT8), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n298), .A2(new_n291), .ZN(new_n333));
  INV_X1    g147(.A(new_n295), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT7), .B1(new_n325), .B2(G953), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n324), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n324), .A2(new_n336), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(G902), .B1(new_n340), .B2(new_n303), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n331), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(G210), .B1(G237), .B2(G902), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n331), .A2(new_n341), .A3(new_n343), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G214), .B1(G237), .B2(G902), .ZN(new_n348));
  NAND2_X1  g162(.A1(G234), .A2(G237), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(G952), .A3(new_n188), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT21), .B(G898), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(G902), .A3(G953), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n347), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT13), .B1(new_n194), .B2(G143), .ZN(new_n356));
  INV_X1    g170(.A(G134), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G128), .B(G143), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT87), .B(G122), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(new_n262), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n262), .A2(G122), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n362), .A2(new_n270), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n270), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n363), .B(KEYINPUT14), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n361), .A2(new_n262), .ZN(new_n368));
  OAI21_X1  g182(.A(G107), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n362), .A2(new_n270), .A3(new_n363), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n359), .B(new_n357), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n374), .A2(new_n250), .A3(G953), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n366), .A2(new_n372), .A3(new_n375), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n237), .ZN(new_n380));
  INV_X1    g194(.A(G478), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT88), .A2(KEYINPUT15), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(KEYINPUT88), .A2(KEYINPUT15), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n377), .B2(new_n378), .ZN(new_n387));
  INV_X1    g201(.A(new_n385), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n391));
  INV_X1    g205(.A(G237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n188), .A3(G214), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n305), .ZN(new_n394));
  NOR2_X1   g208(.A1(G237), .A2(G953), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(G143), .A3(G214), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT18), .A2(G131), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n394), .B2(new_n396), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(G146), .B(new_n211), .C1(new_n215), .C2(KEYINPUT75), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n401), .A2(KEYINPUT84), .A3(new_n228), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT84), .B1(new_n401), .B2(new_n228), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n391), .B(new_n400), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT85), .ZN(new_n406));
  INV_X1    g220(.A(new_n234), .ZN(new_n407));
  INV_X1    g221(.A(new_n396), .ZN(new_n408));
  AOI21_X1  g222(.A(G143), .B1(new_n395), .B2(G214), .ZN(new_n409));
  OAI21_X1  g223(.A(G131), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  INV_X1    g225(.A(G131), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n394), .A2(new_n412), .A3(new_n396), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT17), .B(G131), .C1(new_n408), .C2(new_n409), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n404), .A2(new_n406), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n272), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n406), .A2(new_n404), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT86), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n221), .A2(new_n416), .A3(new_n223), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n419), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n401), .A2(new_n228), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n401), .A2(KEYINPUT84), .A3(new_n228), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n391), .B1(new_n429), .B2(new_n400), .ZN(new_n430));
  INV_X1    g244(.A(new_n404), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n419), .B(new_n423), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT86), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n420), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G475), .B1(new_n434), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n219), .B1(new_n410), .B2(new_n413), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n227), .A2(KEYINPUT19), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n211), .B1(new_n215), .B2(KEYINPUT75), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n439), .B2(KEYINPUT19), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n437), .B1(G146), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n419), .B1(new_n421), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n422), .B1(new_n417), .B2(new_n419), .ZN(new_n444));
  INV_X1    g258(.A(new_n424), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(G475), .A2(G902), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n436), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n442), .B1(new_n433), .B2(new_n424), .ZN(new_n449));
  INV_X1    g263(.A(new_n447), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n449), .A2(KEYINPUT20), .A3(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n390), .B(new_n435), .C1(new_n448), .C2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT11), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n357), .B2(G137), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n357), .A2(G137), .ZN(new_n455));
  INV_X1    g269(.A(G137), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(KEYINPUT11), .A3(G134), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G131), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n454), .A2(new_n457), .A3(new_n412), .A4(new_n455), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n308), .A2(new_n310), .A3(new_n314), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n282), .B2(new_n294), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n314), .A2(KEYINPUT80), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n311), .A2(new_n312), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n309), .B1(new_n465), .B2(new_n194), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT80), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n319), .A2(new_n467), .A3(new_n313), .A4(G128), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n282), .A2(new_n294), .ZN(new_n470));
  OAI22_X1  g284(.A1(new_n463), .A2(KEYINPUT81), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n315), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT81), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n461), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT12), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT0), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n320), .B1(new_n306), .B2(new_n307), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(new_n318), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n479), .A2(KEYINPUT66), .A3(new_n317), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT66), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n311), .A2(new_n312), .A3(G128), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n311), .A2(new_n312), .B1(KEYINPUT0), .B2(G128), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT0), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n317), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n285), .B(new_n283), .C1(new_n480), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n282), .A3(new_n294), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT10), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n466), .B2(new_n314), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n489), .A2(new_n490), .B1(new_n298), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n459), .A2(new_n460), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n487), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G110), .B(G140), .ZN(new_n495));
  INV_X1    g309(.A(G227), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G953), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n495), .B(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT12), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n500), .B(new_n461), .C1(new_n471), .C2(new_n474), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n476), .A2(new_n494), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n487), .A2(new_n492), .A3(new_n493), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n493), .B1(new_n487), .B2(new_n492), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(G902), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G469), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n237), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n472), .A2(new_n473), .B1(new_n298), .B2(new_n488), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n463), .A2(KEYINPUT81), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n493), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n494), .B1(new_n513), .B2(new_n500), .ZN(new_n514));
  INV_X1    g328(.A(new_n501), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n498), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR3_X1    g330(.A1(new_n503), .A2(new_n504), .A3(new_n498), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(G469), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n508), .A2(new_n510), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G221), .B1(new_n374), .B2(G902), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n355), .A2(new_n452), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G472), .A2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n456), .A2(G134), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n357), .A2(G137), .ZN(new_n526));
  OAI21_X1  g340(.A(G131), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n460), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n323), .A2(new_n461), .B1(new_n528), .B2(new_n462), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT64), .B1(new_n529), .B2(KEYINPUT30), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n462), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n484), .A2(new_n485), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(new_n493), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT64), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n461), .B1(new_n480), .B2(new_n486), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n460), .A2(new_n527), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT67), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n460), .A2(new_n527), .A3(KEYINPUT67), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n462), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT68), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n539), .A2(new_n540), .B1(new_n466), .B2(new_n314), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT68), .A3(new_n542), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n538), .A2(KEYINPUT30), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n537), .A2(new_n268), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT31), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT26), .B(G101), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n395), .A2(G210), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT70), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n553), .B(new_n555), .ZN(new_n556));
  AND4_X1   g370(.A1(KEYINPUT68), .A2(new_n541), .A3(new_n542), .A4(new_n462), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT68), .B1(new_n546), .B2(new_n542), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT66), .B1(new_n479), .B2(new_n317), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n484), .A2(new_n485), .A3(new_n481), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n268), .B1(new_n562), .B2(new_n461), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n556), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n549), .A2(new_n550), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT71), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT71), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n549), .A2(new_n567), .A3(new_n550), .A4(new_n564), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT72), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n493), .B1(new_n560), .B2(new_n561), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n541), .A2(new_n542), .A3(new_n462), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n571), .A2(new_n268), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n570), .B1(new_n573), .B2(KEYINPUT28), .ZN(new_n574));
  INV_X1    g388(.A(new_n268), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n538), .A2(new_n575), .A3(new_n543), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT28), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(KEYINPUT72), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n559), .A2(new_n563), .B1(new_n268), .B2(new_n533), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n574), .B(new_n578), .C1(new_n577), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n549), .A2(new_n564), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n580), .A2(new_n556), .B1(new_n581), .B2(KEYINPUT31), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n524), .B1(new_n569), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT73), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI211_X1 g399(.A(KEYINPUT73), .B(new_n524), .C1(new_n569), .C2(new_n582), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT32), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n559), .A2(new_n563), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n549), .A2(new_n556), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n538), .A2(new_n545), .A3(new_n547), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n592), .A2(new_n268), .B1(new_n559), .B2(new_n563), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n574), .B(new_n578), .C1(new_n593), .C2(new_n577), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n594), .A2(KEYINPUT29), .ZN(new_n595));
  INV_X1    g409(.A(new_n556), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n580), .B2(KEYINPUT29), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n591), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g412(.A1(KEYINPUT32), .A2(new_n583), .B1(new_n598), .B2(G472), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n255), .B(new_n522), .C1(new_n587), .C2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  NAND2_X1  g416(.A1(new_n569), .A2(new_n582), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n237), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(KEYINPUT89), .A3(G472), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT89), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n569), .B2(new_n582), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n585), .A2(new_n586), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n252), .A2(new_n254), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n612), .A2(new_n613), .A3(new_n521), .ZN(new_n614));
  INV_X1    g428(.A(new_n348), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n343), .B1(new_n331), .B2(new_n341), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT90), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n347), .B2(new_n617), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n354), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n435), .B1(new_n448), .B2(new_n451), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n379), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT91), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n377), .B(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT92), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n623), .B1(new_n378), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n627), .B2(new_n378), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n624), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n381), .A2(G902), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI22_X1  g446(.A1(new_n630), .A2(new_n632), .B1(G478), .B2(new_n387), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n622), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n621), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n614), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  NAND3_X1  g452(.A1(new_n446), .A2(new_n436), .A3(new_n447), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT20), .B1(new_n449), .B2(new_n450), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n444), .A2(new_n445), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n237), .B1(new_n641), .B2(new_n420), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n639), .A2(new_n640), .B1(new_n642), .B2(G475), .ZN(new_n643));
  INV_X1    g457(.A(new_n390), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n621), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n614), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  OAI22_X1  g463(.A1(new_n224), .A2(new_n231), .B1(KEYINPUT36), .B2(new_n191), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n235), .A2(new_n230), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n653), .A2(KEYINPUT93), .A3(new_n253), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT93), .B1(new_n653), .B2(new_n253), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n249), .A2(new_n251), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT25), .B1(new_n238), .B2(KEYINPUT77), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n246), .B1(new_n658), .B2(new_n242), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n656), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT94), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n252), .A2(KEYINPUT94), .A3(new_n656), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n664), .A2(new_n611), .A3(new_n522), .A4(new_n610), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT95), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT37), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  NAND2_X1  g482(.A1(new_n662), .A2(new_n663), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n603), .A2(new_n523), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT73), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT32), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n583), .A2(new_n584), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n669), .B1(new_n674), .B2(new_n599), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n350), .B1(new_n353), .B2(G900), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT96), .Z(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n643), .A2(new_n644), .A3(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n679), .A2(new_n521), .A3(new_n619), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  XNOR2_X1  g496(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n347), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n622), .A2(new_n644), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n684), .A2(new_n615), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n593), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n237), .B1(new_n687), .B2(new_n596), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n556), .B1(new_n549), .B2(new_n588), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n583), .A2(KEYINPUT32), .B1(G472), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n674), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n660), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n677), .B(KEYINPUT39), .Z(new_n694));
  NAND3_X1  g508(.A1(new_n519), .A2(new_n520), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT40), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n686), .A2(new_n692), .A3(new_n693), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NAND3_X1  g513(.A1(new_n622), .A2(new_n633), .A3(new_n678), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n700), .A2(new_n521), .A3(new_n619), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n675), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  AOI21_X1  g517(.A(new_n613), .B1(new_n674), .B2(new_n599), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n502), .A2(new_n505), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n237), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT98), .B1(new_n506), .B2(new_n507), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n706), .A2(KEYINPUT98), .A3(G469), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT99), .B1(new_n711), .B2(new_n520), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT99), .ZN(new_n713));
  INV_X1    g527(.A(new_n520), .ZN(new_n714));
  AOI211_X1 g528(.A(new_n713), .B(new_n714), .C1(new_n709), .C2(new_n710), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n704), .A2(new_n635), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND3_X1  g533(.A1(new_n704), .A2(new_n646), .A3(new_n716), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  INV_X1    g535(.A(new_n621), .ZN(new_n722));
  INV_X1    g536(.A(new_n452), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n675), .A2(new_n722), .A3(new_n723), .A4(new_n716), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  INV_X1    g539(.A(KEYINPUT100), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n550), .B1(new_n549), .B2(new_n564), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n594), .B2(new_n556), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n524), .B1(new_n569), .B2(new_n728), .ZN(new_n729));
  OAI22_X1  g543(.A1(new_n726), .A2(new_n729), .B1(new_n607), .B2(new_n608), .ZN(new_n730));
  AOI211_X1 g544(.A(KEYINPUT100), .B(new_n524), .C1(new_n569), .C2(new_n728), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n730), .A2(new_n685), .A3(new_n613), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n722), .A3(new_n716), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT101), .B(G122), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G24));
  NOR3_X1   g549(.A1(new_n730), .A2(new_n693), .A3(new_n731), .ZN(new_n736));
  INV_X1    g550(.A(new_n700), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n716), .A2(new_n620), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NAND3_X1  g553(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n520), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n476), .A2(new_n494), .A3(new_n501), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n743), .A2(KEYINPUT102), .A3(new_n498), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT102), .B1(new_n743), .B2(new_n498), .ZN(new_n745));
  OAI211_X1 g559(.A(G469), .B(new_n517), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT103), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n509), .B1(new_n506), .B2(new_n507), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT102), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n516), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n743), .A2(KEYINPUT102), .A3(new_n498), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT103), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n753), .A3(G469), .A4(new_n517), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n747), .A2(new_n748), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT104), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n747), .A2(new_n754), .A3(new_n757), .A4(new_n748), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n742), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n670), .A2(new_n672), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n613), .B1(new_n599), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n759), .A2(KEYINPUT42), .A3(new_n737), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n704), .A2(new_n759), .A3(new_n737), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n763), .A2(KEYINPUT105), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT105), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  INV_X1    g582(.A(new_n679), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n704), .A2(new_n759), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n643), .B2(new_n633), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n633), .B(new_n435), .C1(new_n448), .C2(new_n451), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(KEYINPUT43), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT107), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n643), .A2(new_n772), .A3(new_n633), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT107), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n774), .A2(KEYINPUT43), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n776), .A2(new_n612), .A3(new_n660), .A4(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n740), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(KEYINPUT45), .B(new_n517), .C1(new_n744), .C2(new_n745), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n516), .A2(new_n517), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n507), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n510), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n509), .B1(new_n784), .B2(new_n787), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT46), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n508), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(KEYINPUT106), .A3(new_n520), .A4(new_n694), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n508), .B1(new_n792), .B2(KEYINPUT46), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n790), .B(new_n509), .C1(new_n784), .C2(new_n787), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n520), .B(new_n694), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT106), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n693), .B1(new_n610), .B2(new_n611), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(KEYINPUT44), .A3(new_n780), .A4(new_n776), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n783), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  NOR2_X1   g619(.A1(new_n255), .A2(new_n740), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n737), .A3(new_n674), .A4(new_n599), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n520), .B1(new_n796), .B2(new_n797), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(KEYINPUT47), .B(new_n520), .C1(new_n796), .C2(new_n797), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n210), .ZN(G42));
  NOR3_X1   g627(.A1(new_n692), .A2(new_n613), .A3(new_n350), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n716), .A3(new_n741), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n815), .A2(new_n622), .A3(new_n633), .ZN(new_n816));
  INV_X1    g630(.A(new_n350), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n777), .A2(new_n817), .A3(new_n779), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n818), .A2(new_n613), .A3(new_n731), .A4(new_n730), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n615), .A3(new_n684), .A4(new_n716), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT50), .ZN(new_n821));
  INV_X1    g635(.A(new_n716), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n740), .A3(new_n818), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n816), .B(new_n821), .C1(new_n736), .C2(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n819), .A2(new_n741), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n711), .A2(new_n714), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n810), .A2(new_n811), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(KEYINPUT51), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n188), .A2(G952), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n822), .A2(new_n619), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(new_n819), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n634), .B2(new_n815), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n823), .A2(new_n761), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(KEYINPUT114), .A3(KEYINPUT48), .ZN(new_n835));
  XOR2_X1   g649(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n836));
  AOI211_X1 g650(.A(new_n833), .B(new_n835), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n674), .A2(new_n599), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n839), .B(new_n664), .C1(new_n680), .C2(new_n701), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n678), .A2(new_n520), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n685), .A2(new_n619), .A3(new_n660), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n756), .A2(new_n758), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n692), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n738), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n840), .A2(new_n738), .A3(KEYINPUT52), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n724), .A2(new_n717), .A3(new_n720), .A4(new_n733), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n759), .A2(new_n737), .A3(new_n736), .ZN(new_n852));
  INV_X1    g666(.A(new_n521), .ZN(new_n853));
  OR3_X1    g667(.A1(new_n386), .A2(KEYINPUT108), .A3(new_n389), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT108), .B1(new_n386), .B2(new_n389), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n622), .A2(new_n740), .A3(new_n856), .A4(new_n677), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n839), .A2(new_n853), .A3(new_n664), .A4(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n770), .A2(new_n852), .A3(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n856), .B(new_n435), .C1(new_n448), .C2(new_n451), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n355), .B1(new_n860), .B2(new_n634), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n613), .A2(new_n521), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n611), .A3(new_n610), .A4(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n665), .A2(new_n601), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n767), .A2(new_n849), .A3(new_n851), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT53), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n847), .A2(KEYINPUT109), .A3(new_n848), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT109), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n845), .A2(new_n869), .A3(new_n846), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n767), .A2(new_n872), .A3(new_n851), .A4(new_n865), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n867), .B(KEYINPUT54), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT110), .B1(new_n859), .B2(new_n864), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n665), .A2(new_n601), .A3(new_n863), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n857), .A2(new_n853), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n730), .A2(new_n700), .A3(new_n693), .A4(new_n731), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n675), .A2(new_n877), .B1(new_n878), .B2(new_n759), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT110), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n876), .A2(new_n879), .A3(new_n880), .A4(new_n770), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n875), .A2(new_n881), .A3(KEYINPUT53), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n763), .A2(new_n764), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT105), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n763), .A2(KEYINPUT105), .A3(new_n764), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n850), .B1(new_n887), .B2(new_n762), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n882), .A2(new_n888), .A3(new_n870), .A4(new_n868), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n866), .A2(new_n872), .ZN(new_n890));
  XOR2_X1   g704(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n874), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n810), .A2(new_n811), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT112), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n826), .B(KEYINPUT113), .Z(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n894), .A2(KEYINPUT112), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n825), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT51), .B1(new_n824), .B2(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n838), .A2(new_n893), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n684), .A2(new_n348), .A3(new_n520), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n774), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n711), .B(KEYINPUT49), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n255), .A3(new_n905), .ZN(new_n906));
  OAI22_X1  g720(.A1(new_n901), .A2(new_n902), .B1(new_n692), .B2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n188), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(G210), .A2(G902), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n889), .B2(new_n890), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n304), .A2(new_n330), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n328), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT55), .Z(new_n914));
  OR2_X1    g728(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n909), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n911), .B2(KEYINPUT115), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT115), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n919), .B(new_n910), .C1(new_n889), .C2(new_n890), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n914), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT116), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT116), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n923), .B(new_n914), .C1(new_n918), .C2(new_n920), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n916), .B1(new_n922), .B2(new_n924), .ZN(G51));
  AND3_X1   g739(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n891), .B1(new_n889), .B2(new_n890), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n509), .B(KEYINPUT57), .Z(new_n929));
  OAI21_X1  g743(.A(new_n705), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n889), .A2(new_n890), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n931), .A2(G902), .A3(new_n784), .A4(new_n787), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n908), .B1(new_n930), .B2(new_n932), .ZN(G54));
  NAND4_X1  g747(.A1(new_n931), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n934), .A2(new_n449), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n449), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n935), .A2(new_n936), .A3(new_n908), .ZN(G60));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT59), .Z(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n893), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n630), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT117), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n630), .A2(new_n939), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n926), .B2(new_n927), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n942), .A2(new_n943), .A3(new_n909), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n909), .ZN(new_n947));
  INV_X1    g761(.A(new_n630), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n893), .B2(new_n940), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT117), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(G63));
  XNOR2_X1  g765(.A(KEYINPUT118), .B(KEYINPUT61), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n232), .A2(new_n236), .ZN(new_n954));
  INV_X1    g768(.A(new_n931), .ZN(new_n955));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n954), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n909), .ZN(new_n959));
  INV_X1    g773(.A(new_n653), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n955), .A2(new_n960), .A3(new_n957), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n953), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n961), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n963), .A2(new_n909), .A3(new_n958), .A4(new_n952), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(G66));
  NAND2_X1  g779(.A1(new_n851), .A2(new_n876), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n188), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n351), .B2(new_n325), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT119), .Z(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT120), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n912), .B1(G898), .B2(new_n188), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G69));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n537), .A2(new_n548), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(new_n440), .Z(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n840), .A2(new_n698), .A3(new_n738), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n840), .A2(new_n698), .A3(new_n738), .A4(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n860), .A2(new_n634), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n695), .A2(new_n740), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n839), .A2(new_n255), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT121), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n704), .A2(KEYINPUT121), .A3(new_n983), .A4(new_n984), .ZN(new_n988));
  INV_X1    g802(.A(new_n807), .ZN(new_n989));
  AOI22_X1  g803(.A1(new_n987), .A2(new_n988), .B1(new_n894), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n982), .A2(new_n804), .A3(new_n990), .ZN(new_n991));
  AOI211_X1 g805(.A(KEYINPUT122), .B(new_n977), .C1(new_n991), .C2(new_n188), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT122), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n980), .A2(new_n981), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n804), .A2(new_n990), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n188), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n993), .B1(new_n996), .B2(new_n976), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(G900), .ZN(new_n999));
  OAI21_X1  g813(.A(G953), .B1(new_n496), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(G953), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT123), .Z(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n685), .A2(new_n619), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n761), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n800), .A2(new_n795), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT124), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n800), .A2(new_n795), .A3(new_n1005), .A4(KEYINPUT124), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n840), .A2(new_n738), .ZN(new_n1011));
  INV_X1    g825(.A(new_n770), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1011), .A2(new_n812), .A3(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n767), .A2(new_n1010), .A3(new_n804), .A4(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1003), .B1(new_n1014), .B2(new_n188), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1000), .B1(new_n1015), .B2(new_n976), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n974), .B1(new_n998), .B2(new_n1016), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n804), .A2(new_n990), .ZN(new_n1018));
  AOI21_X1  g832(.A(G953), .B1(new_n1018), .B2(new_n982), .ZN(new_n1019));
  OAI21_X1  g833(.A(KEYINPUT122), .B1(new_n1019), .B2(new_n977), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n977), .B1(new_n991), .B2(new_n188), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n993), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1014), .A2(new_n188), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n1002), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n977), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1023), .A2(KEYINPUT125), .A3(new_n1000), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n976), .B1(new_n1024), .B2(new_n1002), .ZN(new_n1028));
  OAI221_X1 g842(.A(G953), .B1(new_n496), .B2(new_n999), .C1(new_n1028), .C2(new_n1021), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1017), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT126), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1017), .A2(new_n1027), .A3(new_n1029), .A4(KEYINPUT126), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(G72));
  NAND2_X1  g848(.A1(G472), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT63), .Z(new_n1036));
  OAI21_X1  g850(.A(new_n1036), .B1(new_n1014), .B2(new_n966), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(new_n589), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1036), .B1(new_n991), .B2(new_n966), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(new_n689), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1038), .A2(new_n1040), .A3(new_n909), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n867), .B1(new_n871), .B2(new_n873), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1036), .ZN(new_n1043));
  NOR4_X1   g857(.A1(new_n1042), .A2(new_n589), .A3(new_n689), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT127), .ZN(new_n1045));
  OR2_X1    g859(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1041), .B1(new_n1046), .B2(new_n1047), .ZN(G57));
endmodule


