

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  NOR2_X1 U324 ( .A1(n589), .A2(n483), .ZN(n484) );
  XNOR2_X1 U325 ( .A(n413), .B(n339), .ZN(n340) );
  XNOR2_X1 U326 ( .A(n379), .B(n382), .ZN(n383) );
  XNOR2_X1 U327 ( .A(n468), .B(n292), .ZN(n576) );
  NAND2_X1 U328 ( .A1(n545), .A2(n475), .ZN(n468) );
  XNOR2_X1 U329 ( .A(KEYINPUT38), .B(n488), .ZN(n514) );
  XNOR2_X1 U330 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n292) );
  XOR2_X1 U331 ( .A(n348), .B(n347), .Z(n293) );
  XNOR2_X1 U332 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n351) );
  XNOR2_X1 U333 ( .A(n352), .B(n351), .ZN(n374) );
  XNOR2_X1 U334 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n400) );
  INV_X1 U335 ( .A(KEYINPUT20), .ZN(n300) );
  XNOR2_X1 U336 ( .A(n401), .B(n400), .ZN(n539) );
  XNOR2_X1 U337 ( .A(n301), .B(n300), .ZN(n302) );
  INV_X1 U338 ( .A(G134GAT), .ZN(n380) );
  INV_X1 U339 ( .A(n539), .ZN(n540) );
  XNOR2_X1 U340 ( .A(n427), .B(n302), .ZN(n303) );
  XNOR2_X1 U341 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U342 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U343 ( .A(n388), .B(n293), .ZN(n349) );
  XOR2_X1 U344 ( .A(KEYINPUT36), .B(n553), .Z(n589) );
  XNOR2_X1 U345 ( .A(n350), .B(n349), .ZN(n517) );
  NOR2_X1 U346 ( .A1(n545), .A2(n460), .ZN(n574) );
  INV_X1 U347 ( .A(G43GAT), .ZN(n489) );
  XNOR2_X1 U348 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n492) );
  XNOR2_X1 U349 ( .A(n489), .B(KEYINPUT40), .ZN(n490) );
  XNOR2_X1 U350 ( .A(n493), .B(n492), .ZN(G1351GAT) );
  XNOR2_X1 U351 ( .A(n491), .B(n490), .ZN(G1330GAT) );
  XOR2_X1 U352 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n295) );
  XNOR2_X1 U353 ( .A(G176GAT), .B(KEYINPUT84), .ZN(n294) );
  XNOR2_X1 U354 ( .A(n295), .B(n294), .ZN(n307) );
  XOR2_X1 U355 ( .A(G15GAT), .B(G127GAT), .Z(n356) );
  XOR2_X1 U356 ( .A(G99GAT), .B(n356), .Z(n297) );
  XOR2_X1 U357 ( .A(G120GAT), .B(G71GAT), .Z(n330) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(n330), .ZN(n296) );
  XNOR2_X1 U359 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U360 ( .A(n298), .B(G190GAT), .Z(n305) );
  XNOR2_X1 U361 ( .A(G113GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U362 ( .A(n299), .B(KEYINPUT0), .ZN(n427) );
  NAND2_X1 U363 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(n303), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U366 ( .A(n307), .B(n306), .ZN(n312) );
  XOR2_X1 U367 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n309) );
  XNOR2_X1 U368 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n309), .B(n308), .ZN(n311) );
  XOR2_X1 U370 ( .A(G183GAT), .B(KEYINPUT86), .Z(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n412) );
  XNOR2_X2 U372 ( .A(n312), .B(n412), .ZN(n545) );
  INV_X1 U373 ( .A(KEYINPUT41), .ZN(n332) );
  INV_X1 U374 ( .A(G106GAT), .ZN(n313) );
  NAND2_X1 U375 ( .A1(n313), .A2(G92GAT), .ZN(n316) );
  INV_X1 U376 ( .A(G92GAT), .ZN(n314) );
  NAND2_X1 U377 ( .A1(n314), .A2(G106GAT), .ZN(n315) );
  NAND2_X1 U378 ( .A1(n316), .A2(n315), .ZN(n318) );
  XNOR2_X1 U379 ( .A(G99GAT), .B(G85GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n379) );
  XNOR2_X1 U381 ( .A(G148GAT), .B(G78GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n319), .B(G204GAT), .ZN(n451) );
  XNOR2_X1 U383 ( .A(n379), .B(n451), .ZN(n325) );
  XNOR2_X1 U384 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n321) );
  AND2_X1 U385 ( .A1(G230GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U386 ( .A(n321), .B(n320), .ZN(n323) );
  INV_X1 U387 ( .A(KEYINPUT32), .ZN(n322) );
  XNOR2_X1 U388 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U390 ( .A(G57GAT), .B(KEYINPUT13), .Z(n359) );
  XNOR2_X1 U391 ( .A(n326), .B(n359), .ZN(n328) );
  XOR2_X1 U392 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n327) );
  XNOR2_X1 U393 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U395 ( .A(G176GAT), .B(G64GAT), .Z(n410) );
  XNOR2_X1 U396 ( .A(n331), .B(n410), .ZN(n395) );
  XNOR2_X1 U397 ( .A(n332), .B(n395), .ZN(n461) );
  XOR2_X1 U398 ( .A(G141GAT), .B(G113GAT), .Z(n334) );
  XNOR2_X1 U399 ( .A(G50GAT), .B(G36GAT), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U401 ( .A(G197GAT), .B(KEYINPUT70), .Z(n336) );
  XNOR2_X1 U402 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U404 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U405 ( .A(G1GAT), .B(G22GAT), .Z(n369) );
  XOR2_X1 U406 ( .A(n369), .B(KEYINPUT72), .Z(n341) );
  XOR2_X1 U407 ( .A(G169GAT), .B(G8GAT), .Z(n413) );
  NAND2_X1 U408 ( .A1(G229GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U409 ( .A(n343), .B(n342), .ZN(n350) );
  XOR2_X1 U410 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n345) );
  XNOR2_X1 U411 ( .A(G43GAT), .B(G29GAT), .ZN(n344) );
  XNOR2_X1 U412 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U413 ( .A(KEYINPUT71), .B(n346), .ZN(n388) );
  XOR2_X1 U414 ( .A(KEYINPUT67), .B(G15GAT), .Z(n348) );
  XNOR2_X1 U415 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n347) );
  INV_X1 U416 ( .A(n517), .ZN(n578) );
  NAND2_X1 U417 ( .A1(n461), .A2(n578), .ZN(n352) );
  XOR2_X1 U418 ( .A(KEYINPUT81), .B(G78GAT), .Z(n354) );
  XNOR2_X1 U419 ( .A(G71GAT), .B(G64GAT), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U421 ( .A(n355), .B(G155GAT), .Z(n358) );
  XNOR2_X1 U422 ( .A(G8GAT), .B(n356), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n373) );
  XOR2_X1 U424 ( .A(G211GAT), .B(n359), .Z(n361) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U427 ( .A(KEYINPUT79), .B(KEYINPUT82), .Z(n363) );
  XNOR2_X1 U428 ( .A(KEYINPUT12), .B(KEYINPUT83), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U430 ( .A(n365), .B(n364), .Z(n371) );
  XOR2_X1 U431 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n367) );
  XNOR2_X1 U432 ( .A(G183GAT), .B(KEYINPUT80), .ZN(n366) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U436 ( .A(n373), .B(n372), .Z(n585) );
  INV_X1 U437 ( .A(n585), .ZN(n494) );
  NAND2_X1 U438 ( .A1(n374), .A2(n494), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n375), .B(KEYINPUT115), .ZN(n391) );
  XNOR2_X1 U440 ( .A(G36GAT), .B(G190GAT), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n376), .B(G218GAT), .ZN(n407) );
  XOR2_X1 U442 ( .A(n407), .B(KEYINPUT76), .Z(n378) );
  XOR2_X1 U443 ( .A(G50GAT), .B(G162GAT), .Z(n445) );
  XNOR2_X1 U444 ( .A(n445), .B(KEYINPUT10), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n378), .B(n377), .ZN(n384) );
  NAND2_X1 U446 ( .A1(G232GAT), .A2(G233GAT), .ZN(n381) );
  XOR2_X1 U447 ( .A(n384), .B(n383), .Z(n390) );
  XOR2_X1 U448 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n386) );
  XNOR2_X1 U449 ( .A(KEYINPUT11), .B(KEYINPUT77), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U451 ( .A(n388), .B(n387), .Z(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n571) );
  NAND2_X1 U453 ( .A1(n391), .A2(n571), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n392), .B(KEYINPUT47), .ZN(n399) );
  INV_X1 U455 ( .A(KEYINPUT78), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n393), .B(n571), .ZN(n553) );
  NOR2_X1 U457 ( .A1(n589), .A2(n494), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n394), .B(KEYINPUT45), .ZN(n396) );
  INV_X1 U459 ( .A(n395), .ZN(n486) );
  NAND2_X1 U460 ( .A1(n396), .A2(n486), .ZN(n397) );
  NOR2_X1 U461 ( .A1(n578), .A2(n397), .ZN(n398) );
  NOR2_X1 U462 ( .A1(n399), .A2(n398), .ZN(n401) );
  XOR2_X1 U463 ( .A(KEYINPUT79), .B(G204GAT), .Z(n403) );
  NAND2_X1 U464 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n406) );
  XOR2_X1 U466 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n405) );
  XNOR2_X1 U467 ( .A(G197GAT), .B(G211GAT), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n452) );
  XOR2_X1 U469 ( .A(n406), .B(n452), .Z(n409) );
  XNOR2_X1 U470 ( .A(G92GAT), .B(n407), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U472 ( .A(n411), .B(n410), .Z(n415) );
  XOR2_X1 U473 ( .A(n413), .B(n412), .Z(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n533) );
  NOR2_X1 U475 ( .A1(n539), .A2(n533), .ZN(n417) );
  XNOR2_X1 U476 ( .A(KEYINPUT124), .B(KEYINPUT54), .ZN(n416) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(n440) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n423) );
  XOR2_X1 U479 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n419) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(G127GAT), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U482 ( .A(G85GAT), .B(G162GAT), .Z(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n439) );
  XOR2_X1 U485 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n425) );
  XNOR2_X1 U486 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U488 ( .A(G141GAT), .B(n426), .ZN(n457) );
  XNOR2_X1 U489 ( .A(G148GAT), .B(n457), .ZN(n429) );
  XNOR2_X1 U490 ( .A(G1GAT), .B(n427), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n437) );
  XOR2_X1 U492 ( .A(KEYINPUT4), .B(KEYINPUT96), .Z(n431) );
  XNOR2_X1 U493 ( .A(G57GAT), .B(KEYINPUT95), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U495 ( .A(KEYINPUT1), .B(KEYINPUT94), .Z(n433) );
  XNOR2_X1 U496 ( .A(G120GAT), .B(KEYINPUT6), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U498 ( .A(n435), .B(n434), .Z(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n531) );
  NAND2_X1 U501 ( .A1(n440), .A2(n531), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n441), .B(KEYINPUT64), .ZN(n577) );
  XOR2_X1 U503 ( .A(KEYINPUT93), .B(KEYINPUT22), .Z(n443) );
  XNOR2_X1 U504 ( .A(G106GAT), .B(G218GAT), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U506 ( .A(n444), .B(KEYINPUT23), .Z(n447) );
  XNOR2_X1 U507 ( .A(G22GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n456) );
  XOR2_X1 U509 ( .A(KEYINPUT92), .B(KEYINPUT89), .Z(n449) );
  NAND2_X1 U510 ( .A1(G228GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U511 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U512 ( .A(n450), .B(KEYINPUT24), .Z(n454) );
  XNOR2_X1 U513 ( .A(n451), .B(n452), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(n475) );
  NOR2_X1 U517 ( .A1(n577), .A2(n475), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT55), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n461), .B(KEYINPUT110), .ZN(n547) );
  NAND2_X1 U520 ( .A1(n574), .A2(n547), .ZN(n465) );
  XOR2_X1 U521 ( .A(G176GAT), .B(KEYINPUT57), .Z(n463) );
  XOR2_X1 U522 ( .A(KEYINPUT56), .B(KEYINPUT125), .Z(n462) );
  XNOR2_X1 U523 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  INV_X1 U525 ( .A(KEYINPUT37), .ZN(n485) );
  NOR2_X1 U526 ( .A1(n533), .A2(n545), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n475), .A2(n466), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n467), .B(KEYINPUT25), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n533), .B(KEYINPUT27), .ZN(n473) );
  OR2_X1 U530 ( .A1(n473), .A2(n576), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n470), .A2(n469), .ZN(n471) );
  XOR2_X1 U532 ( .A(KEYINPUT101), .B(n471), .Z(n472) );
  NAND2_X1 U533 ( .A1(n472), .A2(n531), .ZN(n480) );
  NOR2_X1 U534 ( .A1(n531), .A2(n473), .ZN(n541) );
  XOR2_X1 U535 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(n543) );
  NAND2_X1 U537 ( .A1(n541), .A2(n543), .ZN(n476) );
  XOR2_X1 U538 ( .A(KEYINPUT98), .B(n476), .Z(n477) );
  NAND2_X1 U539 ( .A1(n477), .A2(n545), .ZN(n478) );
  XOR2_X1 U540 ( .A(KEYINPUT99), .B(n478), .Z(n479) );
  NAND2_X1 U541 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(KEYINPUT102), .ZN(n496) );
  NAND2_X1 U543 ( .A1(n496), .A2(n494), .ZN(n482) );
  XOR2_X1 U544 ( .A(KEYINPUT107), .B(n482), .Z(n483) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(n530) );
  NAND2_X1 U546 ( .A1(n486), .A2(n578), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n487), .B(KEYINPUT75), .ZN(n498) );
  NAND2_X1 U548 ( .A1(n530), .A2(n498), .ZN(n488) );
  NOR2_X1 U549 ( .A1(n514), .A2(n545), .ZN(n491) );
  NAND2_X1 U550 ( .A1(n574), .A2(n553), .ZN(n493) );
  NOR2_X1 U551 ( .A1(n553), .A2(n494), .ZN(n495) );
  XNOR2_X1 U552 ( .A(KEYINPUT16), .B(n495), .ZN(n497) );
  AND2_X1 U553 ( .A1(n497), .A2(n496), .ZN(n519) );
  NAND2_X1 U554 ( .A1(n498), .A2(n519), .ZN(n499) );
  XOR2_X1 U555 ( .A(KEYINPUT103), .B(n499), .Z(n507) );
  NOR2_X1 U556 ( .A1(n531), .A2(n507), .ZN(n500) );
  XOR2_X1 U557 ( .A(G1GAT), .B(n500), .Z(n501) );
  XNOR2_X1 U558 ( .A(KEYINPUT34), .B(n501), .ZN(G1324GAT) );
  NOR2_X1 U559 ( .A1(n533), .A2(n507), .ZN(n502) );
  XOR2_X1 U560 ( .A(G8GAT), .B(n502), .Z(G1325GAT) );
  NOR2_X1 U561 ( .A1(n507), .A2(n545), .ZN(n506) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n504) );
  XNOR2_X1 U563 ( .A(G15GAT), .B(KEYINPUT105), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n506), .B(n505), .ZN(G1326GAT) );
  NOR2_X1 U566 ( .A1(n543), .A2(n507), .ZN(n508) );
  XOR2_X1 U567 ( .A(G22GAT), .B(n508), .Z(G1327GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n510) );
  XNOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT108), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n510), .B(n509), .ZN(n512) );
  NOR2_X1 U571 ( .A1(n514), .A2(n531), .ZN(n511) );
  XOR2_X1 U572 ( .A(n512), .B(n511), .Z(G1328GAT) );
  NOR2_X1 U573 ( .A1(n533), .A2(n514), .ZN(n513) );
  XOR2_X1 U574 ( .A(G36GAT), .B(n513), .Z(G1329GAT) );
  XNOR2_X1 U575 ( .A(G50GAT), .B(KEYINPUT109), .ZN(n516) );
  NOR2_X1 U576 ( .A1(n543), .A2(n514), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n516), .B(n515), .ZN(G1331GAT) );
  NAND2_X1 U578 ( .A1(n547), .A2(n517), .ZN(n518) );
  XNOR2_X1 U579 ( .A(n518), .B(KEYINPUT111), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n529), .A2(n519), .ZN(n526) );
  NOR2_X1 U581 ( .A1(n531), .A2(n526), .ZN(n521) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(KEYINPUT112), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U584 ( .A(G57GAT), .B(n522), .Z(G1332GAT) );
  NOR2_X1 U585 ( .A1(n533), .A2(n526), .ZN(n524) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(KEYINPUT113), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(G1333GAT) );
  NOR2_X1 U588 ( .A1(n545), .A2(n526), .ZN(n525) );
  XOR2_X1 U589 ( .A(G71GAT), .B(n525), .Z(G1334GAT) );
  NOR2_X1 U590 ( .A1(n543), .A2(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1335GAT) );
  NAND2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n536) );
  NOR2_X1 U594 ( .A1(n531), .A2(n536), .ZN(n532) );
  XOR2_X1 U595 ( .A(G85GAT), .B(n532), .Z(G1336GAT) );
  NOR2_X1 U596 ( .A1(n533), .A2(n536), .ZN(n534) );
  XOR2_X1 U597 ( .A(G92GAT), .B(n534), .Z(G1337GAT) );
  NOR2_X1 U598 ( .A1(n545), .A2(n536), .ZN(n535) );
  XOR2_X1 U599 ( .A(G99GAT), .B(n535), .Z(G1338GAT) );
  NOR2_X1 U600 ( .A1(n543), .A2(n536), .ZN(n537) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(n537), .Z(n538) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U604 ( .A(KEYINPUT117), .B(n542), .ZN(n559) );
  NAND2_X1 U605 ( .A1(n543), .A2(n559), .ZN(n544) );
  NOR2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n554) );
  NAND2_X1 U607 ( .A1(n578), .A2(n554), .ZN(n546) );
  XNOR2_X1 U608 ( .A(n546), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(G120GAT), .B(KEYINPUT49), .Z(n549) );
  NAND2_X1 U610 ( .A1(n554), .A2(n547), .ZN(n548) );
  XNOR2_X1 U611 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n551) );
  NAND2_X1 U613 ( .A1(n554), .A2(n585), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n552), .Z(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT120), .Z(n557) );
  XNOR2_X1 U620 ( .A(n558), .B(n557), .ZN(G1343GAT) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(KEYINPUT122), .ZN(n563) );
  INV_X1 U622 ( .A(n576), .ZN(n560) );
  NAND2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT121), .B(n561), .Z(n570) );
  INV_X1 U625 ( .A(n570), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n568), .A2(n578), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n565) );
  NAND2_X1 U629 ( .A1(n568), .A2(n461), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT123), .Z(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n585), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U636 ( .A(G162GAT), .B(n572), .Z(G1347GAT) );
  NAND2_X1 U637 ( .A1(n578), .A2(n574), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n585), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n587) );
  NAND2_X1 U643 ( .A1(n587), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U647 ( .A1(n587), .A2(n395), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n587), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U652 ( .A(n587), .ZN(n588) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

