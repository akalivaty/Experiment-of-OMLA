//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n451, new_n453, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n599, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n647, new_n648, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT69), .Z(G217));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT70), .B(KEYINPUT2), .Z(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NAND2_X1  g036(.A1(new_n457), .A2(G2106), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n475), .A2(G137), .B1(G101), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n469), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n475), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n481), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(KEYINPUT71), .A2(G138), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n481), .B(new_n489), .C1(new_n467), .C2(new_n468), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n481), .A4(new_n489), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n493), .A2(G126), .A3(G2105), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n481), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n492), .A2(new_n494), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n502), .A2(KEYINPUT72), .A3(G651), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT72), .B1(new_n502), .B2(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XOR2_X1   g080(.A(KEYINPUT75), .B(G88), .Z(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT74), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT73), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n507), .B(KEYINPUT5), .C1(new_n508), .C2(KEYINPUT74), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n506), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G50), .A2(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n505), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n512), .A2(G62), .A3(new_n513), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n500), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(G166));
  NAND2_X1  g095(.A1(new_n512), .A2(new_n513), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n505), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT79), .B(G89), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n505), .A2(KEYINPUT76), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n502), .A2(G651), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n530), .B1(new_n500), .B2(KEYINPUT6), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n502), .A2(KEYINPUT72), .A3(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT77), .B(G51), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n528), .A2(G543), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G543), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n539), .A2(new_n507), .B1(KEYINPUT5), .B2(new_n510), .ZN(new_n540));
  INV_X1    g115(.A(new_n513), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n542), .A2(G63), .A3(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT78), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n537), .A2(KEYINPUT78), .A3(new_n543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n527), .B1(new_n546), .B2(new_n547), .ZN(G168));
  AOI21_X1  g123(.A(new_n508), .B1(new_n505), .B2(KEYINPUT76), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n549), .A2(G52), .A3(new_n535), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n512), .A2(G64), .A3(new_n513), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  XOR2_X1   g129(.A(KEYINPUT80), .B(G90), .Z(new_n555));
  NAND2_X1  g130(.A1(new_n522), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n550), .A2(new_n554), .A3(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n521), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n522), .A2(G81), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n528), .A2(G543), .A3(new_n535), .ZN(new_n565));
  INV_X1    g140(.A(G43), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT81), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  AND2_X1   g149(.A1(new_n522), .A2(G91), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT9), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(G543), .B1(new_n533), .B2(new_n534), .ZN(new_n578));
  AOI211_X1 g153(.A(KEYINPUT76), .B(new_n529), .C1(new_n531), .C2(new_n532), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n580), .A2(new_n581), .A3(G53), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n575), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(KEYINPUT73), .B2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT73), .B1(new_n538), .B2(G543), .ZN(new_n586));
  OAI211_X1 g161(.A(KEYINPUT82), .B(new_n513), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT82), .B1(new_n512), .B2(new_n513), .ZN(new_n589));
  OAI21_X1  g164(.A(G65), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G78), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n500), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT83), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI211_X1 g169(.A(KEYINPUT83), .B(new_n500), .C1(new_n590), .C2(new_n591), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n583), .B1(new_n594), .B2(new_n595), .ZN(G299));
  INV_X1    g171(.A(new_n527), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n537), .A2(KEYINPUT78), .A3(new_n543), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT78), .B1(new_n537), .B2(new_n543), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(G286));
  INV_X1    g175(.A(G166), .ZN(G303));
  OR2_X1    g176(.A1(new_n542), .A2(G74), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G87), .B2(new_n522), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n580), .A2(G49), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G288));
  NAND3_X1  g180(.A1(new_n512), .A2(G61), .A3(new_n513), .ZN(new_n606));
  NAND2_X1  g181(.A1(G73), .A2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n500), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n512), .A2(G86), .A3(new_n513), .ZN(new_n610));
  NAND2_X1  g185(.A1(G48), .A2(G543), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n533), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(G305));
  NAND2_X1  g189(.A1(G72), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G60), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n521), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G651), .B1(new_n522), .B2(G85), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n580), .A2(G47), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(G290));
  NAND2_X1  g195(.A1(G301), .A2(G868), .ZN(new_n621));
  NAND4_X1  g196(.A1(new_n533), .A2(G92), .A3(new_n512), .A4(new_n513), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(KEYINPUT84), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n542), .A2(new_n624), .A3(G92), .A4(new_n533), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT10), .ZN(new_n627));
  OAI21_X1  g202(.A(G66), .B1(new_n588), .B2(new_n589), .ZN(new_n628));
  NAND2_X1  g203(.A1(G79), .A2(G543), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT85), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n500), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n549), .A2(G54), .A3(new_n535), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G66), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n540), .B2(new_n541), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n635), .B1(new_n637), .B2(new_n587), .ZN(new_n638));
  INV_X1    g213(.A(new_n630), .ZN(new_n639));
  OAI21_X1  g214(.A(G651), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n580), .A2(G54), .ZN(new_n641));
  AOI21_X1  g216(.A(KEYINPUT86), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n627), .B1(new_n634), .B2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n621), .B1(new_n644), .B2(G868), .ZN(G284));
  OAI21_X1  g220(.A(new_n621), .B1(new_n644), .B2(G868), .ZN(G321));
  INV_X1    g221(.A(G868), .ZN(new_n647));
  NAND2_X1  g222(.A1(G299), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(G168), .ZN(G297));
  OAI21_X1  g224(.A(new_n648), .B1(new_n647), .B2(G168), .ZN(G280));
  INV_X1    g225(.A(G559), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n644), .B1(new_n651), .B2(G860), .ZN(G148));
  OAI21_X1  g227(.A(new_n632), .B1(new_n631), .B2(new_n633), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n640), .A2(KEYINPUT86), .A3(new_n641), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n651), .A3(new_n627), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G868), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g233(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g234(.A1(new_n493), .A2(new_n477), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT12), .Z(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT13), .Z(new_n662));
  INV_X1    g237(.A(G2100), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n475), .A2(G135), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n481), .A2(G111), .ZN(new_n667));
  OAI21_X1  g242(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n668));
  INV_X1    g243(.A(G123), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n493), .A2(G2105), .ZN(new_n670));
  OAI221_X1 g245(.A(new_n666), .B1(new_n667), .B2(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G2096), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n664), .A2(new_n665), .A3(new_n672), .ZN(G156));
  INV_X1    g248(.A(KEYINPUT14), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2427), .B(G2438), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2430), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT15), .B(G2435), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n677), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2451), .B(G2454), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT16), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1341), .B(G1348), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2443), .B(G2446), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(G14), .A3(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G401));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2072), .B(G2078), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n691), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g269(.A(G2084), .B(G2090), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n692), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n690), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n694), .B(new_n696), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n695), .A2(new_n692), .A3(new_n690), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT18), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n698), .A2(new_n699), .A3(new_n695), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G2096), .B(G2100), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(G227));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1956), .B(G2474), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1961), .B(G1966), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1971), .B(G1976), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT19), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n712), .A2(new_n713), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n714), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n717), .A2(new_n718), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT20), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n724), .B1(new_n723), .B2(new_n726), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n711), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n729), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n731), .A2(new_n727), .A3(new_n710), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n709), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(G1981), .B(G1986), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n730), .A2(new_n732), .A3(new_n709), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n735), .ZN(new_n738));
  INV_X1    g313(.A(new_n736), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n733), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(G229));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(G21), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G286), .B2(G16), .ZN(new_n745));
  INV_X1    g320(.A(G1966), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G5), .A2(G16), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT98), .Z(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G301), .B2(new_n743), .ZN(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G29), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n671), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G28), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n753), .B1(new_n755), .B2(G28), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT97), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT31), .B(G11), .Z(new_n761));
  NOR4_X1   g336(.A1(new_n752), .A2(new_n754), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n745), .A2(new_n746), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n747), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(KEYINPUT99), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT91), .B(G16), .Z(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G19), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n568), .B2(new_n767), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(G1341), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n753), .A2(G35), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n487), .B2(G29), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT29), .B(G2090), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(G164), .A2(G29), .ZN(new_n775));
  OR2_X1    g350(.A1(G27), .A2(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(G2078), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND3_X1   g352(.A1(new_n775), .A2(G2078), .A3(new_n776), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n774), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n750), .A2(new_n751), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n769), .A2(G1341), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n770), .A2(new_n779), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n753), .A2(G33), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT25), .Z(new_n785));
  INV_X1    g360(.A(G139), .ZN(new_n786));
  INV_X1    g361(.A(new_n475), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(G115), .A2(G2104), .ZN(new_n789));
  INV_X1    g364(.A(G127), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n469), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n788), .B1(G2105), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n783), .B1(new_n792), .B2(new_n753), .ZN(new_n793));
  INV_X1    g368(.A(G2072), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n477), .A2(G105), .ZN(new_n796));
  INV_X1    g371(.A(G141), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n787), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT26), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G129), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n670), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G29), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n753), .A2(G32), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT27), .B(G1996), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT96), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n753), .A2(G26), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT28), .Z(new_n812));
  AOI22_X1  g387(.A1(new_n482), .A2(G128), .B1(G140), .B2(new_n475), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT94), .B1(G104), .B2(G2105), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(KEYINPUT94), .A2(G104), .A3(G2105), .ZN(new_n816));
  OAI221_X1 g391(.A(G2104), .B1(G116), .B2(new_n481), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT95), .B(G2067), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G34), .ZN(new_n822));
  AOI21_X1  g397(.A(G29), .B1(new_n822), .B2(KEYINPUT24), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(KEYINPUT24), .B2(new_n822), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n479), .B2(new_n753), .ZN(new_n825));
  INV_X1    g400(.A(G2084), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n807), .B1(new_n805), .B2(new_n806), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n826), .B2(new_n825), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n795), .A2(new_n810), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n743), .A2(G4), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n643), .B2(G16), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT93), .B(G1348), .Z(new_n834));
  AOI211_X1 g409(.A(new_n782), .B(new_n831), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n764), .A2(KEYINPUT99), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n833), .A2(new_n834), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n766), .A2(G20), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G299), .B2(G16), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G1956), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n841), .A2(G1956), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n837), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND4_X1   g419(.A1(new_n765), .A2(new_n835), .A3(new_n836), .A4(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n743), .A2(G23), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G288), .B2(G16), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT33), .B(G1976), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(G305), .A2(G16), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT92), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n743), .A2(G6), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT32), .B(G1981), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n767), .A2(G22), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G166), .B2(new_n767), .ZN(new_n859));
  INV_X1    g434(.A(G1971), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n856), .B1(new_n853), .B2(new_n854), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n849), .A2(new_n857), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT34), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  MUX2_X1   g440(.A(G24), .B(G290), .S(new_n767), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G1986), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n753), .A2(G25), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n482), .A2(G119), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n475), .A2(G131), .ZN(new_n870));
  OR2_X1    g445(.A1(G95), .A2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(G2104), .C1(G107), .C2(new_n481), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n868), .B1(new_n874), .B2(new_n753), .ZN(new_n875));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G1991), .Z(new_n876));
  XOR2_X1   g451(.A(new_n875), .B(new_n876), .Z(new_n877));
  NOR2_X1   g452(.A1(new_n867), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n863), .B2(KEYINPUT34), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT36), .B1(new_n865), .B2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n863), .A2(KEYINPUT34), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT36), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n881), .A2(new_n864), .A3(new_n882), .A4(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n845), .A2(new_n884), .ZN(G311));
  AND3_X1   g460(.A1(new_n845), .A2(new_n884), .A3(KEYINPUT101), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT101), .B1(new_n845), .B2(new_n884), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(G150));
  XOR2_X1   g463(.A(KEYINPUT102), .B(G55), .Z(new_n889));
  NAND3_X1  g464(.A1(new_n549), .A2(new_n535), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(G80), .A2(G543), .ZN(new_n891));
  INV_X1    g466(.A(G67), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n521), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G651), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n522), .A2(G93), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(G860), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT37), .Z(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n564), .B2(new_n567), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n580), .A2(G43), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n901), .A2(KEYINPUT103), .A3(new_n562), .A4(new_n563), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n902), .A3(new_n896), .ZN(new_n903));
  INV_X1    g478(.A(new_n896), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n568), .A2(new_n904), .A3(KEYINPUT103), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(KEYINPUT38), .Z(new_n907));
  NAND2_X1  g482(.A1(new_n644), .A2(G559), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT39), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT104), .ZN(new_n911));
  INV_X1    g486(.A(G860), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n909), .B2(KEYINPUT39), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n898), .B1(new_n911), .B2(new_n913), .ZN(G145));
  XNOR2_X1  g489(.A(new_n818), .B(G164), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(new_n792), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n792), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n804), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n804), .A3(new_n918), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n475), .A2(G142), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n481), .A2(G118), .ZN(new_n923));
  OAI21_X1  g498(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n924));
  INV_X1    g499(.A(G130), .ZN(new_n925));
  OAI221_X1 g500(.A(new_n922), .B1(new_n923), .B2(new_n924), .C1(new_n925), .C2(new_n670), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n661), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n661), .A2(new_n926), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(new_n873), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n873), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT105), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n920), .A2(new_n921), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n935));
  INV_X1    g510(.A(new_n932), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n935), .B1(new_n936), .B2(new_n930), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n931), .A2(KEYINPUT105), .A3(new_n932), .ZN(new_n938));
  INV_X1    g513(.A(new_n918), .ZN(new_n939));
  INV_X1    g514(.A(new_n804), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(new_n916), .A3(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n937), .B(new_n938), .C1(new_n919), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n934), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(G160), .B(new_n671), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(G162), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT106), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n934), .A2(new_n942), .A3(new_n948), .A4(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n945), .B(KEYINPUT107), .ZN(new_n951));
  AOI21_X1  g526(.A(G37), .B1(new_n943), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g529(.A(new_n656), .B(new_n906), .Z(new_n955));
  INV_X1    g530(.A(KEYINPUT41), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n643), .A2(G299), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n592), .A2(new_n593), .ZN(new_n958));
  INV_X1    g533(.A(G65), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n637), .B2(new_n587), .ZN(new_n960));
  INV_X1    g535(.A(new_n591), .ZN(new_n961));
  OAI21_X1  g536(.A(G651), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT83), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n655), .A2(new_n627), .B1(new_n964), .B2(new_n583), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n956), .B1(new_n957), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n643), .A2(G299), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n655), .A2(new_n964), .A3(new_n583), .A4(new_n627), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(KEYINPUT41), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n955), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n656), .B(new_n906), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(KEYINPUT108), .A3(new_n968), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT108), .B1(new_n967), .B2(new_n968), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n976), .B1(new_n970), .B2(new_n975), .ZN(new_n979));
  NAND2_X1  g554(.A1(G288), .A2(G290), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n603), .A2(new_n604), .A3(new_n619), .A4(new_n618), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(G303), .B(G305), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n981), .B1(new_n980), .B2(new_n982), .ZN(new_n986));
  MUX2_X1   g561(.A(new_n985), .B(new_n984), .S(new_n986), .Z(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n978), .A2(new_n979), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n970), .A2(new_n975), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT42), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n987), .B1(new_n991), .B2(new_n977), .ZN(new_n992));
  OAI21_X1  g567(.A(G868), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n896), .A2(new_n647), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(G295));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n994), .ZN(G331));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n998));
  NAND2_X1  g573(.A1(G301), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n550), .A2(new_n554), .A3(new_n556), .A4(KEYINPUT110), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(G168), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n597), .B(new_n1000), .C1(new_n598), .C2(new_n599), .ZN(new_n1002));
  INV_X1    g577(.A(new_n999), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n906), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n546), .A2(new_n547), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1007), .A2(new_n597), .A3(new_n1000), .A4(new_n999), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1006), .A2(new_n1008), .A3(new_n905), .A4(new_n903), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(new_n966), .A3(new_n969), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1005), .A2(new_n967), .A3(new_n1009), .A4(new_n968), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n987), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G37), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1009), .B(new_n1005), .C1(new_n973), .C2(new_n974), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n987), .B1(new_n1016), .B2(new_n1011), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n997), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1010), .A2(new_n966), .A3(new_n969), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n957), .B2(new_n965), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1010), .B1(new_n1021), .B2(new_n972), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n988), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1023), .A2(KEYINPUT111), .A3(new_n1014), .A4(new_n1013), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1018), .A2(new_n1024), .A3(KEYINPUT43), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n987), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1015), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1027), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1029), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1015), .A2(new_n1017), .A3(KEYINPUT43), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1026), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1031), .A2(new_n1036), .ZN(G397));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(G1384), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n498), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n498), .B2(new_n1039), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n472), .A2(G40), .A3(new_n478), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n498), .A2(new_n1039), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n1039), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1042), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G2078), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT53), .ZN(new_n1051));
  OAI22_X1  g626(.A1(new_n1043), .A2(G1961), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n1053));
  AND4_X1   g628(.A1(new_n1053), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1053), .B1(new_n1055), .B2(new_n1047), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1050), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1052), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT125), .B1(new_n1059), .B2(G301), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n1059), .B2(G301), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT125), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1049), .A2(KEYINPUT114), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1055), .A2(new_n1053), .A3(new_n1047), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT53), .B1(new_n1066), .B2(new_n1050), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1063), .B(G171), .C1(new_n1067), .C2(new_n1052), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1060), .A2(new_n1062), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(G8), .B1(new_n516), .B2(new_n519), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT55), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n498), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT117), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n498), .A2(new_n1075), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G2090), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1064), .A2(new_n1065), .A3(new_n860), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1072), .B1(new_n1083), .B2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(G8), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1043), .A2(new_n1080), .ZN(new_n1086));
  AOI211_X1 g661(.A(new_n1085), .B(new_n1071), .C1(new_n1082), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1976), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT52), .B1(G288), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1044), .A2(new_n1042), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(new_n1085), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n603), .A2(G1976), .A3(new_n604), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT52), .ZN(new_n1095));
  INV_X1    g670(.A(G1981), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n609), .A2(new_n613), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n505), .B1(new_n610), .B2(new_n611), .ZN(new_n1098));
  OAI21_X1  g673(.A(G1981), .B1(new_n608), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT49), .ZN(new_n1102));
  NAND3_X1  g677(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1091), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1093), .B(new_n1095), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1084), .A2(new_n1087), .A3(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1059), .A2(G301), .ZN(new_n1109));
  AOI211_X1 g684(.A(G171), .B(new_n1052), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1061), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1069), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G299), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n964), .A2(new_n583), .A3(new_n1114), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT56), .B(G2072), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1046), .A2(new_n1048), .A3(new_n1047), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1055), .A2(KEYINPUT121), .A3(new_n1047), .A4(new_n1119), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1122), .B(new_n1123), .C1(new_n1079), .C2(G1956), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1118), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(G1956), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1123), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1128), .A2(new_n1122), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1113), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1118), .A2(new_n1124), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1128), .A2(new_n1117), .A3(new_n1116), .A4(new_n1122), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT61), .ZN(new_n1133));
  INV_X1    g708(.A(G2067), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1090), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n834), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(new_n1043), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT60), .B1(new_n643), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1044), .A2(KEYINPUT50), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1139), .A2(new_n1048), .A3(new_n1073), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1140), .A2(new_n834), .B1(new_n1134), .B2(new_n1090), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n655), .B2(new_n627), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G1996), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1046), .A2(new_n1048), .A3(new_n1144), .A4(new_n1047), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT58), .B(G1341), .Z(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1044), .B2(new_n1042), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n568), .ZN(new_n1149));
  NOR2_X1   g724(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1141), .A2(new_n1152), .A3(new_n655), .A4(new_n627), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1154));
  NAND3_X1  g729(.A1(new_n1148), .A2(new_n568), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1143), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1130), .A2(new_n1133), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n643), .A2(new_n1141), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1129), .B1(new_n1132), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(G1966), .B1(new_n1055), .B2(new_n1047), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT119), .B(G2084), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1162), .A2(new_n1163), .B1(new_n1140), .B2(new_n1164), .ZN(new_n1165));
  AOI211_X1 g740(.A(KEYINPUT118), .B(G1966), .C1(new_n1055), .C2(new_n1047), .ZN(new_n1166));
  OAI211_X1 g741(.A(G8), .B(G286), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT51), .ZN(new_n1168));
  NAND2_X1  g743(.A1(G286), .A2(G8), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(G286), .A2(KEYINPUT124), .A3(G8), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(G8), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(KEYINPUT123), .B(G8), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1168), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT51), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1174), .A2(new_n1179), .A3(new_n1169), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1112), .A2(new_n1161), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1184), .A2(new_n1177), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1168), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1187), .A2(KEYINPUT62), .A3(new_n1180), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1189), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1097), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1194));
  NOR2_X1   g769(.A1(G288), .A2(G1976), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1091), .B(KEYINPUT116), .Z(new_n1197));
  INV_X1    g772(.A(new_n1087), .ZN(new_n1198));
  OAI22_X1  g773(.A1(new_n1196), .A2(new_n1197), .B1(new_n1198), .B2(new_n1107), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1087), .A2(new_n1107), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1084), .ZN(new_n1201));
  OAI211_X1 g776(.A(G8), .B(G168), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT63), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1085), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1200), .B(new_n1207), .C1(new_n1072), .C2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1199), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1183), .A2(new_n1192), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1046), .A2(new_n1042), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(G290), .A2(G1986), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1213), .B1(new_n1214), .B2(KEYINPUT112), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(KEYINPUT112), .B2(new_n1214), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1212), .A2(G1986), .A3(G290), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  XOR2_X1   g793(.A(new_n1218), .B(KEYINPUT113), .Z(new_n1219));
  XNOR2_X1  g794(.A(new_n804), .B(new_n1144), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n818), .B(new_n1134), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n873), .B(new_n876), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1213), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1219), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1211), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1213), .B1(new_n1221), .B2(new_n940), .ZN(new_n1228));
  OR3_X1    g803(.A1(new_n1213), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1229));
  OAI21_X1  g804(.A(KEYINPUT46), .B1(new_n1213), .B2(G1996), .ZN(new_n1230));
  AOI21_X1  g805(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g806(.A(new_n1231), .B(KEYINPUT47), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT48), .ZN(new_n1233));
  AND2_X1   g808(.A1(new_n1216), .A2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g809(.A1(new_n1216), .A2(new_n1233), .ZN(new_n1235));
  NOR3_X1   g810(.A1(new_n1234), .A2(new_n1235), .A3(new_n1225), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n874), .A2(new_n876), .ZN(new_n1237));
  OAI22_X1  g812(.A1(new_n1222), .A2(new_n1237), .B1(G2067), .B2(new_n818), .ZN(new_n1238));
  AOI211_X1 g813(.A(new_n1232), .B(new_n1236), .C1(new_n1212), .C2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1227), .A2(new_n1239), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1242));
  NOR2_X1   g816(.A1(G227), .A2(new_n464), .ZN(new_n1243));
  XNOR2_X1  g817(.A(new_n1243), .B(KEYINPUT126), .ZN(new_n1244));
  NAND2_X1  g818(.A1(new_n1244), .A2(new_n688), .ZN(new_n1245));
  INV_X1    g819(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g820(.A(new_n1242), .B1(new_n741), .B2(new_n1246), .ZN(new_n1247));
  AOI211_X1 g821(.A(KEYINPUT127), .B(new_n1245), .C1(new_n737), .C2(new_n740), .ZN(new_n1248));
  OAI21_X1  g822(.A(new_n953), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NOR2_X1   g823(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1250));
  NOR2_X1   g824(.A1(new_n1249), .A2(new_n1250), .ZN(G308));
  OAI221_X1 g825(.A(new_n953), .B1(new_n1247), .B2(new_n1248), .C1(new_n1034), .C2(new_n1035), .ZN(G225));
endmodule


