

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758;

  AND2_X1 U368 ( .A1(n403), .A2(n404), .ZN(n367) );
  AND2_X1 U369 ( .A1(n378), .A2(n354), .ZN(n464) );
  XNOR2_X1 U370 ( .A(n344), .B(n475), .ZN(n640) );
  XNOR2_X1 U371 ( .A(n379), .B(n353), .ZN(n344) );
  XNOR2_X1 U372 ( .A(n396), .B(n431), .ZN(n430) );
  XNOR2_X1 U373 ( .A(n506), .B(n505), .ZN(n739) );
  XNOR2_X1 U374 ( .A(n466), .B(n509), .ZN(n725) );
  BUF_X1 U375 ( .A(G128), .Z(n653) );
  NOR2_X1 U376 ( .A1(n605), .A2(n685), .ZN(n606) );
  XNOR2_X2 U377 ( .A(n345), .B(KEYINPUT64), .ZN(n625) );
  NAND2_X2 U378 ( .A1(n462), .A2(n622), .ZN(n345) );
  INV_X1 U379 ( .A(G953), .ZN(n745) );
  XOR2_X1 U380 ( .A(n347), .B(n361), .Z(n346) );
  AND2_X2 U381 ( .A1(n388), .A2(n389), .ZN(n383) );
  AND2_X4 U382 ( .A1(n625), .A2(n358), .ZN(n718) );
  NOR2_X2 U383 ( .A1(n662), .A2(n648), .ZN(n618) );
  XNOR2_X2 U384 ( .A(n567), .B(KEYINPUT42), .ZN(n758) );
  NAND2_X2 U385 ( .A1(n405), .A2(n367), .ZN(n402) );
  AND2_X2 U386 ( .A1(n611), .A2(n349), .ZN(n652) );
  XNOR2_X2 U387 ( .A(n450), .B(n531), .ZN(n589) );
  XNOR2_X2 U388 ( .A(n473), .B(G119), .ZN(n396) );
  XNOR2_X2 U389 ( .A(n430), .B(n380), .ZN(n379) );
  INV_X1 U390 ( .A(n613), .ZN(n682) );
  AND2_X1 U391 ( .A1(n578), .A2(n574), .ZN(n659) );
  NOR2_X1 U392 ( .A1(n384), .A2(n383), .ZN(n454) );
  AND2_X1 U393 ( .A1(n386), .A2(n387), .ZN(n385) );
  AND2_X1 U394 ( .A1(n417), .A2(n415), .ZN(n414) );
  AND2_X1 U395 ( .A1(n378), .A2(n682), .ZN(n611) );
  BUF_X1 U396 ( .A(n560), .Z(n685) );
  NOR2_X2 U397 ( .A1(n709), .A2(G902), .ZN(n511) );
  OR2_X1 U398 ( .A1(n626), .A2(G902), .ZN(n447) );
  XNOR2_X1 U399 ( .A(n526), .B(n457), .ZN(n740) );
  XNOR2_X1 U400 ( .A(n399), .B(G146), .ZN(n526) );
  XNOR2_X1 U401 ( .A(KEYINPUT68), .B(G101), .ZN(n510) );
  BUF_X1 U402 ( .A(n401), .Z(n347) );
  NAND2_X1 U403 ( .A1(n377), .A2(n671), .ZN(n401) );
  XNOR2_X1 U404 ( .A(n602), .B(n362), .ZN(n378) );
  NOR2_X1 U405 ( .A1(n461), .A2(n601), .ZN(n602) );
  XNOR2_X2 U406 ( .A(n725), .B(n465), .ZN(n527) );
  INV_X1 U407 ( .A(G125), .ZN(n399) );
  XNOR2_X1 U408 ( .A(G131), .B(G134), .ZN(n489) );
  XOR2_X1 U409 ( .A(G902), .B(KEYINPUT15), .Z(n621) );
  XNOR2_X1 U410 ( .A(n510), .B(KEYINPUT71), .ZN(n465) );
  INV_X1 U411 ( .A(KEYINPUT38), .ZN(n443) );
  XNOR2_X1 U412 ( .A(n688), .B(KEYINPUT6), .ZN(n610) );
  INV_X1 U413 ( .A(n561), .ZN(n468) );
  XNOR2_X1 U414 ( .A(n554), .B(n553), .ZN(n631) );
  XNOR2_X1 U415 ( .A(n458), .B(n740), .ZN(n554) );
  XNOR2_X1 U416 ( .A(KEYINPUT11), .B(KEYINPUT96), .ZN(n460) );
  XNOR2_X1 U417 ( .A(KEYINPUT97), .B(KEYINPUT12), .ZN(n545) );
  XNOR2_X1 U418 ( .A(G143), .B(G131), .ZN(n547) );
  XOR2_X1 U419 ( .A(G146), .B(G107), .Z(n508) );
  XNOR2_X2 U420 ( .A(KEYINPUT4), .B(KEYINPUT69), .ZN(n488) );
  INV_X1 U421 ( .A(KEYINPUT17), .ZN(n520) );
  XNOR2_X1 U422 ( .A(n522), .B(KEYINPUT78), .ZN(n474) );
  XNOR2_X1 U423 ( .A(n526), .B(n429), .ZN(n428) );
  AND2_X1 U424 ( .A1(n560), .A2(n684), .ZN(n382) );
  INV_X1 U425 ( .A(n610), .ZN(n434) );
  INV_X1 U426 ( .A(n535), .ZN(n380) );
  XNOR2_X1 U427 ( .A(n525), .B(KEYINPUT16), .ZN(n431) );
  XNOR2_X1 U428 ( .A(G104), .B(KEYINPUT88), .ZN(n509) );
  XNOR2_X1 U429 ( .A(n408), .B(G110), .ZN(n466) );
  INV_X1 U430 ( .A(KEYINPUT75), .ZN(n408) );
  XNOR2_X1 U431 ( .A(G137), .B(G140), .ZN(n505) );
  XNOR2_X1 U432 ( .A(G475), .B(n557), .ZN(n578) );
  XNOR2_X1 U433 ( .A(n512), .B(G469), .ZN(n478) );
  XNOR2_X1 U434 ( .A(n675), .B(n455), .ZN(n619) );
  INV_X1 U435 ( .A(KEYINPUT81), .ZN(n455) );
  INV_X1 U436 ( .A(n619), .ZN(n435) );
  XNOR2_X1 U437 ( .A(n618), .B(n436), .ZN(n366) );
  INV_X1 U438 ( .A(KEYINPUT94), .ZN(n436) );
  NAND2_X1 U439 ( .A1(n413), .A2(n348), .ZN(n412) );
  INV_X1 U440 ( .A(KEYINPUT104), .ZN(n432) );
  NAND2_X1 U441 ( .A1(n611), .A2(n369), .ZN(n374) );
  AND2_X1 U442 ( .A1(n433), .A2(n432), .ZN(n369) );
  INV_X1 U443 ( .A(KEYINPUT18), .ZN(n429) );
  XNOR2_X1 U444 ( .A(n456), .B(KEYINPUT102), .ZN(n675) );
  NOR2_X1 U445 ( .A1(n661), .A2(n659), .ZN(n456) );
  XNOR2_X1 U446 ( .A(n395), .B(n484), .ZN(n487) );
  XNOR2_X1 U447 ( .A(G137), .B(KEYINPUT74), .ZN(n482) );
  INV_X1 U448 ( .A(KEYINPUT72), .ZN(n525) );
  XOR2_X1 U449 ( .A(KEYINPUT8), .B(n494), .Z(n538) );
  NAND2_X1 U450 ( .A1(n745), .A2(G234), .ZN(n494) );
  XOR2_X1 U451 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n533) );
  XNOR2_X1 U452 ( .A(G134), .B(KEYINPUT100), .ZN(n532) );
  XNOR2_X1 U453 ( .A(n524), .B(G122), .ZN(n535) );
  XNOR2_X1 U454 ( .A(G116), .B(G107), .ZN(n524) );
  NOR2_X1 U455 ( .A1(G953), .A2(G237), .ZN(n551) );
  XNOR2_X1 U456 ( .A(n548), .B(n459), .ZN(n458) );
  XNOR2_X1 U457 ( .A(n545), .B(n460), .ZN(n459) );
  INV_X1 U458 ( .A(KEYINPUT95), .ZN(n546) );
  XNOR2_X1 U459 ( .A(G113), .B(G104), .ZN(n549) );
  XOR2_X1 U460 ( .A(G140), .B(G122), .Z(n550) );
  NAND2_X1 U461 ( .A1(G234), .A2(G237), .ZN(n513) );
  OR2_X1 U462 ( .A1(G237), .A2(G902), .ZN(n529) );
  BUF_X1 U463 ( .A(n624), .Z(n743) );
  INV_X1 U464 ( .A(KEYINPUT10), .ZN(n457) );
  XNOR2_X1 U465 ( .A(n394), .B(n653), .ZN(n393) );
  XNOR2_X1 U466 ( .A(KEYINPUT24), .B(G110), .ZN(n394) );
  XNOR2_X1 U467 ( .A(n441), .B(n392), .ZN(n391) );
  INV_X1 U468 ( .A(KEYINPUT23), .ZN(n441) );
  INV_X1 U469 ( .A(G119), .ZN(n392) );
  AND2_X1 U470 ( .A1(n624), .A2(n621), .ZN(n463) );
  XNOR2_X1 U471 ( .A(n527), .B(n350), .ZN(n451) );
  NOR2_X1 U472 ( .A1(n674), .A2(n376), .ZN(n566) );
  XNOR2_X1 U473 ( .A(n682), .B(KEYINPUT87), .ZN(n604) );
  INV_X1 U474 ( .A(KEYINPUT106), .ZN(n437) );
  XNOR2_X1 U475 ( .A(n608), .B(n607), .ZN(n668) );
  XNOR2_X1 U476 ( .A(n424), .B(n423), .ZN(n575) );
  INV_X1 U477 ( .A(KEYINPUT76), .ZN(n423) );
  INV_X1 U478 ( .A(n382), .ZN(n681) );
  NOR2_X1 U479 ( .A1(n434), .A2(n612), .ZN(n433) );
  XNOR2_X1 U480 ( .A(KEYINPUT86), .B(n627), .ZN(n628) );
  XNOR2_X1 U481 ( .A(n472), .B(n471), .ZN(n720) );
  XNOR2_X1 U482 ( .A(n740), .B(n505), .ZN(n471) );
  XNOR2_X1 U483 ( .A(n495), .B(n390), .ZN(n472) );
  XNOR2_X1 U484 ( .A(n393), .B(n391), .ZN(n390) );
  XNOR2_X1 U485 ( .A(n631), .B(KEYINPUT59), .ZN(n632) );
  XNOR2_X1 U486 ( .A(n558), .B(n559), .ZN(n470) );
  NOR2_X2 U487 ( .A1(n580), .A2(n346), .ZN(n657) );
  AND2_X1 U488 ( .A1(n611), .A2(n433), .ZN(n646) );
  INV_X1 U489 ( .A(KEYINPUT118), .ZN(n445) );
  BUF_X1 U490 ( .A(n755), .Z(n400) );
  AND2_X1 U491 ( .A1(n579), .A2(KEYINPUT80), .ZN(n348) );
  AND2_X1 U492 ( .A1(n603), .A2(n612), .ZN(n349) );
  XOR2_X1 U493 ( .A(n508), .B(n507), .Z(n350) );
  AND2_X1 U494 ( .A1(G214), .A2(n551), .ZN(n351) );
  AND2_X1 U495 ( .A1(n551), .A2(G210), .ZN(n352) );
  XOR2_X1 U496 ( .A(n474), .B(n428), .Z(n353) );
  XOR2_X1 U497 ( .A(n606), .B(KEYINPUT79), .Z(n354) );
  AND2_X1 U498 ( .A1(n578), .A2(n577), .ZN(n355) );
  AND2_X1 U499 ( .A1(G210), .A2(n529), .ZN(n356) );
  AND2_X1 U500 ( .A1(n591), .A2(n584), .ZN(n357) );
  NAND2_X1 U501 ( .A1(n670), .A2(KEYINPUT2), .ZN(n358) );
  AND2_X1 U502 ( .A1(n591), .A2(KEYINPUT48), .ZN(n359) );
  AND2_X1 U503 ( .A1(n435), .A2(n432), .ZN(n360) );
  XNOR2_X1 U504 ( .A(KEYINPUT19), .B(KEYINPUT66), .ZN(n361) );
  XOR2_X1 U505 ( .A(KEYINPUT65), .B(KEYINPUT22), .Z(n362) );
  XNOR2_X1 U506 ( .A(n715), .B(KEYINPUT117), .ZN(n363) );
  XOR2_X1 U507 ( .A(KEYINPUT85), .B(KEYINPUT63), .Z(n364) );
  NOR2_X1 U508 ( .A1(G952), .A2(n745), .ZN(n724) );
  AND2_X1 U509 ( .A1(n572), .A2(n468), .ZN(n467) );
  XNOR2_X1 U510 ( .A(n572), .B(KEYINPUT1), .ZN(n613) );
  XNOR2_X1 U511 ( .A(n426), .B(KEYINPUT77), .ZN(n425) );
  NAND2_X1 U512 ( .A1(n425), .A2(n427), .ZN(n424) );
  BUF_X1 U513 ( .A(n589), .Z(n365) );
  XNOR2_X1 U514 ( .A(n620), .B(KEYINPUT84), .ZN(n404) );
  XNOR2_X1 U515 ( .A(n401), .B(n361), .ZN(n597) );
  NAND2_X1 U516 ( .A1(n366), .A2(n360), .ZN(n368) );
  NAND2_X1 U517 ( .A1(n366), .A2(n435), .ZN(n371) );
  XNOR2_X2 U518 ( .A(n464), .B(KEYINPUT32), .ZN(n755) );
  AND2_X1 U519 ( .A1(n368), .A2(n374), .ZN(n373) );
  NAND2_X1 U520 ( .A1(n373), .A2(n370), .ZN(n403) );
  NAND2_X1 U521 ( .A1(n372), .A2(n371), .ZN(n370) );
  NOR2_X1 U522 ( .A1(n646), .A2(n432), .ZN(n372) );
  INV_X1 U523 ( .A(n375), .ZN(n411) );
  NAND2_X1 U524 ( .A1(n454), .A2(n452), .ZN(n375) );
  NAND2_X1 U525 ( .A1(n375), .A2(n357), .ZN(n409) );
  NOR2_X1 U526 ( .A1(n675), .A2(n376), .ZN(n676) );
  NAND2_X1 U527 ( .A1(n672), .A2(n671), .ZN(n376) );
  XNOR2_X1 U528 ( .A(n377), .B(n443), .ZN(n672) );
  AND2_X1 U529 ( .A1(n575), .A2(n377), .ZN(n576) );
  NOR2_X1 U530 ( .A1(n588), .A2(n377), .ZN(n667) );
  XNOR2_X2 U531 ( .A(n530), .B(n356), .ZN(n377) );
  XNOR2_X1 U532 ( .A(n379), .B(KEYINPUT122), .ZN(n727) );
  NAND2_X1 U533 ( .A1(n467), .A2(n382), .ZN(n426) );
  NOR2_X1 U534 ( .A1(n681), .A2(n381), .ZN(n469) );
  INV_X1 U535 ( .A(n572), .ZN(n381) );
  AND2_X1 U536 ( .A1(n613), .A2(n382), .ZN(n614) );
  NAND2_X1 U537 ( .A1(n385), .A2(n665), .ZN(n384) );
  NAND2_X1 U538 ( .A1(n752), .A2(KEYINPUT46), .ZN(n386) );
  NAND2_X1 U539 ( .A1(n758), .A2(KEYINPUT46), .ZN(n387) );
  NOR2_X1 U540 ( .A1(n752), .A2(KEYINPUT46), .ZN(n388) );
  INV_X1 U541 ( .A(n758), .ZN(n389) );
  XNOR2_X2 U542 ( .A(n449), .B(n470), .ZN(n752) );
  INV_X1 U543 ( .A(n396), .ZN(n395) );
  XNOR2_X1 U544 ( .A(n609), .B(n397), .ZN(n407) );
  INV_X1 U545 ( .A(KEYINPUT44), .ZN(n397) );
  NOR2_X2 U546 ( .A1(n755), .A2(n652), .ZN(n609) );
  NAND2_X1 U547 ( .A1(n398), .A2(n355), .ZN(n476) );
  XNOR2_X1 U548 ( .A(n477), .B(KEYINPUT34), .ZN(n398) );
  XNOR2_X1 U549 ( .A(n739), .B(n451), .ZN(n709) );
  NAND2_X1 U550 ( .A1(n575), .A2(n672), .ZN(n450) );
  NAND2_X1 U551 ( .A1(n589), .A2(n659), .ZN(n449) );
  NOR2_X1 U552 ( .A1(n696), .A2(n580), .ZN(n567) );
  XNOR2_X1 U553 ( .A(n566), .B(KEYINPUT41), .ZN(n696) );
  NOR2_X1 U554 ( .A1(n461), .A2(n668), .ZN(n477) );
  NAND2_X1 U555 ( .A1(n410), .A2(n409), .ZN(n624) );
  NOR2_X1 U556 ( .A1(n570), .A2(n347), .ZN(n571) );
  XNOR2_X1 U557 ( .A(n453), .B(KEYINPUT73), .ZN(n452) );
  XNOR2_X2 U558 ( .A(n402), .B(KEYINPUT45), .ZN(n733) );
  NAND2_X1 U559 ( .A1(n407), .A2(n406), .ZN(n405) );
  NAND2_X1 U560 ( .A1(n609), .A2(n756), .ZN(n406) );
  NAND2_X1 U561 ( .A1(n411), .A2(n359), .ZN(n410) );
  NAND2_X1 U562 ( .A1(n422), .A2(n355), .ZN(n656) );
  NAND2_X1 U563 ( .A1(n414), .A2(n412), .ZN(n480) );
  INV_X1 U564 ( .A(n422), .ZN(n413) );
  NAND2_X1 U565 ( .A1(n422), .A2(n416), .ZN(n415) );
  AND2_X1 U566 ( .A1(n355), .A2(n481), .ZN(n416) );
  NAND2_X1 U567 ( .A1(n420), .A2(n418), .ZN(n417) );
  NAND2_X1 U568 ( .A1(n579), .A2(n419), .ZN(n418) );
  OR2_X1 U569 ( .A1(n355), .A2(n481), .ZN(n419) );
  NAND2_X1 U570 ( .A1(n421), .A2(KEYINPUT80), .ZN(n420) );
  INV_X1 U571 ( .A(n579), .ZN(n421) );
  XNOR2_X1 U572 ( .A(n576), .B(KEYINPUT108), .ZN(n422) );
  INV_X1 U573 ( .A(n519), .ZN(n427) );
  XNOR2_X2 U574 ( .A(n599), .B(KEYINPUT0), .ZN(n461) );
  XNOR2_X1 U575 ( .A(n438), .B(n437), .ZN(n586) );
  AND2_X1 U576 ( .A1(n569), .A2(n659), .ZN(n438) );
  BUF_X1 U577 ( .A(n662), .Z(n439) );
  NAND2_X1 U578 ( .A1(n733), .A2(n463), .ZN(n440) );
  XNOR2_X1 U579 ( .A(n440), .B(KEYINPUT82), .ZN(n462) );
  NOR2_X1 U580 ( .A1(n720), .A2(G902), .ZN(n501) );
  XNOR2_X1 U581 ( .A(n444), .B(n645), .ZN(G51) );
  NAND2_X1 U582 ( .A1(n643), .A2(n644), .ZN(n444) );
  NAND2_X1 U583 ( .A1(n597), .A2(n598), .ZN(n599) );
  XNOR2_X1 U584 ( .A(n446), .B(n445), .ZN(G63) );
  NAND2_X1 U585 ( .A1(n717), .A2(n644), .ZN(n446) );
  XNOR2_X2 U586 ( .A(n447), .B(G472), .ZN(n688) );
  XNOR2_X1 U587 ( .A(n448), .B(n364), .ZN(G57) );
  NAND2_X1 U588 ( .A1(n630), .A2(n644), .ZN(n448) );
  NAND2_X1 U589 ( .A1(n434), .A2(n614), .ZN(n608) );
  XNOR2_X2 U590 ( .A(n521), .B(n489), .ZN(n506) );
  NAND2_X1 U591 ( .A1(n583), .A2(n480), .ZN(n453) );
  NOR2_X1 U592 ( .A1(n461), .A2(n691), .ZN(n616) );
  NOR2_X1 U593 ( .A1(n461), .A2(n617), .ZN(n648) );
  XNOR2_X1 U594 ( .A(n527), .B(n523), .ZN(n475) );
  NAND2_X1 U595 ( .A1(n469), .A2(n603), .ZN(n617) );
  XNOR2_X2 U596 ( .A(G113), .B(KEYINPUT3), .ZN(n473) );
  XNOR2_X2 U597 ( .A(n476), .B(KEYINPUT35), .ZN(n756) );
  XNOR2_X2 U598 ( .A(n511), .B(n478), .ZN(n572) );
  XNOR2_X2 U599 ( .A(n479), .B(n536), .ZN(n521) );
  INV_X1 U600 ( .A(n488), .ZN(n479) );
  INV_X1 U601 ( .A(KEYINPUT80), .ZN(n481) );
  XNOR2_X1 U602 ( .A(n716), .B(n363), .ZN(n717) );
  XNOR2_X1 U603 ( .A(n352), .B(n485), .ZN(n486) );
  XNOR2_X1 U604 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U605 ( .A(n487), .B(n486), .ZN(n491) );
  XNOR2_X1 U606 ( .A(n552), .B(n351), .ZN(n553) );
  BUF_X1 U607 ( .A(n668), .Z(n680) );
  INV_X1 U608 ( .A(KEYINPUT109), .ZN(n559) );
  XNOR2_X1 U609 ( .A(n501), .B(n500), .ZN(n560) );
  XNOR2_X1 U610 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U611 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U612 ( .A(n638), .B(n637), .ZN(G60) );
  INV_X1 U613 ( .A(n724), .ZN(n644) );
  XOR2_X1 U614 ( .A(KEYINPUT30), .B(KEYINPUT107), .Z(n493) );
  XOR2_X1 U615 ( .A(G116), .B(KEYINPUT5), .Z(n483) );
  XNOR2_X1 U616 ( .A(n483), .B(n482), .ZN(n484) );
  INV_X1 U617 ( .A(n510), .ZN(n485) );
  XNOR2_X2 U618 ( .A(G143), .B(G128), .ZN(n536) );
  XNOR2_X1 U619 ( .A(n506), .B(G146), .ZN(n490) );
  XNOR2_X1 U620 ( .A(n491), .B(n490), .ZN(n626) );
  NAND2_X1 U621 ( .A1(G214), .A2(n529), .ZN(n671) );
  NAND2_X1 U622 ( .A1(n688), .A2(n671), .ZN(n492) );
  XNOR2_X1 U623 ( .A(n493), .B(n492), .ZN(n519) );
  NAND2_X1 U624 ( .A1(n538), .A2(G221), .ZN(n495) );
  XOR2_X1 U625 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n499) );
  INV_X1 U626 ( .A(n621), .ZN(n528) );
  NAND2_X1 U627 ( .A1(n528), .A2(G234), .ZN(n496) );
  XNOR2_X1 U628 ( .A(n496), .B(KEYINPUT20), .ZN(n497) );
  XNOR2_X1 U629 ( .A(KEYINPUT90), .B(n497), .ZN(n502) );
  NAND2_X1 U630 ( .A1(G217), .A2(n502), .ZN(n498) );
  XNOR2_X1 U631 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U632 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n504) );
  NAND2_X1 U633 ( .A1(G221), .A2(n502), .ZN(n503) );
  XNOR2_X1 U634 ( .A(n504), .B(n503), .ZN(n684) );
  INV_X1 U635 ( .A(KEYINPUT70), .ZN(n512) );
  NAND2_X1 U636 ( .A1(G227), .A2(n745), .ZN(n507) );
  XNOR2_X1 U637 ( .A(n513), .B(KEYINPUT14), .ZN(n515) );
  NAND2_X1 U638 ( .A1(G952), .A2(n515), .ZN(n514) );
  XOR2_X1 U639 ( .A(KEYINPUT89), .B(n514), .Z(n702) );
  NOR2_X1 U640 ( .A1(G953), .A2(n702), .ZN(n592) );
  NAND2_X1 U641 ( .A1(G902), .A2(n515), .ZN(n593) );
  NOR2_X1 U642 ( .A1(G900), .A2(n593), .ZN(n516) );
  NAND2_X1 U643 ( .A1(G953), .A2(n516), .ZN(n517) );
  XNOR2_X1 U644 ( .A(KEYINPUT105), .B(n517), .ZN(n518) );
  NOR2_X1 U645 ( .A1(n592), .A2(n518), .ZN(n561) );
  XNOR2_X1 U646 ( .A(n521), .B(n520), .ZN(n523) );
  NAND2_X1 U647 ( .A1(G224), .A2(n745), .ZN(n522) );
  NAND2_X1 U648 ( .A1(n640), .A2(n528), .ZN(n530) );
  XOR2_X1 U649 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n531) );
  XNOR2_X1 U650 ( .A(KEYINPUT101), .B(G478), .ZN(n544) );
  XNOR2_X1 U651 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U652 ( .A(n535), .B(n534), .ZN(n542) );
  INV_X1 U653 ( .A(n536), .ZN(n537) );
  XOR2_X1 U654 ( .A(n537), .B(KEYINPUT7), .Z(n540) );
  NAND2_X1 U655 ( .A1(G217), .A2(n538), .ZN(n539) );
  XNOR2_X1 U656 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U657 ( .A(n542), .B(n541), .ZN(n715) );
  NOR2_X1 U658 ( .A1(G902), .A2(n715), .ZN(n543) );
  XNOR2_X1 U659 ( .A(n544), .B(n543), .ZN(n577) );
  INV_X1 U660 ( .A(n577), .ZN(n574) );
  XNOR2_X1 U661 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n556) );
  XNOR2_X1 U662 ( .A(n550), .B(n549), .ZN(n552) );
  NOR2_X1 U663 ( .A1(G902), .A2(n631), .ZN(n555) );
  XNOR2_X1 U664 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U665 ( .A(KEYINPUT40), .B(KEYINPUT110), .Z(n558) );
  NOR2_X1 U666 ( .A1(n561), .A2(n685), .ZN(n562) );
  NAND2_X1 U667 ( .A1(n684), .A2(n562), .ZN(n568) );
  INV_X1 U668 ( .A(n688), .ZN(n603) );
  NOR2_X1 U669 ( .A1(n568), .A2(n603), .ZN(n563) );
  XNOR2_X1 U670 ( .A(n563), .B(KEYINPUT28), .ZN(n564) );
  NAND2_X1 U671 ( .A1(n564), .A2(n572), .ZN(n580) );
  NOR2_X1 U672 ( .A1(n578), .A2(n577), .ZN(n565) );
  XNOR2_X1 U673 ( .A(n565), .B(KEYINPUT103), .ZN(n674) );
  NOR2_X1 U674 ( .A1(n610), .A2(n568), .ZN(n569) );
  XOR2_X1 U675 ( .A(n586), .B(KEYINPUT111), .Z(n570) );
  XNOR2_X1 U676 ( .A(KEYINPUT36), .B(n571), .ZN(n573) );
  NAND2_X1 U677 ( .A1(n573), .A2(n604), .ZN(n665) );
  NOR2_X1 U678 ( .A1(n574), .A2(n578), .ZN(n661) );
  NAND2_X1 U679 ( .A1(KEYINPUT47), .A2(n675), .ZN(n579) );
  XOR2_X1 U680 ( .A(n657), .B(KEYINPUT47), .Z(n582) );
  NAND2_X1 U681 ( .A1(n657), .A2(n619), .ZN(n581) );
  NAND2_X1 U682 ( .A1(n582), .A2(n581), .ZN(n583) );
  INV_X1 U683 ( .A(KEYINPUT48), .ZN(n584) );
  NAND2_X1 U684 ( .A1(n671), .A2(n682), .ZN(n585) );
  NOR2_X1 U685 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U686 ( .A(n587), .B(KEYINPUT43), .ZN(n588) );
  INV_X1 U687 ( .A(n667), .ZN(n590) );
  NAND2_X1 U688 ( .A1(n365), .A2(n661), .ZN(n666) );
  AND2_X1 U689 ( .A1(n590), .A2(n666), .ZN(n591) );
  INV_X1 U690 ( .A(n592), .ZN(n596) );
  INV_X1 U691 ( .A(n593), .ZN(n594) );
  NOR2_X1 U692 ( .A1(G898), .A2(n745), .ZN(n728) );
  NAND2_X1 U693 ( .A1(n594), .A2(n728), .ZN(n595) );
  NAND2_X1 U694 ( .A1(n596), .A2(n595), .ZN(n598) );
  INV_X1 U695 ( .A(n674), .ZN(n600) );
  NAND2_X1 U696 ( .A1(n684), .A2(n600), .ZN(n601) );
  NAND2_X1 U697 ( .A1(n604), .A2(n610), .ZN(n605) );
  INV_X1 U698 ( .A(KEYINPUT33), .ZN(n607) );
  INV_X1 U699 ( .A(n685), .ZN(n612) );
  NAND2_X1 U700 ( .A1(n688), .A2(n614), .ZN(n691) );
  XNOR2_X1 U701 ( .A(KEYINPUT93), .B(KEYINPUT31), .ZN(n615) );
  XNOR2_X1 U702 ( .A(n616), .B(n615), .ZN(n662) );
  NAND2_X1 U703 ( .A1(KEYINPUT44), .A2(n756), .ZN(n620) );
  NAND2_X1 U704 ( .A1(KEYINPUT2), .A2(n621), .ZN(n622) );
  AND2_X1 U705 ( .A1(n733), .A2(n743), .ZN(n670) );
  NAND2_X1 U706 ( .A1(n718), .A2(G472), .ZN(n629) );
  XOR2_X1 U707 ( .A(n626), .B(KEYINPUT62), .Z(n627) );
  XNOR2_X1 U708 ( .A(n629), .B(n628), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n718), .A2(G475), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n634), .A2(n644), .ZN(n638) );
  INV_X1 U712 ( .A(KEYINPUT67), .ZN(n636) );
  INV_X1 U713 ( .A(KEYINPUT60), .ZN(n635) );
  XNOR2_X1 U714 ( .A(n636), .B(n635), .ZN(n637) );
  INV_X1 U715 ( .A(KEYINPUT56), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n718), .A2(G210), .ZN(n642) );
  XOR2_X1 U717 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n639) );
  XNOR2_X1 U718 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n642), .B(n641), .ZN(n643) );
  XOR2_X1 U720 ( .A(n646), .B(G101), .Z(G3) );
  NAND2_X1 U721 ( .A1(n648), .A2(n659), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n647), .B(G104), .ZN(G6) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n650) );
  NAND2_X1 U724 ( .A1(n648), .A2(n661), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U726 ( .A(G107), .B(n651), .ZN(G9) );
  XOR2_X1 U727 ( .A(n652), .B(G110), .Z(G12) );
  XOR2_X1 U728 ( .A(n653), .B(KEYINPUT29), .Z(n655) );
  NAND2_X1 U729 ( .A1(n657), .A2(n661), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n655), .B(n654), .ZN(G30) );
  XNOR2_X1 U731 ( .A(n656), .B(G143), .ZN(G45) );
  NAND2_X1 U732 ( .A1(n657), .A2(n659), .ZN(n658) );
  XNOR2_X1 U733 ( .A(n658), .B(G146), .ZN(G48) );
  NAND2_X1 U734 ( .A1(n439), .A2(n659), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n660), .B(G113), .ZN(G15) );
  NAND2_X1 U736 ( .A1(n439), .A2(n661), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n663), .B(G116), .ZN(G18) );
  XOR2_X1 U738 ( .A(G125), .B(KEYINPUT37), .Z(n664) );
  XNOR2_X1 U739 ( .A(n665), .B(n664), .ZN(G27) );
  XNOR2_X1 U740 ( .A(G134), .B(n666), .ZN(G36) );
  XOR2_X1 U741 ( .A(G140), .B(n667), .Z(G42) );
  NOR2_X1 U742 ( .A1(n696), .A2(n680), .ZN(n669) );
  NOR2_X1 U743 ( .A1(G953), .A2(n669), .ZN(n706) );
  XOR2_X1 U744 ( .A(KEYINPUT2), .B(n670), .Z(n704) );
  XNOR2_X1 U745 ( .A(KEYINPUT114), .B(KEYINPUT52), .ZN(n700) );
  NOR2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n677) );
  NOR2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U749 ( .A(KEYINPUT113), .B(n678), .Z(n679) );
  NOR2_X1 U750 ( .A1(n680), .A2(n679), .ZN(n698) );
  XOR2_X1 U751 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n694) );
  NAND2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U753 ( .A(n683), .B(KEYINPUT50), .ZN(n690) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U755 ( .A(KEYINPUT49), .B(n686), .Z(n687) );
  NOR2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U759 ( .A(n694), .B(n693), .Z(n695) );
  NOR2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U762 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U766 ( .A(n707), .B(KEYINPUT53), .ZN(n708) );
  XNOR2_X1 U767 ( .A(KEYINPUT115), .B(n708), .ZN(G75) );
  XOR2_X1 U768 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n711) );
  XNOR2_X1 U769 ( .A(n709), .B(KEYINPUT116), .ZN(n710) );
  XNOR2_X1 U770 ( .A(n711), .B(n710), .ZN(n713) );
  NAND2_X1 U771 ( .A1(n718), .A2(G469), .ZN(n712) );
  XNOR2_X1 U772 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U773 ( .A1(n724), .A2(n714), .ZN(G54) );
  NAND2_X1 U774 ( .A1(n718), .A2(G478), .ZN(n716) );
  NAND2_X1 U775 ( .A1(n718), .A2(G217), .ZN(n722) );
  INV_X1 U776 ( .A(KEYINPUT119), .ZN(n719) );
  NOR2_X1 U777 ( .A1(n724), .A2(n723), .ZN(G66) );
  XNOR2_X1 U778 ( .A(G101), .B(n725), .ZN(n726) );
  XNOR2_X1 U779 ( .A(n727), .B(n726), .ZN(n729) );
  NOR2_X1 U780 ( .A1(n729), .A2(n728), .ZN(n738) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U782 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U783 ( .A1(n731), .A2(G898), .ZN(n732) );
  XNOR2_X1 U784 ( .A(KEYINPUT120), .B(n732), .ZN(n736) );
  NAND2_X1 U785 ( .A1(n733), .A2(n745), .ZN(n734) );
  XOR2_X1 U786 ( .A(KEYINPUT121), .B(n734), .Z(n735) );
  NAND2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(G69) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U790 ( .A(n741), .B(KEYINPUT123), .ZN(n747) );
  INV_X1 U791 ( .A(n747), .ZN(n742) );
  XNOR2_X1 U792 ( .A(KEYINPUT124), .B(n742), .ZN(n744) );
  XNOR2_X1 U793 ( .A(n744), .B(n743), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(n745), .ZN(n751) );
  XNOR2_X1 U795 ( .A(G227), .B(n747), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n749), .A2(G953), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n751), .A2(n750), .ZN(G72) );
  XNOR2_X1 U799 ( .A(n752), .B(G131), .ZN(n753) );
  XNOR2_X1 U800 ( .A(n753), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U801 ( .A(G119), .B(KEYINPUT126), .Z(n754) );
  XNOR2_X1 U802 ( .A(n400), .B(n754), .ZN(G21) );
  XNOR2_X1 U803 ( .A(n756), .B(G122), .ZN(n757) );
  XNOR2_X1 U804 ( .A(n757), .B(KEYINPUT125), .ZN(G24) );
  XOR2_X1 U805 ( .A(n758), .B(G137), .Z(G39) );
endmodule

