//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n627, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157, new_n1158;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n459), .B1(new_n449), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(G137), .A3(new_n466), .ZN(new_n471));
  INV_X1    g046(.A(G113), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n464), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n473), .B1(new_n470), .B2(G125), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n469), .B(new_n471), .C1(new_n474), .C2(new_n466), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT70), .Z(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n466), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT72), .Z(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n486));
  NOR3_X1   g061(.A1(new_n481), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n470), .B2(new_n466), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n484), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n495), .A2(new_n478), .A3(new_n480), .A4(G138), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n478), .A2(new_n480), .A3(G138), .A4(new_n466), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT73), .B(KEYINPUT4), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n478), .A2(new_n480), .A3(G126), .ZN(new_n502));
  NAND2_X1  g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n466), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n498), .A2(new_n501), .A3(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(KEYINPUT74), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT74), .A3(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n515), .A2(new_n519), .ZN(G166));
  AND3_X1   g095(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT75), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT75), .B1(new_n507), .B2(new_n509), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n525), .B(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(KEYINPUT76), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n531), .B1(new_n512), .B2(new_n513), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n530), .A2(new_n532), .A3(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n507), .A2(new_n509), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n514), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n524), .A2(new_n527), .A3(new_n534), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  INV_X1    g114(.A(new_n521), .ZN(new_n540));
  INV_X1    g115(.A(new_n522), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(G64), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n516), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT78), .B(G52), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n530), .A2(new_n532), .A3(G543), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n528), .A2(new_n529), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n510), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n544), .A2(new_n550), .ZN(G171));
  INV_X1    g126(.A(KEYINPUT80), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n530), .A2(new_n532), .A3(G43), .A4(G543), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n523), .A2(G56), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n516), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n552), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n555), .B(KEYINPUT79), .ZN(new_n562));
  INV_X1    g137(.A(new_n560), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n562), .A2(KEYINPUT80), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  NAND4_X1  g146(.A1(new_n530), .A2(new_n532), .A3(G53), .A4(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(G78), .ZN(new_n574));
  INV_X1    g149(.A(G543), .ZN(new_n575));
  OR3_X1    g150(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT81), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT81), .B1(new_n574), .B2(new_n575), .ZN(new_n577));
  XNOR2_X1  g152(.A(KEYINPUT82), .B(G65), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n535), .C2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n536), .B2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT83), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n573), .A2(KEYINPUT83), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G171), .ZN(G301));
  INV_X1    g161(.A(G166), .ZN(G303));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(new_n521), .B2(new_n522), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n530), .A2(new_n532), .A3(G49), .A4(G543), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n547), .A2(G87), .A3(new_n507), .A4(new_n509), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(G288));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n535), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G651), .ZN(new_n598));
  NAND2_X1  g173(.A1(G48), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G86), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n535), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(new_n547), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n516), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n533), .A2(G47), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT84), .B(G85), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n548), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G290));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n548), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n536), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(new_n516), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n533), .A2(G54), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(G171), .ZN(G321));
  XOR2_X1   g197(.A(G321), .B(KEYINPUT85), .Z(G284));
  NAND2_X1  g198(.A1(G299), .A2(new_n620), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n620), .B2(G168), .ZN(G297));
  XOR2_X1   g200(.A(G297), .B(KEYINPUT86), .Z(G280));
  INV_X1    g201(.A(new_n619), .ZN(new_n627));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G860), .ZN(G148));
  NOR2_X1   g204(.A1(new_n619), .A2(G559), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n565), .B2(G868), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n490), .A2(G135), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(G111), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n464), .B1(new_n637), .B2(G2105), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n482), .A2(G123), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT88), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n468), .A2(new_n470), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT87), .B(G2100), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT15), .B(G2435), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(G14), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT17), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n672), .B(new_n673), .C1(new_n671), .C2(new_n667), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n673), .B2(new_n672), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT90), .B(G2096), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT91), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n686), .B1(new_n689), .B2(KEYINPUT20), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n683), .A2(new_n685), .A3(new_n687), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n690), .B(new_n691), .C1(KEYINPUT20), .C2(new_n689), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1991), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT92), .B(G1986), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n692), .B(new_n698), .ZN(G229));
  XNOR2_X1  g274(.A(KEYINPUT31), .B(G11), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G19), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n565), .B2(new_n701), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT95), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1341), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n490), .A2(G139), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT96), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT97), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G2105), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT25), .Z(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G29), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G29), .B2(G33), .ZN(new_n716));
  INV_X1    g291(.A(G2072), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G27), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G164), .B2(new_n719), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G2078), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n490), .A2(G141), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT26), .Z(new_n725));
  AOI22_X1  g300(.A1(new_n482), .A2(G129), .B1(G105), .B2(new_n468), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G32), .B(new_n727), .S(G29), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT27), .B(G1996), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n490), .A2(G140), .ZN(new_n731));
  OR2_X1    g306(.A1(G104), .A2(G2105), .ZN(new_n732));
  INV_X1    g307(.A(G116), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n464), .B1(new_n733), .B2(G2105), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n482), .A2(G128), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n719), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n719), .A2(G26), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT28), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(KEYINPUT28), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g314(.A1(G5), .A2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G171), .B2(G16), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n739), .A2(G2067), .B1(G1961), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n718), .A2(new_n722), .A3(new_n730), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n716), .A2(new_n717), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n627), .A2(new_n701), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G4), .B2(new_n701), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n741), .A2(G1961), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n746), .A2(new_n747), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n744), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n739), .A2(G2067), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n701), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n701), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT98), .B(G1966), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n743), .A2(new_n751), .A3(new_n752), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT99), .B(KEYINPUT23), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n701), .A2(G20), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G299), .B2(G16), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1956), .ZN(new_n762));
  INV_X1    g337(.A(G28), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT30), .B2(new_n763), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n765), .B1(new_n640), .B2(new_n719), .C1(new_n721), .C2(G2078), .ZN(new_n766));
  OR2_X1    g341(.A1(KEYINPUT24), .A2(G34), .ZN(new_n767));
  NAND2_X1  g342(.A1(KEYINPUT24), .A2(G34), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n767), .A2(new_n719), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G160), .B2(new_n719), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n766), .B1(new_n770), .B2(G2084), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n719), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n719), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT29), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n771), .B1(G2084), .B2(new_n770), .C1(new_n774), .C2(G2090), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G2090), .B2(new_n774), .ZN(new_n776));
  AND4_X1   g351(.A1(new_n705), .A2(new_n757), .A3(new_n762), .A4(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(G95), .A2(G2105), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n464), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n780), .B1(new_n779), .B2(new_n778), .C1(G107), .C2(new_n466), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n482), .A2(G119), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n490), .A2(G131), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G25), .B(new_n785), .S(G29), .Z(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT35), .B(G1991), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n701), .A2(G24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n609), .B2(new_n701), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n788), .B1(G1986), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n701), .A2(G23), .ZN(new_n792));
  INV_X1    g367(.A(G288), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n701), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT33), .Z(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G1976), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(G1976), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n701), .A2(G6), .ZN(new_n798));
  INV_X1    g373(.A(G305), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n701), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT32), .B(G1981), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n701), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n701), .ZN(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n796), .A2(new_n797), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n791), .B1(G1986), .B2(new_n790), .C1(new_n807), .C2(KEYINPUT34), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT94), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT36), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n807), .A2(KEYINPUT34), .ZN(new_n811));
  AND3_X1   g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n810), .B1(new_n809), .B2(new_n811), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n700), .B(new_n777), .C1(new_n812), .C2(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  NAND2_X1  g390(.A1(new_n523), .A2(G67), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT100), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n816), .A2(KEYINPUT100), .A3(new_n817), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n820), .A2(G651), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n533), .A2(G55), .B1(G93), .B2(new_n536), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n561), .A2(new_n564), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n822), .B(new_n823), .C1(new_n560), .C2(new_n557), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n619), .A2(new_n628), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n829));
  XOR2_X1   g404(.A(new_n828), .B(new_n829), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n827), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT101), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n822), .A2(new_n823), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n836), .ZN(G145));
  NOR2_X1   g412(.A1(new_n713), .A2(new_n644), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n731), .A2(new_n735), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT73), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(KEYINPUT4), .A3(G138), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n497), .B1(new_n481), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(new_n466), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n502), .A2(new_n503), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G2105), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n499), .A2(new_n500), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n840), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n490), .A2(G142), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n482), .A2(G130), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n854), .B(new_n855), .C1(G118), .C2(new_n466), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n850), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n849), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n713), .A2(new_n644), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n849), .A2(new_n857), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n839), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n860), .ZN(new_n863));
  INV_X1    g438(.A(new_n861), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n863), .A2(new_n838), .B1(new_n864), .B2(new_n858), .ZN(new_n865));
  AOI21_X1  g440(.A(G160), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n640), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n862), .A2(new_n865), .A3(G160), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n640), .B1(new_n871), .B2(new_n866), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n785), .B(new_n727), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n492), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n870), .A2(new_n872), .A3(new_n875), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT103), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n877), .A2(new_n882), .A3(new_n878), .A4(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g460(.A1(new_n834), .A2(G868), .ZN(new_n886));
  XNOR2_X1  g461(.A(G166), .B(G288), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n799), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n609), .B(KEYINPUT104), .Z(new_n889));
  XOR2_X1   g464(.A(new_n888), .B(new_n889), .Z(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT105), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n896), .A2(KEYINPUT106), .ZN(new_n897));
  INV_X1    g472(.A(new_n584), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT83), .B1(new_n573), .B2(new_n580), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n619), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n583), .A2(new_n627), .A3(new_n584), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT41), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n902), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n827), .B(new_n631), .ZN(new_n908));
  MUX2_X1   g483(.A(new_n906), .B(new_n907), .S(new_n908), .Z(new_n909));
  NOR2_X1   g484(.A1(new_n897), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n896), .A2(KEYINPUT106), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n886), .B1(new_n912), .B2(G868), .ZN(G295));
  AOI21_X1  g488(.A(new_n886), .B1(new_n912), .B2(G868), .ZN(G331));
  OAI21_X1  g489(.A(KEYINPUT107), .B1(new_n544), .B2(new_n550), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n544), .A2(KEYINPUT107), .A3(new_n550), .ZN(new_n917));
  OAI21_X1  g492(.A(G168), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(G286), .A3(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n824), .B2(new_n826), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n557), .A2(new_n552), .A3(new_n560), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT80), .B1(new_n562), .B2(new_n563), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n834), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n925), .A2(new_n825), .A3(new_n920), .A4(new_n918), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n906), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n922), .A2(new_n926), .A3(new_n907), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G37), .B1(new_n930), .B2(new_n891), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n891), .B2(new_n930), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n905), .A2(KEYINPUT108), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n903), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n902), .A2(KEYINPUT108), .A3(KEYINPUT41), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n936), .A2(new_n937), .B1(new_n922), .B2(new_n926), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n929), .B1(new_n938), .B2(KEYINPUT109), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n937), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(KEYINPUT109), .A3(new_n927), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n890), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n943), .A2(new_n931), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n933), .B(KEYINPUT44), .C1(new_n934), .C2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n931), .A3(new_n934), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n943), .A2(new_n931), .A3(KEYINPUT110), .A4(new_n934), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n951), .A2(KEYINPUT111), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT111), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(G397));
  OR2_X1    g530(.A1(new_n785), .A2(new_n787), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT125), .Z(new_n957));
  INV_X1    g532(.A(G1996), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n727), .B(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G2067), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n840), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n957), .A2(new_n962), .B1(G2067), .B2(new_n840), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT112), .B(G1384), .Z(new_n964));
  NAND2_X1  g539(.A1(new_n848), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G40), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT113), .B1(new_n475), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n469), .A2(new_n471), .ZN(new_n970));
  INV_X1    g545(.A(G125), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n481), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(G2105), .B1(new_n972), .B2(new_n473), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n970), .A2(new_n973), .A3(new_n974), .A4(G40), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n969), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n967), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n963), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n961), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n979), .B2(new_n727), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT46), .ZN(new_n981));
  INV_X1    g556(.A(new_n977), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(new_n982), .B2(G1996), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n977), .A2(KEYINPUT46), .A3(new_n958), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n980), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT47), .Z(new_n986));
  NAND2_X1  g561(.A1(new_n785), .A2(new_n787), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n959), .A2(new_n961), .A3(new_n987), .A4(new_n956), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n977), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT126), .Z(new_n990));
  NOR2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n977), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n993));
  XNOR2_X1  g568(.A(new_n992), .B(new_n993), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n978), .B(new_n986), .C1(new_n990), .C2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n515), .B2(new_n519), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT55), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n848), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n848), .B2(new_n999), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n976), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT114), .B(G2090), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n848), .A2(new_n999), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n966), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n848), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n969), .A3(new_n975), .A4(new_n1006), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1002), .A2(new_n1003), .B1(new_n1007), .B2(new_n805), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n997), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n805), .ZN(new_n1011));
  INV_X1    g586(.A(new_n976), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n848), .A2(new_n998), .A3(new_n999), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1003), .ZN(new_n1015));
  AOI211_X1 g590(.A(new_n1009), .B(new_n997), .C1(new_n1011), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n498), .A2(new_n504), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1384), .B1(new_n1019), .B2(new_n847), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(new_n969), .A3(new_n975), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n590), .A2(new_n593), .A3(G1976), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT115), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n590), .A2(new_n593), .A3(new_n1024), .A4(G1976), .ZN(new_n1025));
  AND4_X1   g600(.A1(G8), .A2(new_n1021), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n793), .A2(G1976), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1026), .A2(KEYINPUT116), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1020), .A2(new_n969), .A3(new_n975), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n1009), .ZN(new_n1032));
  AND2_X1   g607(.A1(G305), .A2(G1981), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  OR3_X1    g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1030), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1021), .A2(new_n1023), .A3(G8), .A4(new_n1025), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1040), .A2(KEYINPUT52), .A3(new_n1028), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n1040), .B2(KEYINPUT52), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT118), .B(new_n997), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n848), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1047), .A2(KEYINPUT119), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(KEYINPUT119), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n976), .B1(new_n966), .B2(new_n1004), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1966), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1013), .A2(new_n969), .A3(new_n975), .A4(new_n1014), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2084), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(G168), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1018), .A2(new_n1045), .A3(new_n1046), .A4(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1044), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1038), .A4(new_n1030), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1030), .B(new_n1038), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT117), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1010), .A2(KEYINPUT63), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1055), .A2(new_n1016), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1062), .A2(new_n1064), .A3(new_n1016), .ZN(new_n1069));
  INV_X1    g644(.A(G1976), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1038), .A2(new_n1070), .A3(new_n793), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1032), .B1(new_n1071), .B2(new_n1034), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n1021), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT121), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1012), .A2(new_n958), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1021), .A2(new_n1078), .A3(new_n1074), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1080), .A2(KEYINPUT59), .A3(new_n565), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT59), .B1(new_n1080), .B2(new_n565), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1053), .A2(new_n747), .B1(new_n1031), .B2(new_n960), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1084), .A2(KEYINPUT60), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1053), .A2(new_n747), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1031), .A2(new_n960), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(KEYINPUT60), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(KEYINPUT122), .A3(new_n619), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1086), .A2(new_n1090), .A3(KEYINPUT60), .A4(new_n1087), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n627), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1084), .B2(KEYINPUT60), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1085), .B(new_n1089), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT61), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n581), .B(KEYINPUT57), .Z(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1051), .A2(new_n1006), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1956), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1053), .A2(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1096), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1095), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1096), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(KEYINPUT61), .A3(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1083), .A2(new_n1094), .A3(new_n1103), .A4(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1084), .A2(new_n619), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1107), .B1(new_n1102), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1052), .A2(G286), .A3(new_n1054), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n1113), .B2(new_n1009), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1005), .A2(new_n969), .A3(new_n975), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1116), .A2(G1966), .B1(G2084), .B2(new_n1053), .ZN(new_n1117));
  OAI21_X1  g692(.A(G8), .B1(new_n1117), .B2(G286), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1117), .B2(G286), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1114), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1010), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1063), .B1(KEYINPUT118), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1007), .B2(G2078), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1002), .A2(G1961), .ZN(new_n1126));
  XNOR2_X1  g701(.A(G171), .B(KEYINPUT54), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n475), .A2(new_n968), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1124), .A2(G2078), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n967), .A2(new_n1128), .A3(new_n1006), .A4(new_n1129), .ZN(new_n1130));
  AND4_X1   g705(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1116), .A2(new_n1129), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1127), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1121), .A2(new_n1018), .A3(new_n1123), .A4(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1068), .B(new_n1073), .C1(new_n1112), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT123), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1121), .B(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1123), .A2(new_n1018), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1140), .A2(G171), .A3(new_n1133), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1143), .A2(new_n1141), .A3(new_n1121), .A4(new_n1135), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n1073), .A4(new_n1068), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1138), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  AND2_X1   g723(.A1(G290), .A2(G1986), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n988), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n977), .B1(new_n1150), .B2(new_n991), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1148), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n995), .B1(new_n1152), .B2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g729(.A(new_n678), .B1(new_n661), .B2(new_n662), .ZN(new_n1156));
  AOI21_X1  g730(.A(new_n1156), .B1(new_n881), .B2(new_n883), .ZN(new_n1157));
  NOR2_X1   g731(.A1(G229), .A2(new_n461), .ZN(new_n1158));
  NAND3_X1  g732(.A1(new_n1157), .A2(new_n951), .A3(new_n1158), .ZN(G225));
  INV_X1    g733(.A(G225), .ZN(G308));
endmodule


