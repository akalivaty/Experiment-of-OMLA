

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U560 ( .A1(G2105), .A2(G2104), .ZN(n905) );
  AND2_X1 U561 ( .A1(n594), .A2(n593), .ZN(n527) );
  XNOR2_X1 U562 ( .A(KEYINPUT30), .B(KEYINPUT91), .ZN(n662) );
  XNOR2_X1 U563 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X1 U564 ( .A1(n716), .A2(n598), .ZN(n656) );
  NAND2_X1 U565 ( .A1(n684), .A2(G8), .ZN(n714) );
  NOR2_X1 U566 ( .A1(G543), .A2(G651), .ZN(n811) );
  NOR2_X1 U567 ( .A1(G651), .A2(n540), .ZN(n807) );
  XNOR2_X1 U568 ( .A(n772), .B(KEYINPUT102), .ZN(n773) );
  XNOR2_X1 U569 ( .A(n774), .B(n773), .ZN(G329) );
  INV_X1 U570 ( .A(G651), .ZN(n532) );
  NOR2_X1 U571 ( .A1(G543), .A2(n532), .ZN(n528) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n528), .Z(n529) );
  XNOR2_X1 U573 ( .A(KEYINPUT68), .B(n529), .ZN(n808) );
  NAND2_X1 U574 ( .A1(n808), .A2(G61), .ZN(n538) );
  NAND2_X1 U575 ( .A1(G86), .A2(n811), .ZN(n531) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n540) );
  NAND2_X1 U577 ( .A1(G48), .A2(n807), .ZN(n530) );
  NAND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n536) );
  OR2_X1 U579 ( .A1(n532), .A2(n540), .ZN(n533) );
  XNOR2_X1 U580 ( .A(KEYINPUT67), .B(n533), .ZN(n812) );
  NAND2_X1 U581 ( .A1(n812), .A2(G73), .ZN(n534) );
  XOR2_X1 U582 ( .A(KEYINPUT2), .B(n534), .Z(n535) );
  NOR2_X1 U583 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U584 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U585 ( .A(n539), .B(KEYINPUT78), .ZN(G305) );
  NAND2_X1 U586 ( .A1(G87), .A2(n540), .ZN(n542) );
  NAND2_X1 U587 ( .A1(G74), .A2(G651), .ZN(n541) );
  NAND2_X1 U588 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U589 ( .A1(n808), .A2(n543), .ZN(n545) );
  NAND2_X1 U590 ( .A1(n807), .A2(G49), .ZN(n544) );
  NAND2_X1 U591 ( .A1(n545), .A2(n544), .ZN(G288) );
  NAND2_X1 U592 ( .A1(G52), .A2(n807), .ZN(n547) );
  NAND2_X1 U593 ( .A1(G64), .A2(n808), .ZN(n546) );
  NAND2_X1 U594 ( .A1(n547), .A2(n546), .ZN(n552) );
  NAND2_X1 U595 ( .A1(G90), .A2(n811), .ZN(n549) );
  NAND2_X1 U596 ( .A1(G77), .A2(n812), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n550), .Z(n551) );
  NOR2_X1 U599 ( .A1(n552), .A2(n551), .ZN(G171) );
  INV_X1 U600 ( .A(G171), .ZN(G301) );
  NAND2_X1 U601 ( .A1(G51), .A2(n807), .ZN(n554) );
  NAND2_X1 U602 ( .A1(G63), .A2(n808), .ZN(n553) );
  NAND2_X1 U603 ( .A1(n554), .A2(n553), .ZN(n556) );
  XOR2_X1 U604 ( .A(KEYINPUT73), .B(KEYINPUT6), .Z(n555) );
  XNOR2_X1 U605 ( .A(n556), .B(n555), .ZN(n564) );
  XNOR2_X1 U606 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n562) );
  NAND2_X1 U607 ( .A1(n811), .A2(G89), .ZN(n557) );
  XNOR2_X1 U608 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U609 ( .A1(G76), .A2(n812), .ZN(n558) );
  NAND2_X1 U610 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U611 ( .A(n560), .B(KEYINPUT5), .ZN(n561) );
  XNOR2_X1 U612 ( .A(n562), .B(n561), .ZN(n563) );
  NOR2_X1 U613 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U614 ( .A(KEYINPUT7), .B(n565), .Z(G168) );
  XOR2_X1 U615 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U616 ( .A1(n812), .A2(G75), .ZN(n567) );
  NAND2_X1 U617 ( .A1(n811), .A2(G88), .ZN(n566) );
  NAND2_X1 U618 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U619 ( .A1(G50), .A2(n807), .ZN(n569) );
  NAND2_X1 U620 ( .A1(G62), .A2(n808), .ZN(n568) );
  NAND2_X1 U621 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U622 ( .A1(n571), .A2(n570), .ZN(G166) );
  INV_X1 U623 ( .A(G166), .ZN(G303) );
  NAND2_X1 U624 ( .A1(G85), .A2(n811), .ZN(n573) );
  NAND2_X1 U625 ( .A1(G72), .A2(n812), .ZN(n572) );
  NAND2_X1 U626 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U627 ( .A1(G47), .A2(n807), .ZN(n575) );
  NAND2_X1 U628 ( .A1(G60), .A2(n808), .ZN(n574) );
  NAND2_X1 U629 ( .A1(n575), .A2(n574), .ZN(n576) );
  OR2_X1 U630 ( .A1(n577), .A2(n576), .ZN(G290) );
  XNOR2_X1 U631 ( .A(G305), .B(G1981), .ZN(n993) );
  INV_X1 U632 ( .A(KEYINPUT33), .ZN(n695) );
  NOR2_X1 U633 ( .A1(G2105), .A2(G2104), .ZN(n578) );
  XOR2_X1 U634 ( .A(KEYINPUT17), .B(n578), .Z(n579) );
  XNOR2_X1 U635 ( .A(KEYINPUT66), .B(n579), .ZN(n719) );
  NAND2_X1 U636 ( .A1(n719), .A2(G137), .ZN(n777) );
  AND2_X1 U637 ( .A1(n777), .A2(G40), .ZN(n588) );
  XOR2_X1 U638 ( .A(KEYINPUT64), .B(KEYINPUT23), .Z(n582) );
  INV_X1 U639 ( .A(G2105), .ZN(n580) );
  AND2_X1 U640 ( .A1(n580), .A2(G2104), .ZN(n900) );
  NAND2_X1 U641 ( .A1(G101), .A2(n900), .ZN(n581) );
  XNOR2_X1 U642 ( .A(n582), .B(n581), .ZN(n585) );
  NAND2_X1 U643 ( .A1(G113), .A2(n905), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT65), .B(n583), .Z(n584) );
  NAND2_X1 U645 ( .A1(n585), .A2(n584), .ZN(n780) );
  INV_X1 U646 ( .A(n780), .ZN(n586) );
  INV_X1 U647 ( .A(G2104), .ZN(n591) );
  AND2_X1 U648 ( .A1(n591), .A2(G2105), .ZN(n904) );
  NAND2_X1 U649 ( .A1(G125), .A2(n904), .ZN(n778) );
  AND2_X1 U650 ( .A1(n586), .A2(n778), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(n716) );
  INV_X1 U652 ( .A(G1384), .ZN(n589) );
  AND2_X1 U653 ( .A1(G138), .A2(n589), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n719), .A2(n590), .ZN(n597) );
  AND2_X1 U655 ( .A1(n591), .A2(G126), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G2105), .A2(n592), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G114), .A2(n905), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n900), .A2(G102), .ZN(n595) );
  AND2_X1 U659 ( .A1(n527), .A2(n595), .ZN(n775) );
  OR2_X1 U660 ( .A1(G1384), .A2(n775), .ZN(n596) );
  NAND2_X1 U661 ( .A1(n597), .A2(n596), .ZN(n717) );
  INV_X1 U662 ( .A(n717), .ZN(n598) );
  INV_X1 U663 ( .A(n656), .ZN(n684) );
  INV_X1 U664 ( .A(n714), .ZN(n707) );
  NOR2_X1 U665 ( .A1(G1976), .A2(G288), .ZN(n694) );
  NAND2_X1 U666 ( .A1(n707), .A2(n694), .ZN(n599) );
  NOR2_X1 U667 ( .A1(n695), .A2(n599), .ZN(n600) );
  XOR2_X1 U668 ( .A(n600), .B(KEYINPUT96), .Z(n701) );
  NAND2_X1 U669 ( .A1(G53), .A2(n807), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G65), .A2(n808), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G91), .A2(n811), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G78), .A2(n812), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U675 ( .A1(n606), .A2(n605), .ZN(n1001) );
  NAND2_X1 U676 ( .A1(n656), .A2(G2072), .ZN(n607) );
  XNOR2_X1 U677 ( .A(n607), .B(KEYINPUT27), .ZN(n609) );
  AND2_X1 U678 ( .A1(G1956), .A2(n684), .ZN(n608) );
  NOR2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n611) );
  NOR2_X1 U680 ( .A1(n1001), .A2(n611), .ZN(n610) );
  XOR2_X1 U681 ( .A(n610), .B(KEYINPUT28), .Z(n649) );
  NAND2_X1 U682 ( .A1(n1001), .A2(n611), .ZN(n647) );
  INV_X1 U683 ( .A(G2067), .ZN(n969) );
  NOR2_X1 U684 ( .A1(n684), .A2(n969), .ZN(n613) );
  AND2_X1 U685 ( .A1(n684), .A2(G1348), .ZN(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n623) );
  NAND2_X1 U687 ( .A1(G79), .A2(n812), .ZN(n615) );
  NAND2_X1 U688 ( .A1(G54), .A2(n807), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U690 ( .A(KEYINPUT70), .B(n616), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G92), .A2(n811), .ZN(n617) );
  XNOR2_X1 U692 ( .A(KEYINPUT69), .B(n617), .ZN(n618) );
  NOR2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G66), .A2(n808), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U696 ( .A(KEYINPUT15), .B(n622), .ZN(n995) );
  OR2_X1 U697 ( .A1(n623), .A2(n995), .ZN(n645) );
  NAND2_X1 U698 ( .A1(n623), .A2(n995), .ZN(n643) );
  NAND2_X1 U699 ( .A1(n808), .A2(G56), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT14), .B(n624), .Z(n630) );
  NAND2_X1 U701 ( .A1(n811), .A2(G81), .ZN(n625) );
  XNOR2_X1 U702 ( .A(n625), .B(KEYINPUT12), .ZN(n627) );
  NAND2_X1 U703 ( .A1(G68), .A2(n812), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U705 ( .A(KEYINPUT13), .B(n628), .Z(n629) );
  NOR2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n807), .A2(G43), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n996) );
  AND2_X1 U709 ( .A1(n684), .A2(G1341), .ZN(n636) );
  AND2_X1 U710 ( .A1(n636), .A2(KEYINPUT26), .ZN(n633) );
  NOR2_X1 U711 ( .A1(KEYINPUT90), .A2(n633), .ZN(n634) );
  NOR2_X1 U712 ( .A1(n996), .A2(n634), .ZN(n641) );
  XOR2_X1 U713 ( .A(G1996), .B(KEYINPUT89), .Z(n977) );
  NAND2_X1 U714 ( .A1(n656), .A2(n977), .ZN(n635) );
  XNOR2_X1 U715 ( .A(KEYINPUT26), .B(n635), .ZN(n638) );
  INV_X1 U716 ( .A(n636), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U718 ( .A1(KEYINPUT90), .A2(n639), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n650), .B(KEYINPUT29), .ZN(n654) );
  NOR2_X1 U725 ( .A1(n656), .A2(G1961), .ZN(n652) );
  XOR2_X1 U726 ( .A(G2078), .B(KEYINPUT25), .Z(n971) );
  NOR2_X1 U727 ( .A1(n684), .A2(n971), .ZN(n651) );
  NOR2_X1 U728 ( .A1(n652), .A2(n651), .ZN(n666) );
  NOR2_X1 U729 ( .A1(G301), .A2(n666), .ZN(n653) );
  OR2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n671) );
  INV_X1 U731 ( .A(G8), .ZN(n659) );
  INV_X1 U732 ( .A(G2084), .ZN(n655) );
  AND2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U734 ( .A(n657), .B(KEYINPUT88), .ZN(n658) );
  OR2_X1 U735 ( .A1(n659), .A2(n658), .ZN(n661) );
  NOR2_X1 U736 ( .A1(G1966), .A2(n714), .ZN(n660) );
  NOR2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n663) );
  NOR2_X1 U738 ( .A1(G168), .A2(n664), .ZN(n665) );
  XOR2_X1 U739 ( .A(KEYINPUT92), .B(n665), .Z(n668) );
  NAND2_X1 U740 ( .A1(n666), .A2(G301), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U742 ( .A(KEYINPUT31), .B(n669), .ZN(n670) );
  AND2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n672), .B(KEYINPUT93), .ZN(n682) );
  AND2_X1 U745 ( .A1(G286), .A2(G8), .ZN(n673) );
  NAND2_X1 U746 ( .A1(n682), .A2(n673), .ZN(n680) );
  NOR2_X1 U747 ( .A1(G2090), .A2(n684), .ZN(n674) );
  XNOR2_X1 U748 ( .A(KEYINPUT95), .B(n674), .ZN(n677) );
  NOR2_X1 U749 ( .A1(G1971), .A2(n714), .ZN(n675) );
  NOR2_X1 U750 ( .A1(G166), .A2(n675), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n677), .A2(n676), .ZN(n678) );
  OR2_X1 U752 ( .A1(n659), .A2(n678), .ZN(n679) );
  AND2_X1 U753 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n681), .B(KEYINPUT32), .ZN(n692) );
  XNOR2_X1 U755 ( .A(KEYINPUT94), .B(n682), .ZN(n690) );
  NAND2_X1 U756 ( .A1(G1966), .A2(KEYINPUT88), .ZN(n683) );
  NAND2_X1 U757 ( .A1(n683), .A2(n684), .ZN(n687) );
  XOR2_X1 U758 ( .A(KEYINPUT88), .B(G2084), .Z(n685) );
  NAND2_X1 U759 ( .A1(n685), .A2(n656), .ZN(n686) );
  NAND2_X1 U760 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U761 ( .A1(n688), .A2(G8), .ZN(n689) );
  NAND2_X1 U762 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n705) );
  NOR2_X1 U764 ( .A1(G1971), .A2(G303), .ZN(n693) );
  NOR2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n1004) );
  AND2_X1 U766 ( .A1(n1004), .A2(n695), .ZN(n696) );
  NAND2_X1 U767 ( .A1(n705), .A2(n696), .ZN(n699) );
  AND2_X1 U768 ( .A1(G1976), .A2(G288), .ZN(n1006) );
  NOR2_X1 U769 ( .A1(n1006), .A2(n714), .ZN(n697) );
  OR2_X1 U770 ( .A1(KEYINPUT33), .A2(n697), .ZN(n698) );
  AND2_X1 U771 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U773 ( .A1(n993), .A2(n702), .ZN(n710) );
  NOR2_X1 U774 ( .A1(G2090), .A2(G303), .ZN(n703) );
  NAND2_X1 U775 ( .A1(G8), .A2(n703), .ZN(n704) );
  NAND2_X1 U776 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U777 ( .A(n706), .B(KEYINPUT97), .ZN(n708) );
  NOR2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U779 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U780 ( .A(n711), .B(KEYINPUT98), .ZN(n762) );
  NOR2_X1 U781 ( .A1(G305), .A2(G1981), .ZN(n712) );
  XOR2_X1 U782 ( .A(n712), .B(KEYINPUT24), .Z(n713) );
  NOR2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U784 ( .A(KEYINPUT87), .B(n715), .ZN(n760) );
  NOR2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U786 ( .A(KEYINPUT83), .B(n718), .Z(n764) );
  NAND2_X1 U787 ( .A1(G119), .A2(n904), .ZN(n722) );
  INV_X1 U788 ( .A(n719), .ZN(n720) );
  INV_X1 U789 ( .A(n720), .ZN(n901) );
  NAND2_X1 U790 ( .A1(G131), .A2(n901), .ZN(n721) );
  NAND2_X1 U791 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U792 ( .A1(G95), .A2(n900), .ZN(n724) );
  NAND2_X1 U793 ( .A1(G107), .A2(n905), .ZN(n723) );
  NAND2_X1 U794 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n890) );
  NAND2_X1 U796 ( .A1(G1991), .A2(n890), .ZN(n736) );
  NAND2_X1 U797 ( .A1(G129), .A2(n904), .ZN(n728) );
  NAND2_X1 U798 ( .A1(G141), .A2(n901), .ZN(n727) );
  NAND2_X1 U799 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U800 ( .A1(G105), .A2(n900), .ZN(n729) );
  XNOR2_X1 U801 ( .A(n729), .B(KEYINPUT85), .ZN(n730) );
  XNOR2_X1 U802 ( .A(n730), .B(KEYINPUT38), .ZN(n731) );
  NOR2_X1 U803 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U804 ( .A1(n905), .A2(G117), .ZN(n733) );
  NAND2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n891) );
  NAND2_X1 U806 ( .A1(G1996), .A2(n891), .ZN(n735) );
  NAND2_X1 U807 ( .A1(n736), .A2(n735), .ZN(n950) );
  NAND2_X1 U808 ( .A1(n950), .A2(n764), .ZN(n737) );
  XOR2_X1 U809 ( .A(KEYINPUT86), .B(n737), .Z(n763) );
  NOR2_X1 U810 ( .A1(G1986), .A2(G290), .ZN(n738) );
  NOR2_X1 U811 ( .A1(G1991), .A2(n890), .ZN(n947) );
  NOR2_X1 U812 ( .A1(n738), .A2(n947), .ZN(n739) );
  NOR2_X1 U813 ( .A1(n763), .A2(n739), .ZN(n741) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n891), .ZN(n740) );
  XOR2_X1 U815 ( .A(KEYINPUT99), .B(n740), .Z(n954) );
  NOR2_X1 U816 ( .A1(n741), .A2(n954), .ZN(n742) );
  XNOR2_X1 U817 ( .A(n742), .B(KEYINPUT39), .ZN(n743) );
  XNOR2_X1 U818 ( .A(n743), .B(KEYINPUT100), .ZN(n754) );
  NAND2_X1 U819 ( .A1(n900), .A2(G104), .ZN(n745) );
  NAND2_X1 U820 ( .A1(G140), .A2(n901), .ZN(n744) );
  NAND2_X1 U821 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U822 ( .A(KEYINPUT34), .B(n746), .ZN(n752) );
  NAND2_X1 U823 ( .A1(G128), .A2(n904), .ZN(n748) );
  NAND2_X1 U824 ( .A1(G116), .A2(n905), .ZN(n747) );
  NAND2_X1 U825 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U826 ( .A(KEYINPUT84), .B(n749), .Z(n750) );
  XNOR2_X1 U827 ( .A(KEYINPUT35), .B(n750), .ZN(n751) );
  NOR2_X1 U828 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U829 ( .A(KEYINPUT36), .B(n753), .ZN(n912) );
  XNOR2_X1 U830 ( .A(G2067), .B(KEYINPUT37), .ZN(n755) );
  OR2_X1 U831 ( .A1(n912), .A2(n755), .ZN(n961) );
  NAND2_X1 U832 ( .A1(n754), .A2(n961), .ZN(n756) );
  NAND2_X1 U833 ( .A1(n912), .A2(n755), .ZN(n960) );
  NAND2_X1 U834 ( .A1(n756), .A2(n960), .ZN(n757) );
  NAND2_X1 U835 ( .A1(n764), .A2(n757), .ZN(n758) );
  XNOR2_X1 U836 ( .A(n758), .B(KEYINPUT101), .ZN(n769) );
  INV_X1 U837 ( .A(n769), .ZN(n759) );
  AND2_X1 U838 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U839 ( .A1(n762), .A2(n761), .ZN(n771) );
  INV_X1 U840 ( .A(n763), .ZN(n767) );
  XOR2_X1 U841 ( .A(G1986), .B(G290), .Z(n1010) );
  NAND2_X1 U842 ( .A1(n961), .A2(n1010), .ZN(n765) );
  NAND2_X1 U843 ( .A1(n765), .A2(n764), .ZN(n766) );
  AND2_X1 U844 ( .A1(n767), .A2(n766), .ZN(n768) );
  OR2_X1 U845 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U846 ( .A1(n771), .A2(n770), .ZN(n774) );
  INV_X1 U847 ( .A(KEYINPUT40), .ZN(n772) );
  NAND2_X1 U848 ( .A1(n901), .A2(G138), .ZN(n776) );
  AND2_X1 U849 ( .A1(n776), .A2(n775), .ZN(G164) );
  INV_X1 U850 ( .A(G96), .ZN(G221) );
  AND2_X1 U851 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U852 ( .A(G132), .ZN(G219) );
  INV_X1 U853 ( .A(G82), .ZN(G220) );
  INV_X1 U854 ( .A(G57), .ZN(G237) );
  NAND2_X1 U855 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U856 ( .A1(n780), .A2(n779), .ZN(G160) );
  NAND2_X1 U857 ( .A1(G7), .A2(G661), .ZN(n781) );
  XNOR2_X1 U858 ( .A(n781), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U859 ( .A(G223), .ZN(n845) );
  NAND2_X1 U860 ( .A1(n845), .A2(G567), .ZN(n782) );
  XOR2_X1 U861 ( .A(KEYINPUT11), .B(n782), .Z(G234) );
  INV_X1 U862 ( .A(G860), .ZN(n806) );
  OR2_X1 U863 ( .A1(n996), .A2(n806), .ZN(G153) );
  NAND2_X1 U864 ( .A1(G868), .A2(G301), .ZN(n784) );
  BUF_X1 U865 ( .A(n995), .Z(n919) );
  OR2_X1 U866 ( .A1(n919), .A2(G868), .ZN(n783) );
  NAND2_X1 U867 ( .A1(n784), .A2(n783), .ZN(G284) );
  INV_X1 U868 ( .A(n1001), .ZN(G299) );
  XOR2_X1 U869 ( .A(KEYINPUT74), .B(G868), .Z(n785) );
  NOR2_X1 U870 ( .A1(G286), .A2(n785), .ZN(n787) );
  NOR2_X1 U871 ( .A1(G868), .A2(G299), .ZN(n786) );
  NOR2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U873 ( .A(KEYINPUT75), .B(n788), .Z(G297) );
  NAND2_X1 U874 ( .A1(n806), .A2(G559), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n789), .A2(n919), .ZN(n790) );
  XNOR2_X1 U876 ( .A(n790), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U877 ( .A1(G868), .A2(n996), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n919), .A2(G868), .ZN(n791) );
  NOR2_X1 U879 ( .A1(G559), .A2(n791), .ZN(n792) );
  NOR2_X1 U880 ( .A1(n793), .A2(n792), .ZN(G282) );
  NAND2_X1 U881 ( .A1(n904), .A2(G123), .ZN(n794) );
  XNOR2_X1 U882 ( .A(n794), .B(KEYINPUT18), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G99), .A2(n900), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n905), .A2(G111), .ZN(n798) );
  NAND2_X1 U886 ( .A1(G135), .A2(n901), .ZN(n797) );
  NAND2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n946) );
  XNOR2_X1 U889 ( .A(n946), .B(G2096), .ZN(n801) );
  XNOR2_X1 U890 ( .A(n801), .B(KEYINPUT76), .ZN(n803) );
  INV_X1 U891 ( .A(G2100), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n803), .A2(n802), .ZN(G156) );
  XNOR2_X1 U893 ( .A(n996), .B(KEYINPUT77), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n919), .A2(G559), .ZN(n804) );
  XNOR2_X1 U895 ( .A(n805), .B(n804), .ZN(n824) );
  NAND2_X1 U896 ( .A1(n806), .A2(n824), .ZN(n817) );
  NAND2_X1 U897 ( .A1(G55), .A2(n807), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G67), .A2(n808), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n816) );
  NAND2_X1 U900 ( .A1(G93), .A2(n811), .ZN(n814) );
  NAND2_X1 U901 ( .A1(G80), .A2(n812), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U903 ( .A1(n816), .A2(n815), .ZN(n827) );
  XOR2_X1 U904 ( .A(n817), .B(n827), .Z(G145) );
  XNOR2_X1 U905 ( .A(n1001), .B(n827), .ZN(n820) );
  XOR2_X1 U906 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n818) );
  XNOR2_X1 U907 ( .A(G288), .B(n818), .ZN(n819) );
  XNOR2_X1 U908 ( .A(n820), .B(n819), .ZN(n821) );
  XNOR2_X1 U909 ( .A(G290), .B(n821), .ZN(n823) );
  XNOR2_X1 U910 ( .A(G166), .B(G305), .ZN(n822) );
  XNOR2_X1 U911 ( .A(n823), .B(n822), .ZN(n916) );
  XOR2_X1 U912 ( .A(n916), .B(KEYINPUT80), .Z(n825) );
  XNOR2_X1 U913 ( .A(n825), .B(n824), .ZN(n826) );
  NAND2_X1 U914 ( .A1(n826), .A2(G868), .ZN(n829) );
  OR2_X1 U915 ( .A1(n827), .A2(G868), .ZN(n828) );
  NAND2_X1 U916 ( .A1(n829), .A2(n828), .ZN(G295) );
  NAND2_X1 U917 ( .A1(G2084), .A2(G2078), .ZN(n830) );
  XOR2_X1 U918 ( .A(KEYINPUT20), .B(n830), .Z(n831) );
  NAND2_X1 U919 ( .A1(G2090), .A2(n831), .ZN(n832) );
  XNOR2_X1 U920 ( .A(KEYINPUT21), .B(n832), .ZN(n833) );
  NAND2_X1 U921 ( .A1(n833), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U922 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U923 ( .A1(G69), .A2(G120), .ZN(n834) );
  NOR2_X1 U924 ( .A1(G237), .A2(n834), .ZN(n835) );
  NAND2_X1 U925 ( .A1(G108), .A2(n835), .ZN(n849) );
  NAND2_X1 U926 ( .A1(G567), .A2(n849), .ZN(n836) );
  XOR2_X1 U927 ( .A(KEYINPUT82), .B(n836), .Z(n842) );
  NOR2_X1 U928 ( .A1(G220), .A2(G219), .ZN(n837) );
  XOR2_X1 U929 ( .A(KEYINPUT22), .B(n837), .Z(n838) );
  NOR2_X1 U930 ( .A1(G218), .A2(n838), .ZN(n839) );
  XNOR2_X1 U931 ( .A(n839), .B(KEYINPUT81), .ZN(n840) );
  OR2_X1 U932 ( .A1(G221), .A2(n840), .ZN(n850) );
  AND2_X1 U933 ( .A1(n850), .A2(G2106), .ZN(n841) );
  NOR2_X1 U934 ( .A1(n842), .A2(n841), .ZN(G319) );
  INV_X1 U935 ( .A(G319), .ZN(n844) );
  NAND2_X1 U936 ( .A1(G483), .A2(G661), .ZN(n843) );
  NOR2_X1 U937 ( .A1(n844), .A2(n843), .ZN(n848) );
  NAND2_X1 U938 ( .A1(n848), .A2(G36), .ZN(G176) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n845), .ZN(G217) );
  AND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U941 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U943 ( .A1(n848), .A2(n847), .ZN(G188) );
  INV_X1 U945 ( .A(G120), .ZN(G236) );
  INV_X1 U946 ( .A(G69), .ZN(G235) );
  NOR2_X1 U947 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U948 ( .A(KEYINPUT104), .B(n851), .ZN(G325) );
  INV_X1 U949 ( .A(G325), .ZN(G261) );
  XOR2_X1 U950 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n853) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(G2678), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U953 ( .A(KEYINPUT105), .B(G2072), .Z(n855) );
  XNOR2_X1 U954 ( .A(G2090), .B(G2067), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U956 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U957 ( .A(G2096), .B(G2100), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U959 ( .A(G2078), .B(n860), .ZN(n861) );
  XOR2_X1 U960 ( .A(n861), .B(G2084), .Z(G227) );
  XOR2_X1 U961 ( .A(G1976), .B(G1956), .Z(n863) );
  XNOR2_X1 U962 ( .A(G1966), .B(G1961), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U964 ( .A(G1986), .B(G1971), .Z(n865) );
  XNOR2_X1 U965 ( .A(G1991), .B(G1996), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U967 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U968 ( .A(KEYINPUT107), .B(G2474), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n871) );
  XOR2_X1 U970 ( .A(G1981), .B(KEYINPUT41), .Z(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U972 ( .A1(G124), .A2(n904), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n872), .B(KEYINPUT108), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G100), .A2(n900), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n905), .A2(G112), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G136), .A2(n901), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U980 ( .A1(n879), .A2(n878), .ZN(G162) );
  NAND2_X1 U981 ( .A1(G118), .A2(n905), .ZN(n888) );
  NAND2_X1 U982 ( .A1(n904), .A2(G130), .ZN(n880) );
  XNOR2_X1 U983 ( .A(KEYINPUT109), .B(n880), .ZN(n886) );
  NAND2_X1 U984 ( .A1(n900), .A2(G106), .ZN(n882) );
  NAND2_X1 U985 ( .A1(G142), .A2(n901), .ZN(n881) );
  NAND2_X1 U986 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U987 ( .A(KEYINPUT110), .B(n883), .Z(n884) );
  XNOR2_X1 U988 ( .A(KEYINPUT45), .B(n884), .ZN(n885) );
  NOR2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n889), .B(n946), .ZN(n894) );
  XNOR2_X1 U992 ( .A(G164), .B(n890), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(n894), .B(n893), .Z(n899) );
  XOR2_X1 U995 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n896) );
  XNOR2_X1 U996 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n895) );
  XNOR2_X1 U997 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U998 ( .A(G162), .B(n897), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n911) );
  NAND2_X1 U1000 ( .A1(n900), .A2(G103), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(G139), .A2(n901), .ZN(n902) );
  NAND2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n910) );
  NAND2_X1 U1003 ( .A1(G127), .A2(n904), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(G115), .A2(n905), .ZN(n906) );
  NAND2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1006 ( .A(KEYINPUT47), .B(n908), .Z(n909) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n940) );
  XOR2_X1 U1008 ( .A(n911), .B(n940), .Z(n914) );
  XOR2_X1 U1009 ( .A(G160), .B(n912), .Z(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n915), .ZN(G395) );
  XNOR2_X1 U1012 ( .A(n916), .B(KEYINPUT113), .ZN(n918) );
  XNOR2_X1 U1013 ( .A(n996), .B(G286), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n918), .B(n917), .ZN(n921) );
  XOR2_X1 U1015 ( .A(n919), .B(G301), .Z(n920) );
  XNOR2_X1 U1016 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n922), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(KEYINPUT114), .B(n923), .ZN(G397) );
  XOR2_X1 U1019 ( .A(G2454), .B(G2435), .Z(n925) );
  XNOR2_X1 U1020 ( .A(G2438), .B(G2427), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(n925), .B(n924), .ZN(n932) );
  XOR2_X1 U1022 ( .A(KEYINPUT103), .B(G2446), .Z(n927) );
  XNOR2_X1 U1023 ( .A(G2443), .B(G2430), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(n927), .B(n926), .ZN(n928) );
  XOR2_X1 U1025 ( .A(n928), .B(G2451), .Z(n930) );
  XNOR2_X1 U1026 ( .A(G1341), .B(G1348), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(n930), .B(n929), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n932), .B(n931), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n933), .A2(G14), .ZN(n939) );
  NAND2_X1 U1030 ( .A1(G319), .A2(n939), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(G227), .A2(G229), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(KEYINPUT49), .B(n934), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(G395), .A2(G397), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(G225) );
  INV_X1 U1036 ( .A(G225), .ZN(G308) );
  INV_X1 U1037 ( .A(G108), .ZN(G238) );
  INV_X1 U1038 ( .A(n939), .ZN(G401) );
  XNOR2_X1 U1039 ( .A(G2072), .B(n940), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(G164), .B(G2078), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(n941), .B(KEYINPUT116), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(n944), .B(KEYINPUT117), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT50), .B(n945), .ZN(n959) );
  XNOR2_X1 U1045 ( .A(G160), .B(G2084), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(KEYINPUT115), .B(n948), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n957) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(n955), .B(KEYINPUT51), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT52), .B(n964), .ZN(n965) );
  INV_X1 U1058 ( .A(KEYINPUT55), .ZN(n988) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n988), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n966), .A2(G29), .ZN(n1051) );
  XNOR2_X1 U1061 ( .A(G2090), .B(G35), .ZN(n983) );
  XNOR2_X1 U1062 ( .A(G1991), .B(G25), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G33), .B(G2072), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(G26), .B(n969), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n970), .A2(G28), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(G27), .B(n971), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(KEYINPUT118), .B(n972), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n980) );
  XOR2_X1 U1071 ( .A(G32), .B(n977), .Z(n978) );
  XNOR2_X1 U1072 ( .A(KEYINPUT119), .B(n978), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(KEYINPUT53), .B(n981), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(G34), .B(KEYINPUT54), .ZN(n984) );
  XOR2_X1 U1077 ( .A(n984), .B(G2084), .Z(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(n988), .B(n987), .ZN(n990) );
  INV_X1 U1080 ( .A(G29), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(G11), .A2(n991), .ZN(n1049) );
  XNOR2_X1 U1083 ( .A(G16), .B(KEYINPUT56), .ZN(n1018) );
  XOR2_X1 U1084 ( .A(G168), .B(G1966), .Z(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1086 ( .A(KEYINPUT57), .B(n994), .Z(n1016) );
  XNOR2_X1 U1087 ( .A(n995), .B(G1348), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(G301), .B(G1961), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n996), .B(G1341), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1014) );
  XNOR2_X1 U1092 ( .A(G1956), .B(n1001), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1002), .B(KEYINPUT120), .ZN(n1008) );
  NAND2_X1 U1094 ( .A1(G1971), .A2(G303), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT121), .B(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT122), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1047) );
  INV_X1 U1104 ( .A(G16), .ZN(n1045) );
  XNOR2_X1 U1105 ( .A(G1971), .B(G22), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(G24), .B(G1986), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XOR2_X1 U1108 ( .A(G1976), .B(G23), .Z(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n1023) );
  XNOR2_X1 U1111 ( .A(n1024), .B(n1023), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(G1966), .B(G21), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(G1961), .B(G5), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1041) );
  XNOR2_X1 U1116 ( .A(KEYINPUT59), .B(G1348), .ZN(n1029) );
  XNOR2_X1 U1117 ( .A(n1029), .B(G4), .ZN(n1037) );
  XOR2_X1 U1118 ( .A(G1981), .B(G6), .Z(n1030) );
  XNOR2_X1 U1119 ( .A(KEYINPUT123), .B(n1030), .ZN(n1032) );
  XNOR2_X1 U1120 ( .A(G19), .B(G1341), .ZN(n1031) );
  NOR2_X1 U1121 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1122 ( .A(KEYINPUT124), .B(n1033), .Z(n1035) );
  XNOR2_X1 U1123 ( .A(G1956), .B(G20), .ZN(n1034) );
  NOR2_X1 U1124 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1125 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XOR2_X1 U1126 ( .A(KEYINPUT125), .B(n1038), .Z(n1039) );
  XNOR2_X1 U1127 ( .A(KEYINPUT60), .B(n1039), .ZN(n1040) );
  NOR2_X1 U1128 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XOR2_X1 U1129 ( .A(n1042), .B(KEYINPUT61), .Z(n1043) );
  XNOR2_X1 U1130 ( .A(KEYINPUT127), .B(n1043), .ZN(n1044) );
  NAND2_X1 U1131 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NAND2_X1 U1132 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NOR2_X1 U1133 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  NAND2_X1 U1134 ( .A1(n1051), .A2(n1050), .ZN(n1052) );
  XOR2_X1 U1135 ( .A(KEYINPUT62), .B(n1052), .Z(G311) );
  INV_X1 U1136 ( .A(G311), .ZN(G150) );
endmodule

