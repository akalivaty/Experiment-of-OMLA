//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936;
  NAND2_X1  g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT7), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT8), .ZN(new_n204));
  AND2_X1   g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205));
  OAI221_X1 g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .C1(G85gat), .C2(G92gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G99gat), .B(G106gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT93), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT85), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT85), .ZN(new_n214));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215));
  AOI211_X1 g014(.A(new_n211), .B(new_n214), .C1(KEYINPUT15), .C2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n213), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT14), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n216), .B(new_n218), .C1(KEYINPUT15), .C2(new_n215), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n212), .B2(new_n213), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(KEYINPUT15), .A3(new_n215), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n209), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n219), .A2(new_n221), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT17), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n223), .B(new_n224), .C1(new_n209), .C2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G190gat), .B(G218gat), .Z(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT94), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT92), .ZN(new_n235));
  XOR2_X1   g034(.A(G134gat), .B(G162gat), .Z(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n230), .A2(new_n232), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n233), .A2(KEYINPUT95), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n237), .B(KEYINPUT95), .Z(new_n240));
  AND2_X1   g039(.A1(new_n230), .A2(new_n232), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n230), .A2(new_n232), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(G71gat), .A2(G78gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(G71gat), .A2(G78gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G57gat), .B(G64gat), .Z(new_n248));
  INV_X1    g047(.A(KEYINPUT90), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(KEYINPUT9), .B2(new_n245), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n251), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT21), .ZN(new_n255));
  XNOR2_X1  g054(.A(G127gat), .B(G155gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G231gat), .A2(G233gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT91), .ZN(new_n259));
  INV_X1    g058(.A(G183gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G211gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n257), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G15gat), .B(G22gat), .ZN(new_n265));
  INV_X1    g064(.A(G1gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(KEYINPUT16), .A3(new_n266), .ZN(new_n267));
  OAI221_X1 g066(.A(new_n267), .B1(KEYINPUT86), .B2(G8gat), .C1(new_n266), .C2(new_n265), .ZN(new_n268));
  NAND2_X1  g067(.A1(KEYINPUT86), .A2(G8gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  INV_X1    g069(.A(KEYINPUT21), .ZN(new_n271));
  INV_X1    g070(.A(new_n254), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n264), .A2(new_n275), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n244), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT10), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n209), .A2(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n208), .A2(new_n254), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n208), .A2(new_n254), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G230gat), .A2(G233gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n288), .B1(new_n284), .B2(new_n285), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G120gat), .B(G148gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G176gat), .B(G204gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n289), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n288), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n283), .B2(new_n286), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n294), .B1(new_n298), .B2(new_n290), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n280), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT89), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT36), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT32), .ZN(new_n305));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(KEYINPUT65), .A3(new_n308), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  AND2_X1   g116(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT28), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n320), .B2(new_n321), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n306), .B(new_n316), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT66), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT27), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n260), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n330));
  AOI21_X1  g129(.A(G190gat), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT28), .B1(new_n331), .B2(KEYINPUT64), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n334), .A2(KEYINPUT66), .A3(new_n306), .A4(new_n316), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G113gat), .B(G120gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(KEYINPUT1), .ZN(new_n338));
  XOR2_X1   g137(.A(G127gat), .B(G134gat), .Z(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT24), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(G183gat), .A3(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n306), .A2(KEYINPUT24), .ZN(new_n344));
  NOR2_X1   g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n308), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR3_X1   g147(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n341), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n343), .A2(new_n308), .ZN(new_n352));
  INV_X1    g151(.A(new_n345), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(KEYINPUT24), .A3(new_n306), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n313), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n347), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n352), .A2(new_n354), .A3(new_n357), .A4(KEYINPUT25), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n351), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n340), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n325), .A2(new_n326), .ZN(new_n364));
  INV_X1    g163(.A(new_n306), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n332), .B2(new_n333), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT66), .B1(new_n366), .B2(new_n316), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n360), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n340), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n359), .B1(new_n327), .B2(new_n335), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(KEYINPUT67), .A3(new_n340), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n363), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n305), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT33), .B1(new_n373), .B2(new_n375), .ZN(new_n377));
  XNOR2_X1  g176(.A(G15gat), .B(G43gat), .ZN(new_n378));
  INV_X1    g177(.A(G99gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT68), .B(G71gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n376), .A2(new_n377), .A3(new_n383), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n383), .A2(KEYINPUT69), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(KEYINPUT69), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(KEYINPUT33), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n376), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n363), .A2(new_n374), .A3(new_n370), .A4(new_n372), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT34), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n384), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT34), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n389), .B(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n375), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT32), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n397), .A3(new_n382), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n376), .A2(new_n387), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n393), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n304), .B1(new_n391), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n390), .B1(new_n384), .B2(new_n388), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(new_n399), .A3(new_n393), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(KEYINPUT36), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  INV_X1    g205(.A(G85gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT0), .B(G57gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(G155gat), .ZN(new_n413));
  INV_X1    g212(.A(G162gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT75), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT75), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n415), .A2(new_n419), .A3(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G141gat), .B(G148gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n414), .A2(KEYINPUT76), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(G162gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n425), .A3(G155gat), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n422), .B1(new_n426), .B2(KEYINPUT2), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n421), .A2(new_n427), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n422), .A2(KEYINPUT2), .ZN(new_n429));
  INV_X1    g228(.A(new_n417), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n369), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n421), .A2(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n340), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n412), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(KEYINPUT4), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT4), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n340), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT3), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n340), .B1(new_n440), .B2(new_n434), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n432), .A2(KEYINPUT3), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n437), .A2(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n436), .B1(new_n443), .B2(new_n412), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT5), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT5), .B1(new_n443), .B2(new_n412), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n411), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n443), .A2(new_n412), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n445), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n450), .B(new_n410), .C1(new_n445), .C2(new_n444), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n446), .A2(new_n447), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n454), .A2(KEYINPUT77), .A3(KEYINPUT6), .A4(new_n410), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT77), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n451), .B2(new_n452), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n453), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G211gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n462), .A3(G218gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT70), .B(KEYINPUT22), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G197gat), .B(G204gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(G211gat), .B(G218gat), .Z(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(new_n470), .A3(new_n466), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT72), .B1(new_n336), .B2(new_n360), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT72), .ZN(new_n476));
  AOI211_X1 g275(.A(new_n476), .B(new_n359), .C1(new_n327), .C2(new_n335), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT73), .ZN(new_n479));
  NAND2_X1  g278(.A1(G226gat), .A2(G233gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n480), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n368), .A2(new_n476), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n371), .A2(KEYINPUT72), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n482), .B1(new_n485), .B2(new_n474), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n360), .A2(new_n325), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT73), .B1(new_n488), .B2(new_n480), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n473), .B(new_n481), .C1(new_n486), .C2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n474), .A3(new_n480), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(new_n485), .B2(new_n480), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n472), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G64gat), .B(G92gat), .Z(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT74), .ZN(new_n496));
  XNOR2_X1  g295(.A(G8gat), .B(G36gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n496), .B(new_n497), .Z(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n490), .A2(new_n493), .A3(new_n498), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(KEYINPUT30), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n490), .A2(new_n503), .A3(new_n493), .A4(new_n498), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n459), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G78gat), .B(G106gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(G22gat), .B(G50gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT31), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G228gat), .ZN(new_n511));
  INV_X1    g310(.A(G233gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n434), .A2(new_n440), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n472), .B1(new_n514), .B2(new_n474), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n465), .A2(new_n470), .A3(new_n466), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n470), .B1(new_n465), .B2(new_n466), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT79), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n467), .A2(new_n518), .A3(new_n468), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n474), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT80), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n469), .A2(KEYINPUT79), .A3(new_n471), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT29), .B1(new_n517), .B2(new_n518), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT80), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n440), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n432), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n515), .B1(new_n528), .B2(KEYINPUT81), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n523), .A2(new_n524), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT3), .B1(new_n530), .B2(KEYINPUT80), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n434), .B1(new_n531), .B2(new_n526), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT81), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n513), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n440), .B1(new_n473), .B2(KEYINPUT29), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n432), .ZN(new_n537));
  INV_X1    g336(.A(new_n513), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n515), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT82), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n539), .A3(KEYINPUT82), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n535), .A2(KEYINPUT78), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT78), .ZN(new_n546));
  INV_X1    g345(.A(new_n515), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n532), .B2(new_n533), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n528), .A2(KEYINPUT81), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n538), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n544), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n510), .B1(new_n545), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT78), .B1(new_n535), .B2(new_n544), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(new_n551), .A3(new_n546), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n509), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n405), .B1(new_n505), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT83), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n554), .A2(new_n555), .A3(new_n509), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n509), .B1(new_n554), .B2(new_n555), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n501), .A2(new_n453), .A3(new_n455), .A4(new_n457), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT37), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n490), .A2(new_n564), .A3(new_n493), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n472), .B(new_n481), .C1(new_n486), .C2(new_n489), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n492), .B2(new_n473), .ZN(new_n567));
  AOI211_X1 g366(.A(KEYINPUT38), .B(new_n498), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n563), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n499), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n564), .B1(new_n490), .B2(new_n493), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT38), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n562), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n443), .A2(new_n412), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n410), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n433), .A2(new_n412), .A3(new_n435), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT39), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT40), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n581), .A2(new_n451), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n502), .A2(new_n583), .A3(new_n504), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n558), .A2(new_n559), .B1(new_n573), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n405), .B(KEYINPUT83), .C1(new_n505), .C2(new_n557), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n502), .A2(new_n504), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n458), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n391), .A2(new_n400), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n557), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT35), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n505), .A2(new_n592), .A3(new_n589), .A4(new_n557), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n585), .A2(new_n586), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n226), .A2(new_n270), .A3(new_n228), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n270), .A2(new_n225), .ZN(new_n596));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT18), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT87), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G113gat), .B(G141gat), .ZN(new_n601));
  INV_X1    g400(.A(G197gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT11), .B(G169gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n270), .B(new_n225), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n597), .B(KEYINPUT13), .Z(new_n609));
  AOI22_X1  g408(.A1(new_n598), .A2(new_n599), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT18), .A4(new_n597), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n610), .B(new_n611), .C1(new_n600), .C2(new_n606), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT88), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT88), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n303), .B1(new_n594), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n557), .B1(new_n587), .B2(new_n458), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n402), .A2(KEYINPUT36), .A3(new_n403), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT36), .B1(new_n402), .B2(new_n403), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n559), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n569), .A2(new_n572), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n557), .A3(new_n584), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n586), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n591), .A2(new_n593), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n632), .A2(KEYINPUT89), .A3(new_n620), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n302), .B1(new_n622), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n459), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G1gat), .ZN(G1324gat));
  INV_X1    g435(.A(KEYINPUT42), .ZN(new_n637));
  INV_X1    g436(.A(new_n587), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n244), .A2(new_n279), .A3(new_n300), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT89), .B1(new_n632), .B2(new_n620), .ZN(new_n640));
  AOI211_X1 g439(.A(new_n303), .B(new_n621), .C1(new_n630), .C2(new_n631), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT16), .B(G8gat), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n637), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT96), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(KEYINPUT96), .B(new_n637), .C1(new_n642), .C2(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n634), .A2(KEYINPUT42), .A3(new_n638), .A4(new_n643), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI211_X1 g451(.A(new_n587), .B(new_n302), .C1(new_n622), .C2(new_n633), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n653), .A2(KEYINPUT97), .A3(KEYINPUT42), .A4(new_n643), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n642), .A2(G8gat), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n649), .A2(new_n655), .A3(new_n656), .ZN(G1325gat));
  AOI21_X1  g456(.A(G15gat), .B1(new_n634), .B2(new_n589), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n626), .A2(G15gat), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n634), .B2(new_n659), .ZN(G1326gat));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n634), .A2(new_n661), .A3(new_n562), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n562), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT98), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT43), .B(G22gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  NAND2_X1  g466(.A1(new_n622), .A2(new_n633), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n279), .A2(new_n301), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n239), .A2(new_n243), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n668), .A2(new_n212), .A3(new_n459), .A4(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n672), .A2(KEYINPUT45), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(KEYINPUT45), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n623), .A2(new_n626), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n629), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n670), .B1(new_n676), .B2(new_n631), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(KEYINPUT44), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n632), .A2(KEYINPUT44), .A3(new_n244), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n669), .A2(new_n615), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n680), .A2(new_n459), .A3(new_n681), .ZN(new_n682));
  OAI22_X1  g481(.A1(new_n673), .A2(new_n674), .B1(new_n212), .B2(new_n682), .ZN(G1328gat));
  NAND3_X1  g482(.A1(new_n680), .A2(new_n638), .A3(new_n681), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n587), .A2(G36gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n668), .A2(new_n671), .A3(new_n685), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n684), .A2(G36gat), .B1(new_n686), .B2(KEYINPUT46), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(KEYINPUT46), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(KEYINPUT99), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n686), .A2(new_n690), .A3(KEYINPUT46), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n687), .B1(new_n689), .B2(new_n691), .ZN(G1329gat));
  NOR2_X1   g491(.A1(KEYINPUT100), .A2(KEYINPUT47), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n678), .A2(new_n626), .A3(new_n679), .A4(new_n681), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(G43gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(KEYINPUT100), .A2(KEYINPUT47), .ZN(new_n696));
  INV_X1    g495(.A(G43gat), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n668), .A2(new_n697), .A3(new_n589), .A4(new_n671), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n696), .B1(new_n695), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(G1330gat));
  NAND4_X1  g500(.A1(new_n678), .A2(new_n562), .A3(new_n679), .A4(new_n681), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G50gat), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n557), .A2(G50gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n668), .A2(new_n671), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1331gat));
  NAND3_X1  g507(.A1(new_n280), .A2(new_n615), .A3(new_n300), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT101), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n631), .B2(new_n676), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n459), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT103), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT102), .B(G57gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1332gat));
  AOI21_X1  g514(.A(new_n587), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT104), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1333gat));
  AOI21_X1  g519(.A(G71gat), .B1(new_n711), .B2(new_n589), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n626), .A2(G71gat), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n711), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g523(.A1(new_n711), .A2(new_n562), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT105), .B(G78gat), .Z(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1335gat));
  NOR3_X1   g526(.A1(new_n617), .A2(new_n301), .A3(new_n278), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n678), .A2(new_n679), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G85gat), .B1(new_n730), .B2(new_n458), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n617), .A2(new_n278), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n677), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT51), .B1(new_n677), .B2(new_n732), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n459), .A2(new_n407), .A3(new_n300), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n731), .B1(new_n737), .B2(new_n738), .ZN(G1336gat));
  NAND2_X1  g538(.A1(new_n729), .A2(new_n638), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n734), .A2(KEYINPUT106), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n677), .A2(new_n732), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n677), .B2(new_n732), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n587), .A2(G92gat), .A3(new_n301), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n740), .A2(G92gat), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n740), .A2(G92gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n745), .B1(new_n735), .B2(new_n736), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n747), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n750), .ZN(G1337gat));
  OAI21_X1  g550(.A(G99gat), .B1(new_n730), .B2(new_n405), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n589), .A2(new_n379), .A3(new_n300), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n737), .B2(new_n753), .ZN(G1338gat));
  NAND4_X1  g553(.A1(new_n678), .A2(new_n562), .A3(new_n679), .A4(new_n728), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G106gat), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n557), .A2(G106gat), .A3(new_n301), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n756), .B(new_n757), .C1(new_n737), .C2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n742), .B2(new_n743), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT107), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n763), .B(new_n758), .C1(new_n742), .C2(new_n743), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n762), .A2(new_n756), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n765), .B2(new_n757), .ZN(G1339gat));
  NAND2_X1  g565(.A1(new_n639), .A2(new_n615), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n610), .A2(new_n606), .A3(new_n611), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n608), .A2(new_n609), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n597), .B1(new_n595), .B2(new_n596), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n605), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n300), .A2(KEYINPUT109), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(new_n772), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n301), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n283), .A2(new_n297), .A3(new_n286), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n778), .A2(new_n298), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n294), .B1(new_n289), .B2(KEYINPUT54), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n295), .B1(new_n298), .B2(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n289), .A2(KEYINPUT54), .ZN(new_n784));
  OAI211_X1 g583(.A(KEYINPUT55), .B(new_n783), .C1(new_n784), .C2(new_n778), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n782), .A2(new_n296), .A3(new_n785), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n773), .B(new_n776), .C1(new_n786), .C2(new_n615), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n670), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n786), .A2(new_n670), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n775), .B(KEYINPUT108), .Z(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n768), .B1(new_n792), .B2(new_n279), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n793), .A2(new_n458), .A3(new_n590), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n587), .ZN(new_n795));
  OAI21_X1  g594(.A(G113gat), .B1(new_n795), .B2(new_n621), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n615), .A2(G113gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT110), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n795), .B2(new_n798), .ZN(G1340gat));
  NOR2_X1   g598(.A1(new_n795), .A2(new_n301), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT111), .B(G120gat), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1341gat));
  NOR2_X1   g601(.A1(new_n795), .A2(new_n279), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(G127gat), .Z(G1342gat));
  INV_X1    g603(.A(G134gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n587), .A2(new_n244), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT112), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n794), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n794), .A2(KEYINPUT113), .A3(new_n805), .A4(new_n808), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G134gat), .B1(new_n795), .B2(new_n670), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n811), .A2(new_n813), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(KEYINPUT56), .ZN(new_n818));
  AOI211_X1 g617(.A(KEYINPUT114), .B(new_n812), .C1(new_n811), .C2(new_n813), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n814), .B(new_n815), .C1(new_n818), .C2(new_n819), .ZN(G1343gat));
  NOR2_X1   g619(.A1(new_n793), .A2(new_n458), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n405), .A2(new_n562), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(KEYINPUT116), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(KEYINPUT116), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n821), .A2(new_n587), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n825), .A2(G141gat), .A3(new_n621), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n827), .B2(KEYINPUT58), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n626), .A2(new_n638), .A3(new_n458), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n562), .A2(KEYINPUT57), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n786), .B1(new_n616), .B2(new_n619), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n301), .A2(new_n775), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n670), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n278), .B1(new_n834), .B2(new_n791), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n831), .B1(new_n835), .B2(new_n768), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n787), .A2(new_n670), .B1(new_n789), .B2(new_n790), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n767), .B1(new_n837), .B2(new_n278), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT57), .B1(new_n838), .B2(new_n562), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI211_X1 g640(.A(KEYINPUT115), .B(KEYINPUT57), .C1(new_n838), .C2(new_n562), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n830), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n829), .B(G141gat), .C1(new_n843), .C2(new_n621), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n617), .B(new_n830), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n827), .A2(new_n826), .B1(new_n846), .B2(G141gat), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n829), .B2(new_n847), .ZN(G1344gat));
  OAI211_X1 g647(.A(new_n300), .B(new_n830), .C1(new_n841), .C2(new_n842), .ZN(new_n849));
  INV_X1    g648(.A(G148gat), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(KEYINPUT59), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT57), .B1(new_n793), .B2(new_n557), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n557), .A2(KEYINPUT57), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n302), .A2(new_n620), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n835), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n853), .A2(new_n300), .A3(new_n830), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G148gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT59), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n825), .A2(G148gat), .A3(new_n301), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(KEYINPUT118), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864));
  AOI22_X1  g663(.A1(new_n849), .A2(new_n851), .B1(new_n858), .B2(KEYINPUT59), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n861), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n866), .ZN(G1345gat));
  OR3_X1    g666(.A1(new_n843), .A2(new_n413), .A3(new_n279), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n413), .B1(new_n825), .B2(new_n279), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(G1346gat));
  NAND2_X1  g669(.A1(new_n423), .A2(new_n425), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n807), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n670), .A2(new_n871), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n843), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n875), .B(new_n876), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n590), .A2(new_n587), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n838), .A2(new_n458), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G169gat), .B1(new_n879), .B2(new_n621), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT120), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n615), .A2(G169gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n879), .B2(new_n882), .ZN(G1348gat));
  NOR2_X1   g682(.A1(new_n879), .A2(new_n301), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(G176gat), .Z(G1349gat));
  NOR2_X1   g684(.A1(new_n793), .A2(new_n459), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887));
  AOI211_X1 g686(.A(new_n319), .B(new_n318), .C1(new_n887), .C2(G183gat), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n886), .A2(new_n278), .A3(new_n878), .A4(new_n888), .ZN(new_n889));
  OAI22_X1  g688(.A1(new_n879), .A2(new_n279), .B1(new_n887), .B2(new_n260), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT122), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n889), .A2(new_n890), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n895), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(new_n892), .A3(new_n891), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT123), .B1(new_n896), .B2(new_n892), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(G1350gat));
  NOR2_X1   g700(.A1(new_n879), .A2(new_n670), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n317), .ZN(new_n904));
  XOR2_X1   g703(.A(KEYINPUT61), .B(G190gat), .Z(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n902), .B2(new_n905), .ZN(G1351gat));
  NAND3_X1  g705(.A1(new_n405), .A2(new_n638), .A3(new_n562), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT124), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(KEYINPUT124), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n886), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n602), .A3(new_n617), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n853), .A2(new_n856), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n626), .A2(new_n459), .A3(new_n587), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n915), .A2(new_n620), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n912), .B1(new_n916), .B2(new_n602), .ZN(G1352gat));
  XOR2_X1   g716(.A(KEYINPUT125), .B(G204gat), .Z(new_n918));
  OR3_X1    g717(.A1(new_n910), .A2(new_n301), .A3(new_n918), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n919), .A2(KEYINPUT62), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n913), .A2(new_n300), .A3(new_n914), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n918), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(KEYINPUT62), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(G1353gat));
  NAND2_X1  g723(.A1(new_n460), .A2(new_n462), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n911), .A2(new_n925), .A3(new_n278), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n853), .A2(new_n278), .A3(new_n856), .A4(new_n914), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n927), .B2(G211gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT126), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n932), .B(new_n926), .C1(new_n928), .C2(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1354gat));
  AOI21_X1  g733(.A(G218gat), .B1(new_n911), .B2(new_n244), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n244), .A2(G218gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n915), .B2(new_n936), .ZN(G1355gat));
endmodule


