//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n206), .B(new_n212), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT64), .Z(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(new_n215), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G87), .B(G97), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G107), .ZN(new_n236));
  INV_X1    g0036(.A(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  NAND2_X1  g0042(.A1(G33), .A2(G41), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n243), .A2(G1), .A3(G13), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT3), .B(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G222), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n246), .B1(new_n247), .B2(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  OR2_X1    g0049(.A1(KEYINPUT67), .A2(G223), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT67), .A2(G223), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n245), .B1(G77), .B2(new_n246), .C1(new_n248), .C2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  INV_X1    g0058(.A(new_n209), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(new_n243), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n257), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n245), .A2(new_n256), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n253), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G169), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n209), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n210), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G150), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n273), .A2(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G50), .A2(G58), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n210), .B1(new_n279), .B2(new_n216), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n272), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G50), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n283), .A2(new_n272), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT68), .ZN(new_n289));
  OAI21_X1  g0089(.A(G50), .B1(new_n210), .B2(G1), .ZN(new_n290));
  XOR2_X1   g0090(.A(new_n290), .B(KEYINPUT69), .Z(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n270), .A2(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n294), .A2(KEYINPUT70), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(KEYINPUT70), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n295), .B(new_n296), .C1(G179), .C2(new_n268), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT74), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT73), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT68), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n288), .B(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n291), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n299), .B1(new_n303), .B2(new_n286), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n287), .A2(new_n292), .A3(KEYINPUT73), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT9), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n298), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n304), .A2(KEYINPUT74), .A3(new_n305), .A4(KEYINPUT9), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n268), .A2(G200), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n268), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n306), .B2(new_n307), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n310), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n310), .B2(new_n315), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n297), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(G232), .A2(G1698), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n249), .A2(G238), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n246), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(G107), .B2(new_n246), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n244), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n323), .B2(new_n322), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n266), .A2(G244), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n325), .A2(new_n265), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(G169), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n273), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT15), .B(G87), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  OR3_X1    g0133(.A1(new_n332), .A2(new_n333), .A3(new_n274), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n332), .B2(new_n274), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n272), .ZN(new_n337));
  INV_X1    g0137(.A(G77), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n283), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n272), .B1(new_n261), .B2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G77), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n337), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n343), .B1(new_n327), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n327), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n342), .B1(new_n327), .B2(G190), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n329), .A2(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n276), .A2(G50), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT76), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n350), .B(new_n351), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n274), .A2(new_n338), .B1(new_n210), .B2(G68), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n272), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT11), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n355), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(KEYINPUT77), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n282), .A2(G68), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT12), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(G68), .B2(new_n340), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT77), .B1(new_n356), .B2(new_n357), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT3), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G33), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G232), .A2(G1698), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT75), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT75), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n246), .A2(new_n372), .A3(G232), .A4(G1698), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G97), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n365), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G226), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(G1698), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n246), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n244), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n244), .A2(G238), .A3(new_n262), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n265), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT13), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n382), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT13), .ZN(new_n385));
  INV_X1    g0185(.A(new_n378), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n369), .A2(new_n386), .B1(new_n365), .B2(new_n375), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n373), .B2(new_n371), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n384), .B(new_n385), .C1(new_n388), .C2(new_n244), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n383), .A2(G190), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n383), .A2(new_n389), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G200), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n364), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n383), .A2(new_n389), .A3(G179), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n269), .B1(new_n383), .B2(new_n389), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT14), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(new_n396), .A3(G169), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT78), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(KEYINPUT78), .A3(new_n396), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n349), .B(new_n393), .C1(new_n364), .C2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(KEYINPUT81), .A2(KEYINPUT17), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n273), .B1(new_n261), .B2(G20), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n301), .A2(new_n406), .B1(new_n282), .B2(new_n330), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(G20), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n365), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n368), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT79), .B1(new_n365), .B2(KEYINPUT3), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n409), .B1(new_n246), .B2(G20), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n216), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n214), .A2(new_n216), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G58), .A2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(G20), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n276), .A2(G159), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n408), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n272), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n369), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n415), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n421), .B1(new_n425), .B2(G68), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n423), .B1(new_n426), .B2(KEYINPUT16), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n407), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n377), .A2(G1698), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n246), .B(new_n429), .C1(G223), .C2(G1698), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n245), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n266), .A2(G232), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n433), .A2(new_n313), .A3(new_n265), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n265), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n244), .B1(new_n430), .B2(new_n431), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n346), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n404), .B1(new_n428), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT7), .B1(new_n369), .B2(new_n210), .ZN(new_n441));
  AOI211_X1 g0241(.A(new_n409), .B(G20), .C1(new_n366), .C2(new_n368), .ZN(new_n442));
  OAI21_X1  g0242(.A(G68), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n421), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(KEYINPUT16), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n422), .A2(new_n445), .A3(new_n272), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n289), .A2(new_n405), .B1(new_n283), .B2(new_n273), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT81), .B(KEYINPUT17), .ZN(new_n448));
  AND4_X1   g0248(.A1(new_n446), .A2(new_n439), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n440), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n447), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT80), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n446), .A2(KEYINPUT80), .A3(new_n447), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n433), .A2(G179), .A3(new_n265), .A4(new_n434), .ZN(new_n455));
  OAI21_X1  g0255(.A(G169), .B1(new_n436), .B2(new_n437), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT18), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n453), .A2(KEYINPUT18), .A3(new_n454), .A4(new_n457), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n450), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n366), .A2(new_n368), .A3(G244), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT4), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(G1698), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n467), .A2(new_n366), .A3(new_n368), .A4(G244), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n246), .A2(G250), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n249), .B1(new_n471), .B2(KEYINPUT4), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n245), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n261), .B(G45), .C1(new_n254), .C2(KEYINPUT5), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n260), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n255), .A2(G1), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n254), .A2(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n475), .A2(G41), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G257), .A3(new_n244), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n473), .A2(new_n344), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G250), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT4), .B1(new_n369), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G1698), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n468), .A2(new_n469), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n466), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n484), .B1(new_n491), .B2(new_n245), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n486), .B1(new_n492), .B2(G169), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n282), .A2(G97), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n261), .A2(G33), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n423), .A2(new_n282), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n496), .B2(G97), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(KEYINPUT6), .B2(G97), .ZN(new_n500));
  XNOR2_X1  g0300(.A(KEYINPUT82), .B(G107), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n500), .A2(new_n501), .ZN(new_n503));
  OAI21_X1  g0303(.A(G20), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n277), .A2(new_n338), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n414), .A2(new_n415), .ZN(new_n507));
  INV_X1    g0307(.A(G107), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n504), .B(new_n506), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n498), .B1(new_n509), .B2(new_n272), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT84), .B1(new_n493), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n500), .A2(new_n501), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n500), .A2(new_n501), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n210), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n508), .B1(new_n414), .B2(new_n415), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n514), .A2(new_n515), .A3(new_n505), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n497), .B1(new_n516), .B2(new_n423), .ZN(new_n517));
  AOI21_X1  g0317(.A(G169), .B1(new_n473), .B2(new_n485), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT84), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n486), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n511), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n366), .A2(new_n368), .A3(G250), .A4(new_n249), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G294), .ZN(new_n524));
  AND2_X1   g0324(.A1(G257), .A2(G1698), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n366), .A2(new_n368), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n244), .B1(new_n527), .B2(KEYINPUT92), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT92), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n523), .A2(new_n526), .A3(new_n529), .A4(new_n524), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n482), .A2(G264), .A3(new_n244), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n478), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n346), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(G190), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT25), .B1(new_n282), .B2(G107), .ZN(new_n536));
  OR3_X1    g0336(.A1(new_n282), .A2(KEYINPUT25), .A3(G107), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n288), .A2(new_n495), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(new_n508), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n539), .B(KEYINPUT91), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT23), .ZN(new_n543));
  AOI21_X1  g0343(.A(G20), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(KEYINPUT90), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(KEYINPUT23), .A2(G107), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n546), .B(new_n547), .C1(KEYINPUT90), .C2(new_n545), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n366), .A2(new_n368), .A3(new_n210), .A4(G87), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(KEYINPUT22), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT88), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n246), .A2(KEYINPUT88), .A3(new_n210), .A4(G87), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT22), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n550), .B1(new_n554), .B2(KEYINPUT89), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT89), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n552), .A2(new_n553), .A3(new_n556), .A4(KEYINPUT22), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n541), .B(new_n548), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n548), .B1(new_n555), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n272), .B1(new_n559), .B2(KEYINPUT24), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n535), .B(new_n540), .C1(new_n558), .C2(new_n560), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n332), .A2(new_n283), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n246), .A2(new_n210), .A3(G68), .ZN(new_n563));
  INV_X1    g0363(.A(G87), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n375), .A3(new_n508), .ZN(new_n565));
  OAI211_X1 g0365(.A(KEYINPUT19), .B(new_n565), .C1(new_n376), .C2(G20), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n274), .B2(new_n375), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n562), .B1(new_n569), .B2(new_n272), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n496), .A2(G87), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n217), .A2(G1698), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(new_n366), .A3(new_n368), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT85), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT85), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n246), .A2(new_n576), .A3(new_n573), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n366), .A2(new_n368), .A3(G244), .A4(G1698), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n542), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n244), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n479), .A2(new_n258), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n487), .B1(new_n255), .B2(G1), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n244), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(G200), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n580), .B1(new_n577), .B2(new_n575), .ZN(new_n588));
  OAI211_X1 g0388(.A(G190), .B(new_n585), .C1(new_n588), .C2(new_n244), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n572), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n473), .A2(new_n485), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G200), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT83), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n492), .B2(G190), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n593), .A2(new_n473), .A3(G190), .A4(new_n485), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n510), .B(new_n592), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n522), .A2(new_n561), .A3(new_n590), .A4(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n540), .B1(new_n560), .B2(new_n558), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT93), .ZN(new_n599));
  INV_X1    g0399(.A(new_n532), .ZN(new_n600));
  INV_X1    g0400(.A(new_n478), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n600), .B(new_n601), .C1(new_n528), .C2(new_n530), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n599), .B1(new_n602), .B2(new_n269), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n533), .A2(KEYINPUT93), .A3(G169), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(G179), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n269), .B1(new_n582), .B2(new_n586), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n570), .B1(new_n332), .B2(new_n538), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n344), .B(new_n585), .C1(new_n588), .C2(new_n244), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(G270), .B(new_n244), .C1(new_n474), .C2(new_n476), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT86), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT86), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n482), .A2(new_n614), .A3(G270), .A4(new_n244), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G303), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n244), .B1(new_n369), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n249), .A2(G257), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G264), .A2(G1698), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n246), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n618), .A2(new_n621), .B1(new_n260), .B2(new_n477), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n288), .A2(G116), .A3(new_n495), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n283), .A2(new_n237), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n271), .A2(new_n209), .B1(G20), .B2(new_n237), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n469), .B(new_n210), .C1(G33), .C2(new_n375), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n626), .A2(KEYINPUT20), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT20), .B1(new_n626), .B2(new_n627), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n624), .B(new_n625), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n623), .A2(G169), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT21), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(KEYINPUT87), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n616), .A2(G179), .A3(new_n622), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n630), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n632), .B1(new_n631), .B2(KEYINPUT87), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n623), .A2(new_n313), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n346), .B1(new_n616), .B2(new_n622), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n639), .A2(new_n630), .A3(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n637), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n607), .A2(new_n611), .A3(new_n642), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n597), .A2(new_n643), .ZN(new_n644));
  NOR4_X1   g0444(.A1(new_n318), .A2(new_n403), .A3(new_n463), .A4(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n297), .ZN(new_n646));
  INV_X1    g0446(.A(new_n450), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n329), .A2(new_n345), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n649), .A2(new_n393), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n402), .A2(new_n364), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n451), .A2(new_n457), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT18), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n316), .A2(new_n317), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n646), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n318), .A2(new_n403), .A3(new_n463), .ZN(new_n659));
  INV_X1    g0459(.A(new_n638), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n636), .A3(new_n633), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n598), .B2(new_n606), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n597), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g0463(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n664));
  NAND2_X1  g0464(.A1(new_n590), .A2(new_n611), .ZN(new_n665));
  AOI211_X1 g0465(.A(new_n664), .B(new_n665), .C1(new_n511), .C2(new_n521), .ZN(new_n666));
  INV_X1    g0466(.A(new_n665), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n493), .A2(new_n510), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT26), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n611), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n659), .B1(new_n663), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n658), .A2(new_n671), .ZN(G369));
  NOR2_X1   g0472(.A1(new_n637), .A2(new_n638), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n261), .A2(new_n210), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n540), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n554), .A2(KEYINPUT89), .ZN(new_n683));
  INV_X1    g0483(.A(new_n550), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(new_n557), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n548), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n423), .B1(new_n687), .B2(new_n541), .ZN(new_n688));
  INV_X1    g0488(.A(new_n558), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n682), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n679), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n561), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n607), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n607), .A2(new_n679), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT96), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT96), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n681), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n694), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n698), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n630), .A2(new_n679), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT95), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n642), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n673), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n700), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n204), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n565), .A2(G116), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n207), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n691), .B1(new_n663), .B2(new_n670), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT100), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AND4_X1   g0520(.A1(new_n590), .A2(new_n596), .A3(new_n511), .A4(new_n521), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n673), .B1(new_n690), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n723), .A3(new_n561), .ZN(new_n724));
  INV_X1    g0524(.A(new_n611), .ZN(new_n725));
  INV_X1    g0525(.A(new_n664), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n473), .A2(new_n344), .A3(new_n485), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n518), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n520), .B1(new_n728), .B2(new_n517), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n493), .A2(new_n510), .A3(KEYINPUT84), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n667), .B(new_n726), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT26), .ZN(new_n732));
  INV_X1    g0532(.A(new_n668), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n732), .B1(new_n733), .B2(new_n665), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n725), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n679), .B1(new_n724), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT100), .B1(new_n736), .B2(KEYINPUT29), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n511), .A2(new_n521), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n726), .B1(new_n738), .B2(new_n667), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n733), .A2(new_n665), .A3(new_n732), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n611), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT29), .B(new_n691), .C1(new_n663), .C2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n720), .A2(new_n737), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G330), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT31), .B1(new_n597), .B2(new_n643), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n582), .A2(new_n586), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n600), .B1(new_n528), .B2(new_n530), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n492), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n634), .A2(KEYINPUT97), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT97), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n616), .A2(new_n622), .A3(new_n750), .A4(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n748), .A2(KEYINPUT30), .A3(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n623), .B(new_n344), .C1(new_n582), .C2(new_n586), .ZN(new_n754));
  OAI21_X1  g0554(.A(KEYINPUT98), .B1(new_n602), .B2(new_n492), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT98), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n533), .A2(new_n591), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n754), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT31), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT99), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n492), .A2(new_n746), .A3(new_n747), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n751), .B2(new_n749), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n761), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n748), .A2(new_n752), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT30), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n765), .A2(KEYINPUT99), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n759), .A2(new_n760), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n679), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n745), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n759), .B1(KEYINPUT30), .B2(new_n763), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n691), .A2(new_n760), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n744), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n743), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n716), .B1(new_n777), .B2(G1), .ZN(G364));
  AND2_X1   g0578(.A1(new_n210), .A2(G13), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G45), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n712), .A2(G1), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n707), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G330), .B2(new_n705), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n781), .B(KEYINPUT101), .Z(new_n785));
  NAND2_X1  g0585(.A1(new_n246), .A2(new_n204), .ZN(new_n786));
  INV_X1    g0586(.A(G355), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n786), .A2(new_n787), .B1(G116), .B2(new_n204), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n710), .A2(new_n246), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n255), .B2(new_n208), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n241), .A2(G45), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(G20), .B1(KEYINPUT102), .B2(G169), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(KEYINPUT102), .A2(G169), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n209), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n785), .B1(new_n793), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n210), .A2(new_n313), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n344), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n246), .B1(new_n807), .B2(G322), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G179), .A2(G200), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n210), .B1(new_n809), .B2(G190), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G190), .ZN(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT33), .B(G317), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n811), .A2(G294), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n812), .A2(new_n313), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G326), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n808), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G283), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n210), .A2(G190), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n346), .A2(G179), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n805), .A2(new_n820), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n819), .A2(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n804), .A2(new_n821), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n820), .A2(new_n809), .ZN(new_n827));
  INV_X1    g0627(.A(G329), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n826), .A2(new_n617), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n818), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n831), .A2(KEYINPUT104), .ZN(new_n832));
  INV_X1    g0632(.A(new_n827), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G159), .ZN(new_n834));
  XOR2_X1   g0634(.A(KEYINPUT103), .B(KEYINPUT32), .Z(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n369), .B(new_n836), .C1(G58), .C2(new_n807), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n811), .A2(G97), .B1(G50), .B2(new_n816), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n834), .A2(new_n835), .B1(new_n813), .B2(G68), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n338), .A2(new_n823), .B1(new_n822), .B2(new_n508), .ZN(new_n840));
  INV_X1    g0640(.A(new_n826), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(G87), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n831), .A2(KEYINPUT104), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n832), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n803), .B1(new_n845), .B2(new_n797), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n800), .B(KEYINPUT105), .Z(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n705), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n784), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  NAND2_X1  g0650(.A1(new_n327), .A2(new_n344), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n342), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n852), .A2(new_n328), .A3(new_n679), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n347), .A2(new_n348), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n342), .A2(new_n679), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n853), .B1(new_n856), .B2(new_n648), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n717), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n691), .C1(new_n663), .C2(new_n670), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n782), .B1(new_n861), .B2(new_n775), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n775), .B2(new_n861), .ZN(new_n863));
  INV_X1    g0663(.A(new_n785), .ZN(new_n864));
  INV_X1    g0664(.A(new_n797), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n799), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT106), .Z(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n864), .B1(new_n338), .B2(new_n868), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n369), .B1(new_n810), .B2(new_n375), .C1(new_n508), .C2(new_n826), .ZN(new_n870));
  INV_X1    g0670(.A(new_n813), .ZN(new_n871));
  INV_X1    g0671(.A(new_n816), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n871), .A2(new_n819), .B1(new_n872), .B2(new_n617), .ZN(new_n873));
  INV_X1    g0673(.A(G294), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n806), .A2(new_n874), .B1(new_n823), .B2(new_n237), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n822), .A2(new_n564), .B1(new_n827), .B2(new_n824), .ZN(new_n876));
  NOR4_X1   g0676(.A1(new_n870), .A2(new_n873), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n823), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G143), .A2(new_n807), .B1(new_n878), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(G137), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n879), .B1(new_n872), .B2(new_n880), .C1(new_n275), .C2(new_n871), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT34), .ZN(new_n882));
  INV_X1    g0682(.A(new_n822), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(G68), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n284), .B2(new_n826), .ZN(new_n885));
  INV_X1    g0685(.A(G132), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n246), .B1(new_n827), .B2(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT107), .Z(new_n888));
  AOI211_X1 g0688(.A(new_n885), .B(new_n888), .C1(G58), .C2(new_n811), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n877), .B1(new_n882), .B2(new_n889), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n869), .B1(new_n865), .B2(new_n890), .C1(new_n857), .C2(new_n799), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n863), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(G384));
  NOR2_X1   g0693(.A1(new_n502), .A2(new_n503), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(G116), .A3(new_n211), .A4(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT36), .Z(new_n899));
  OAI211_X1 g0699(.A(new_n208), .B(G77), .C1(new_n214), .C2(new_n216), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n284), .A2(G68), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n261), .B(G13), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n677), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n453), .A2(new_n454), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT37), .B1(new_n428), .B2(new_n439), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n458), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n439), .A2(new_n446), .A3(new_n447), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n426), .A2(KEYINPUT16), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n407), .B1(new_n909), .B2(new_n427), .ZN(new_n910));
  INV_X1    g0710(.A(new_n457), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n910), .A2(new_n677), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT37), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n913), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n915), .B1(new_n462), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(KEYINPUT38), .B(new_n915), .C1(new_n462), .C2(new_n916), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(KEYINPUT108), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n853), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n860), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT108), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n917), .A2(new_n924), .A3(new_n918), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n679), .B1(new_n362), .B2(new_n363), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(new_n393), .C1(new_n402), .C2(new_n364), .ZN(new_n927));
  INV_X1    g0727(.A(new_n926), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n400), .A2(new_n401), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n929), .B2(new_n397), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n921), .A2(new_n923), .A3(new_n925), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n654), .A2(new_n677), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT109), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT109), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n932), .A2(new_n936), .A3(new_n933), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n921), .A2(KEYINPUT39), .A3(new_n925), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n905), .B1(new_n655), .B2(new_n647), .ZN(new_n939));
  INV_X1    g0739(.A(new_n907), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT37), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n653), .A2(new_n908), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n942), .B2(new_n905), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n918), .B1(new_n939), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(new_n920), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n938), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n651), .A2(new_n691), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT110), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n935), .A2(new_n937), .A3(new_n952), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n720), .A2(new_n737), .A3(new_n659), .A4(new_n742), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n954), .A2(new_n658), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n953), .B(new_n955), .Z(new_n956));
  INV_X1    g0756(.A(new_n772), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT99), .B1(new_n765), .B2(new_n766), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n761), .B(KEYINPUT30), .C1(new_n748), .C2(new_n752), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n957), .B1(new_n960), .B2(new_n759), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n745), .B2(new_n769), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n931), .A2(new_n857), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n921), .A3(new_n925), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT40), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n945), .B2(new_n920), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n965), .A2(new_n966), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n770), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n659), .B1(new_n970), .B2(new_n961), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n971), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(G330), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n956), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n261), .B2(new_n779), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n956), .A2(new_n974), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n903), .B1(new_n976), .B2(new_n977), .ZN(G367));
  OAI211_X1 g0778(.A(new_n522), .B(new_n596), .C1(new_n510), .C2(new_n691), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n668), .A2(new_n679), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n598), .A3(new_n606), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n679), .B1(new_n982), .B2(new_n522), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n699), .A2(new_n981), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n983), .B1(new_n984), .B2(KEYINPUT42), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT42), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n699), .A2(new_n986), .A3(new_n981), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n572), .A2(new_n691), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n665), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n725), .A2(new_n988), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n985), .A2(new_n987), .B1(KEYINPUT43), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(KEYINPUT43), .B2(new_n991), .ZN(new_n993));
  INV_X1    g0793(.A(new_n981), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n708), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT43), .ZN(new_n996));
  INV_X1    g0796(.A(new_n991), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n985), .A2(new_n996), .A3(new_n997), .A4(new_n987), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n993), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n995), .B1(new_n993), .B2(new_n998), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n711), .B(KEYINPUT41), .Z(new_n1002));
  INV_X1    g0802(.A(new_n708), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT45), .B1(new_n700), .B2(new_n981), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT45), .ZN(new_n1005));
  NOR4_X1   g0805(.A1(new_n699), .A2(new_n1005), .A3(new_n694), .A4(new_n994), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n981), .B1(KEYINPUT111), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n699), .B2(new_n694), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT112), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1009), .B(new_n1012), .C1(new_n699), .C2(new_n694), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1003), .B1(new_n1007), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n701), .A2(new_n680), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1018), .A2(new_n695), .A3(new_n981), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n1005), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1022), .A2(new_n708), .A3(new_n1015), .A4(new_n1014), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n697), .A2(new_n698), .A3(new_n681), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n706), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1018), .A2(new_n707), .A3(new_n1024), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(new_n776), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1017), .A2(new_n1023), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1002), .B1(new_n1030), .B2(new_n777), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n780), .A2(G1), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1001), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n991), .A2(new_n847), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n232), .A2(new_n789), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n801), .C1(new_n204), .C2(new_n332), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n822), .A2(new_n338), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n810), .A2(new_n216), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n369), .ZN(new_n1039));
  INV_X1    g0839(.A(G143), .ZN(new_n1040));
  INV_X1    g0840(.A(G159), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n872), .C1(new_n1041), .C2(new_n871), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n806), .A2(new_n275), .B1(new_n823), .B2(new_n284), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n826), .A2(new_n214), .B1(new_n827), .B2(new_n880), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT113), .Z(new_n1046));
  NAND2_X1  g0846(.A1(new_n833), .A2(G317), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n375), .B2(new_n822), .C1(new_n819), .C2(new_n823), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n826), .A2(new_n237), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(KEYINPUT46), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n508), .B2(new_n810), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1049), .A2(KEYINPUT46), .B1(new_n824), .B2(new_n872), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n369), .B1(new_n806), .B2(new_n617), .C1(new_n874), .C2(new_n871), .ZN(new_n1053));
  NOR4_X1   g0853(.A1(new_n1048), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1046), .A2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT47), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n785), .B(new_n1036), .C1(new_n1056), .C2(new_n865), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1034), .B1(new_n1057), .B2(KEYINPUT114), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(KEYINPUT114), .B2(new_n1057), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1033), .A2(new_n1059), .ZN(G387));
  INV_X1    g0860(.A(new_n1028), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n701), .A2(new_n847), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n786), .A2(new_n713), .B1(G107), .B2(new_n204), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n229), .A2(G45), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n273), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT50), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n330), .B2(new_n284), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n713), .B(new_n255), .C1(new_n216), .C2(new_n338), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1065), .B(new_n1067), .C1(KEYINPUT115), .C2(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(KEYINPUT115), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n790), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1063), .B1(new_n1064), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n785), .B1(new_n1072), .B2(new_n802), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n826), .A2(new_n874), .B1(new_n810), .B2(new_n819), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G317), .A2(new_n807), .B1(new_n878), .B2(G303), .ZN(new_n1075));
  INV_X1    g0875(.A(G322), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1075), .B1(new_n872), .B2(new_n1076), .C1(new_n824), .C2(new_n871), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT48), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT49), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n822), .A2(new_n237), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n246), .B(new_n1084), .C1(G326), .C2(new_n833), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n246), .B1(new_n822), .B2(new_n375), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n330), .B2(new_n813), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G77), .A2(new_n841), .B1(new_n833), .B2(G150), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G50), .A2(new_n807), .B1(new_n878), .B2(G68), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n810), .A2(new_n332), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n816), .B2(G159), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1086), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1073), .B1(new_n1094), .B2(new_n797), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1061), .A2(new_n1032), .B1(new_n1062), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1029), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n711), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1061), .A2(new_n777), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(G393));
  NAND3_X1  g0900(.A1(new_n1017), .A2(new_n1023), .A3(new_n1032), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n994), .A2(new_n800), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT116), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n238), .A2(new_n790), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n801), .B1(new_n375), .B2(new_n204), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n785), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n872), .A2(new_n275), .B1(new_n806), .B2(new_n1041), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT51), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n810), .A2(new_n338), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n246), .B1(new_n822), .B2(new_n564), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(G50), .C2(new_n813), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n823), .A2(new_n273), .B1(new_n827), .B2(new_n1040), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G68), .B2(new_n841), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1108), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT117), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n807), .A2(G311), .B1(G317), .B2(new_n816), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT52), .Z(new_n1118));
  OAI22_X1  g0918(.A1(new_n823), .A2(new_n874), .B1(new_n827), .B2(new_n1076), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G283), .B2(new_n841), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n369), .B1(new_n822), .B2(new_n508), .C1(new_n871), .C2(new_n617), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G116), .B2(new_n811), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1118), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1116), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1106), .B1(new_n1125), .B2(new_n797), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1103), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1101), .A2(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1030), .A2(new_n711), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1017), .A2(new_n1023), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1097), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1128), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(G390));
  AOI21_X1  g0933(.A(new_n853), .B1(new_n736), .B2(new_n857), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n931), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n950), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n938), .A2(new_n1136), .A3(new_n947), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n945), .A2(new_n920), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n741), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n679), .B1(new_n1139), .B2(new_n724), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n856), .A2(new_n648), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n853), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n950), .B(new_n1138), .C1(new_n1142), .C2(new_n1135), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n962), .A2(new_n963), .A3(new_n744), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n774), .A2(new_n857), .A3(new_n931), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1137), .A2(new_n1143), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n659), .B(G330), .C1(new_n970), .C2(new_n961), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n954), .A2(new_n1150), .A3(new_n658), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n931), .B1(new_n774), .B2(new_n857), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n923), .B1(new_n1152), .B2(new_n1145), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n962), .A2(new_n744), .A3(new_n858), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1147), .B(new_n1142), .C1(new_n931), .C2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1151), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1149), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1146), .A2(new_n1156), .A3(new_n1148), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n711), .A3(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1146), .A2(new_n1032), .A3(new_n1148), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT54), .B(G143), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n823), .A2(new_n1162), .B1(new_n827), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n841), .A2(G150), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT53), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(G50), .C2(new_n883), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n246), .B1(new_n806), .B2(new_n886), .ZN(new_n1168));
  INV_X1    g0968(.A(G128), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n871), .A2(new_n880), .B1(new_n872), .B2(new_n1169), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(G159), .C2(new_n811), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n369), .B1(new_n826), .B2(new_n564), .C1(new_n819), .C2(new_n872), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n884), .B1(new_n375), .B2(new_n823), .C1(new_n874), .C2(new_n827), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(G107), .C2(new_n813), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1109), .B1(G116), .B2(new_n807), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT118), .Z(new_n1176));
  AOI22_X1  g0976(.A1(new_n1167), .A2(new_n1171), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n785), .B1(new_n330), .B2(new_n867), .C1(new_n1177), .C2(new_n865), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT119), .Z(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n948), .B2(new_n799), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1161), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1160), .A2(new_n1181), .ZN(G378));
  NAND2_X1  g0982(.A1(new_n965), .A2(new_n966), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n967), .A2(new_n964), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n318), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1185), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n297), .B(new_n1187), .C1(new_n316), .C2(new_n317), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n306), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n677), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1186), .A2(new_n306), .A3(new_n904), .A4(new_n1188), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AND4_X1   g0993(.A1(G330), .A2(new_n1183), .A3(new_n1184), .A4(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n968), .B2(G330), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n953), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1183), .A2(G330), .A3(new_n1184), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1193), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n934), .A2(KEYINPUT109), .B1(new_n948), .B2(new_n951), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n968), .A2(G330), .A3(new_n1193), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1199), .A2(new_n937), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1151), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1196), .A2(new_n1202), .B1(new_n1159), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n711), .B1(new_n1204), .B2(KEYINPUT57), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1196), .A2(new_n1202), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1159), .A2(new_n1203), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1206), .A2(KEYINPUT57), .A3(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1198), .A2(new_n798), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n806), .A2(new_n508), .B1(new_n827), .B2(new_n819), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n332), .A2(new_n823), .B1(new_n822), .B2(new_n214), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G41), .B(new_n246), .C1(new_n841), .C2(G77), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1211), .B(new_n1212), .C1(new_n1213), .C2(KEYINPUT120), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n872), .A2(new_n237), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1038), .B(new_n1215), .C1(G97), .C2(new_n813), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(KEYINPUT120), .C2(new_n1213), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT58), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n254), .B1(new_n367), .B2(new_n365), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1217), .A2(new_n1218), .B1(new_n284), .B2(new_n1219), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n872), .A2(new_n1163), .B1(new_n810), .B2(new_n275), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n878), .A2(G137), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n1169), .B2(new_n806), .C1(new_n826), .C2(new_n1162), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(G132), .C2(new_n813), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n365), .B(new_n254), .C1(new_n822), .C2(new_n1041), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G124), .B2(new_n833), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT59), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1228), .B1(new_n1224), .B2(new_n1229), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1220), .B1(new_n1218), .B2(new_n1217), .C1(new_n1226), .C2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n797), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n782), .B1(new_n867), .B2(G50), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT121), .Z(new_n1234));
  NAND3_X1  g1034(.A1(new_n1210), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1206), .B2(new_n1032), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1209), .A2(new_n1237), .ZN(G375));
  NAND2_X1  g1038(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1135), .A2(new_n798), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n785), .B1(new_n867), .B2(G68), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n806), .A2(new_n880), .B1(new_n827), .B2(new_n1169), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n886), .A2(new_n872), .B1(new_n871), .B2(new_n1162), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(G159), .C2(new_n841), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n823), .A2(new_n275), .B1(new_n810), .B2(new_n284), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT123), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n246), .B1(new_n822), .B2(new_n214), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT124), .Z(new_n1248));
  NAND3_X1  g1048(.A1(new_n1244), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n872), .A2(new_n874), .B1(new_n823), .B2(new_n508), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G116), .B2(new_n813), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n1251), .B(KEYINPUT122), .Z(new_n1252));
  NOR3_X1   g1052(.A1(new_n1037), .A2(new_n1091), .A3(new_n246), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(G97), .A2(new_n841), .B1(new_n833), .B2(G303), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(new_n819), .C2(new_n806), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1249), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1241), .B1(new_n1256), .B2(new_n797), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1239), .A2(new_n1032), .B1(new_n1240), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1002), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1157), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1239), .A2(new_n1203), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(G381));
  INV_X1    g1062(.A(G375), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1033), .A2(new_n1132), .A3(new_n1059), .ZN(new_n1264));
  OR2_X1    g1064(.A1(G393), .A2(G396), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1265), .A2(G378), .A3(G384), .A4(G381), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .ZN(G407));
  INV_X1    g1067(.A(G378), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n678), .A2(G213), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1263), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(KEYINPUT125), .Z(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(G213), .A3(G407), .ZN(G409));
  XNOR2_X1  g1073(.A(G393), .B(new_n849), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1132), .B1(new_n1033), .B2(new_n1059), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1264), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G387), .A2(G390), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1033), .A2(new_n1132), .A3(new_n1059), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1274), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1196), .A2(new_n1202), .A3(KEYINPUT126), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT126), .B1(new_n1196), .B2(new_n1202), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1032), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1206), .A2(new_n1259), .A3(new_n1207), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1235), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1268), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1237), .C1(new_n1205), .C2(new_n1208), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1270), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n712), .B(new_n1156), .C1(new_n1261), .C2(KEYINPUT60), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(KEYINPUT60), .B2(new_n1261), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(G384), .A3(new_n1258), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G384), .B1(new_n1292), .B2(new_n1258), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT62), .B1(new_n1290), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1299), .B2(new_n1269), .ZN(new_n1300));
  AOI211_X1 g1100(.A(KEYINPUT127), .B(new_n1270), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1296), .A2(KEYINPUT62), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1297), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1270), .A2(G2897), .ZN(new_n1305));
  OR3_X1    g1105(.A1(new_n1294), .A2(new_n1295), .A3(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1305), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1281), .B1(new_n1304), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1302), .A2(KEYINPUT63), .A3(new_n1296), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1281), .A2(KEYINPUT61), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1290), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1296), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1308), .A2(new_n1316), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1313), .A2(new_n1314), .A3(new_n1318), .A4(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1312), .A2(new_n1320), .ZN(G405));
  NAND2_X1  g1121(.A1(G375), .A2(new_n1268), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1289), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1296), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1322), .A2(new_n1289), .A3(new_n1317), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1281), .ZN(G402));
endmodule


