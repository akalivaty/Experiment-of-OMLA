//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT69), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n454), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT70), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT72), .A3(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2104), .ZN(new_n479));
  AND4_X1   g054(.A1(new_n464), .A2(new_n474), .A3(new_n476), .A4(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT73), .B1(new_n480), .B2(G137), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n474), .A2(new_n476), .A3(new_n479), .A4(new_n464), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT73), .ZN(new_n483));
  INV_X1    g058(.A(G137), .ZN(new_n484));
  NOR3_X1   g059(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n472), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT74), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n474), .A2(new_n476), .A3(new_n479), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n488), .A2(KEYINPUT73), .A3(G137), .A4(new_n464), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n483), .B1(new_n482), .B2(new_n484), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT74), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(new_n472), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n468), .B1(new_n487), .B2(new_n493), .ZN(G160));
  NAND2_X1  g069(.A1(new_n488), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G124), .ZN(new_n496));
  NOR2_X1   g071(.A1(G100), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(new_n464), .B2(G112), .ZN(new_n498));
  OAI22_X1  g073(.A1(new_n495), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n480), .A2(KEYINPUT75), .A3(G136), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT75), .B1(new_n480), .B2(G136), .ZN(new_n501));
  OR3_X1    g076(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G162));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT4), .B1(new_n482), .B2(new_n504), .ZN(new_n505));
  NOR3_X1   g080(.A1(new_n504), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n465), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT76), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT76), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n465), .A2(new_n509), .A3(new_n506), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n505), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n474), .A2(new_n476), .A3(new_n479), .A4(G126), .ZN(new_n512));
  NAND2_X1  g087(.A1(G114), .A2(G2104), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n469), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n514), .A2(G2105), .B1(G102), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n511), .A2(new_n516), .A3(KEYINPUT77), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(G164));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT78), .B(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT6), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT6), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G50), .ZN(new_n528));
  INV_X1    g103(.A(new_n523), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G75), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n522), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n522), .A2(KEYINPUT5), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n522), .A2(KEYINPUT5), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n527), .A2(G88), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n529), .A2(G62), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n531), .A2(new_n537), .ZN(G166));
  XNOR2_X1  g113(.A(KEYINPUT80), .B(G89), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n527), .A2(new_n539), .B1(G63), .B2(G651), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n534), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n524), .A2(new_n526), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n522), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G51), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT79), .B(KEYINPUT7), .Z(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n545), .B(new_n546), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n541), .A2(new_n544), .A3(new_n547), .ZN(G168));
  INV_X1    g123(.A(new_n534), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n549), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n523), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n542), .A2(new_n534), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n543), .A2(G52), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n534), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n543), .A2(G43), .B1(new_n529), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n552), .A2(G81), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND3_X1  g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  XOR2_X1   g141(.A(KEYINPUT81), .B(KEYINPUT8), .Z(new_n567));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G188));
  AOI22_X1  g145(.A1(new_n549), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n525), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n524), .A2(KEYINPUT82), .A3(G543), .A4(new_n526), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OR3_X1    g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n552), .A2(G91), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n574), .B1(new_n573), .B2(new_n575), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n572), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(G299));
  NAND3_X1  g154(.A1(new_n541), .A2(new_n544), .A3(new_n547), .ZN(G286));
  INV_X1    g155(.A(G166), .ZN(G303));
  NAND2_X1  g156(.A1(new_n527), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G49), .ZN(new_n583));
  OR3_X1    g158(.A1(new_n582), .A2(KEYINPUT83), .A3(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n549), .A2(G74), .ZN(new_n585));
  AOI22_X1  g160(.A1(G87), .A2(new_n552), .B1(new_n585), .B2(G651), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT83), .B1(new_n582), .B2(new_n583), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n543), .A2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n552), .A2(G86), .ZN(new_n591));
  INV_X1    g166(.A(G73), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT84), .B1(new_n592), .B2(new_n522), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n592), .A2(new_n522), .A3(KEYINPUT84), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n593), .B(new_n594), .C1(new_n534), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(new_n529), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n590), .A2(new_n591), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n552), .A2(G85), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n543), .A2(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n549), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n523), .C2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n552), .A2(G92), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(KEYINPUT10), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n534), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n543), .A2(G54), .B1(G651), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n604), .A2(KEYINPUT10), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  OR2_X1    g195(.A1(new_n562), .A2(G868), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n611), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g199(.A(new_n495), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n625), .A2(KEYINPUT85), .A3(G123), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(new_n464), .B2(G111), .ZN(new_n627));
  INV_X1    g202(.A(G99), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n464), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n480), .B2(G135), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n495), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n626), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n465), .A2(new_n515), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2435), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2438), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2451), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n651), .B(new_n652), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G14), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2096), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(G2100), .Z(new_n664));
  INV_X1    g239(.A(KEYINPUT17), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n658), .B2(new_n659), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n661), .B1(new_n660), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT88), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT19), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  INV_X1    g255(.A(new_n678), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n672), .A2(new_n681), .A3(new_n675), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT90), .B(KEYINPUT91), .Z(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n690), .ZN(G229));
  NOR2_X1   g266(.A1(G16), .A2(G23), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n588), .B2(G16), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G22), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G1971), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n695), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT34), .Z(new_n705));
  MUX2_X1   g280(.A(G24), .B(G290), .S(G16), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT92), .ZN(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  INV_X1    g287(.A(G131), .ZN(new_n713));
  NOR2_X1   g288(.A1(G95), .A2(G2105), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(new_n464), .B2(G107), .ZN(new_n715));
  OAI22_X1  g290(.A1(new_n482), .A2(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n625), .B2(G119), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n712), .B1(new_n717), .B2(new_n711), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT35), .B(G1991), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NOR4_X1   g296(.A1(new_n709), .A2(new_n710), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n705), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT36), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT36), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n705), .A2(new_n726), .A3(new_n722), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n711), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n711), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G2090), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT101), .Z(new_n733));
  NOR2_X1   g308(.A1(G29), .A2(G33), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G139), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n515), .A2(G103), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  AOI22_X1  g312(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT95), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n735), .B(new_n737), .C1(new_n739), .C2(new_n464), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT96), .Z(new_n741));
  AOI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(G29), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G2072), .Z(new_n743));
  NAND2_X1  g318(.A1(G168), .A2(G16), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G16), .B2(G21), .ZN(new_n745));
  INV_X1    g320(.A(G1966), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G32), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n480), .A2(G141), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT26), .Z(new_n751));
  INV_X1    g326(.A(G129), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n495), .B2(new_n752), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n749), .B(new_n753), .C1(G105), .C2(new_n515), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT27), .B(G1996), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G28), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT99), .Z(new_n760));
  OAI211_X1 g335(.A(new_n760), .B(new_n711), .C1(new_n758), .C2(G28), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n747), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n755), .A2(new_n756), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n634), .A2(new_n711), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n731), .A2(G2090), .ZN(new_n766));
  INV_X1    g341(.A(G2078), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n519), .A2(G29), .A3(new_n520), .ZN(new_n768));
  INV_X1    g343(.A(G27), .ZN(new_n769));
  OAI21_X1  g344(.A(KEYINPUT100), .B1(new_n769), .B2(G29), .ZN(new_n770));
  OR3_X1    g345(.A1(new_n769), .A2(KEYINPUT100), .A3(G29), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n766), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n733), .A2(new_n743), .A3(new_n765), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G4), .A2(G16), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n612), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT94), .B(G1348), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n696), .A2(G19), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n562), .B2(new_n696), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G1341), .Z(new_n782));
  XOR2_X1   g357(.A(KEYINPUT31), .B(G11), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT98), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n782), .B(new_n784), .C1(new_n746), .C2(new_n745), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n777), .A2(new_n778), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n775), .A2(new_n779), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n772), .A2(G2078), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n711), .A2(G26), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n791));
  INV_X1    g366(.A(G140), .ZN(new_n792));
  INV_X1    g367(.A(G128), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n791), .B1(new_n792), .B2(new_n482), .C1(new_n495), .C2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(new_n711), .ZN(new_n796));
  MUX2_X1   g371(.A(new_n789), .B(new_n796), .S(KEYINPUT28), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2067), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n696), .A2(G5), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G171), .B2(new_n696), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1961), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n728), .A2(new_n787), .A3(new_n788), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(new_n711), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G160), .B2(new_n711), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2084), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n696), .A2(KEYINPUT23), .A3(G20), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT23), .ZN(new_n810));
  INV_X1    g385(.A(G20), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G16), .ZN(new_n812));
  INV_X1    g387(.A(G299), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n809), .B(new_n812), .C1(new_n813), .C2(new_n696), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT102), .B(G1956), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n803), .A2(new_n808), .A3(new_n817), .ZN(G311));
  OR3_X1    g393(.A1(new_n803), .A2(new_n808), .A3(new_n817), .ZN(G150));
  NAND2_X1  g394(.A1(new_n552), .A2(G93), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n543), .A2(G55), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n549), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n820), .B(new_n821), .C1(new_n523), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  OR2_X1    g400(.A1(new_n562), .A2(new_n823), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n562), .A2(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n611), .A2(new_n619), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n825), .B1(new_n832), .B2(G860), .ZN(G145));
  XNOR2_X1  g408(.A(new_n517), .B(new_n794), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n754), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT103), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(KEYINPUT103), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n741), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT104), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n835), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n740), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n839), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n845));
  INV_X1    g420(.A(G106), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n464), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n625), .B2(G130), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n849));
  INV_X1    g424(.A(G142), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n482), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n480), .A2(KEYINPUT105), .A3(G142), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n848), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(new_n637), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n717), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n844), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(G160), .B(new_n634), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n502), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n844), .A2(new_n856), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT106), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n844), .A2(new_n863), .A3(new_n855), .ZN(new_n864));
  INV_X1    g439(.A(new_n859), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n855), .A2(new_n863), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n840), .A2(new_n842), .A3(new_n843), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT40), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT40), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n861), .A2(new_n871), .A3(new_n862), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(G395));
  NAND2_X1  g448(.A1(new_n823), .A2(new_n615), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n588), .B(G290), .ZN(new_n875));
  XNOR2_X1  g450(.A(G166), .B(G305), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT107), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(KEYINPUT42), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(KEYINPUT42), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n828), .B(new_n622), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n611), .B(new_n813), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n885), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n886), .B1(new_n889), .B2(new_n884), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n883), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n874), .B1(new_n891), .B2(new_n615), .ZN(G295));
  OAI21_X1  g467(.A(new_n874), .B1(new_n891), .B2(new_n615), .ZN(G331));
  NOR2_X1   g468(.A1(G168), .A2(G301), .ZN(new_n894));
  NOR2_X1   g469(.A1(G286), .A2(G171), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n828), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n828), .B1(new_n894), .B2(new_n895), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n885), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n900), .A2(KEYINPUT108), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n899), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n888), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n900), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n906), .B2(new_n879), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n879), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT43), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT110), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n914), .A3(KEYINPUT43), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n906), .A2(new_n879), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT108), .B1(new_n903), .B2(new_n900), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n909), .B1(new_n918), .B2(new_n901), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n919), .A3(new_n862), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT44), .B1(new_n920), .B2(KEYINPUT43), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n907), .A2(new_n923), .A3(new_n910), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI22_X1  g500(.A1(new_n916), .A2(new_n921), .B1(KEYINPUT44), .B2(new_n925), .ZN(G397));
  INV_X1    g501(.A(G8), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT114), .ZN(new_n928));
  INV_X1    g503(.A(new_n468), .ZN(new_n929));
  XNOR2_X1  g504(.A(KEYINPUT112), .B(G40), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n492), .B1(new_n491), .B2(new_n472), .ZN(new_n931));
  AOI211_X1 g506(.A(KEYINPUT74), .B(new_n471), .C1(new_n489), .C2(new_n490), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n934));
  INV_X1    g509(.A(G1384), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n519), .A2(new_n935), .A3(new_n520), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G1384), .B1(new_n511), .B2(new_n516), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT45), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n928), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n934), .ZN(new_n941));
  INV_X1    g516(.A(new_n933), .ZN(new_n942));
  AND4_X1   g517(.A1(new_n928), .A2(new_n941), .A3(new_n942), .A4(new_n939), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n699), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n933), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n936), .A2(KEYINPUT50), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(G2090), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n927), .B1(new_n944), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(G166), .A2(new_n927), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT55), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n957), .B(new_n958), .C1(KEYINPUT55), .C2(new_n954), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT63), .B1(new_n953), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n941), .A2(new_n942), .A3(new_n939), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT114), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n941), .A2(new_n942), .A3(new_n928), .A4(new_n939), .ZN(new_n963));
  AOI21_X1  g538(.A(G1971), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(G8), .B(new_n959), .C1(new_n964), .C2(new_n951), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n517), .A2(new_n935), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n933), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(new_n927), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n588), .A2(G1976), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n971));
  NAND2_X1  g546(.A1(G305), .A2(G1981), .ZN(new_n972));
  INV_X1    g547(.A(G1981), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n590), .A2(new_n591), .A3(new_n973), .A4(new_n597), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT116), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT49), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n972), .B(KEYINPUT49), .C1(new_n976), .C2(new_n977), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n968), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1976), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(G288), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n984), .A2(new_n968), .A3(new_n969), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n971), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n965), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n960), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT119), .B(G2084), .Z(new_n989));
  NAND3_X1  g564(.A1(new_n948), .A2(new_n989), .A3(new_n949), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT120), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n966), .A2(new_n934), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n942), .B(new_n993), .C1(new_n934), .C2(new_n936), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n746), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n948), .A2(KEYINPUT120), .A3(new_n989), .A4(new_n949), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n997), .A2(G8), .A3(G168), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n519), .A2(new_n945), .A3(new_n935), .A4(new_n520), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n966), .A2(KEYINPUT50), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(G160), .A3(new_n930), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT118), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G2090), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n942), .A2(KEYINPUT118), .A3(new_n1000), .A4(new_n999), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(G8), .B1(new_n964), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n959), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(new_n965), .A3(new_n986), .A4(new_n998), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT63), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n988), .A2(new_n998), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n965), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n986), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n982), .A2(new_n983), .A3(new_n588), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n976), .A2(new_n977), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT117), .ZN(new_n1018));
  INV_X1    g593(.A(new_n968), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT121), .B1(new_n1012), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n997), .A2(G286), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n992), .A2(new_n995), .A3(G168), .A4(new_n996), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1022), .A2(KEYINPUT51), .A3(G8), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(G8), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT62), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n927), .B1(new_n944), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n965), .B(new_n986), .C1(new_n1031), .C2(new_n959), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n962), .A2(new_n767), .A3(new_n963), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OR3_X1    g610(.A1(new_n994), .A2(new_n1034), .A3(G2078), .ZN(new_n1036));
  INV_X1    g611(.A(new_n950), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1037), .A2(G1961), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1032), .A2(G301), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1029), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n966), .B(KEYINPUT111), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n934), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1034), .A2(G2078), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n939), .A2(G40), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1043), .A2(G160), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1035), .A2(new_n1038), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT126), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1035), .A2(KEYINPUT126), .A3(new_n1038), .A4(new_n1046), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(G171), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1039), .B2(G301), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1032), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1035), .A2(G301), .A3(new_n1038), .A4(new_n1046), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n1039), .B2(G301), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1028), .B1(new_n1056), .B2(new_n1052), .ZN(new_n1057));
  INV_X1    g632(.A(G1956), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1001), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n576), .A2(new_n1060), .A3(new_n578), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n813), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(G299), .A2(new_n1062), .A3(new_n1061), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n941), .A2(new_n942), .A3(new_n939), .A4(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1059), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1059), .A2(new_n1068), .A3(KEYINPUT61), .A4(new_n1066), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1348), .ZN(new_n1074));
  INV_X1    g649(.A(new_n949), .ZN(new_n1075));
  NAND3_X1  g650(.A1(G160), .A2(new_n930), .A3(new_n946), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n933), .A2(G2067), .A3(new_n966), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(KEYINPUT60), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT60), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1348), .B1(new_n948), .B2(new_n949), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n1078), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1083), .A3(new_n612), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1059), .A2(new_n1068), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1066), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1077), .A2(KEYINPUT60), .A3(new_n611), .A4(new_n1079), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1073), .A2(new_n1084), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT58), .B(G1341), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n961), .A2(G1996), .B1(new_n967), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n562), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n562), .A3(new_n1093), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1099));
  AOI211_X1 g674(.A(KEYINPUT123), .B(new_n1066), .C1(new_n1059), .C2(new_n1068), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n611), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1069), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1089), .A2(new_n1097), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT125), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n1106));
  OAI221_X1 g681(.A(new_n1106), .B1(new_n1102), .B2(new_n1103), .C1(new_n1089), .C2(new_n1097), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1054), .A2(new_n1057), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n998), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1011), .B1(new_n1032), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(G8), .B1(new_n964), .B2(new_n951), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1011), .B1(new_n1111), .B2(new_n1008), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1112), .A2(new_n965), .A3(new_n986), .A4(new_n998), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1017), .B(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1117), .A2(new_n968), .B1(new_n1013), .B2(new_n986), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1021), .A2(new_n1041), .A3(new_n1108), .A4(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1042), .A2(new_n934), .A3(new_n942), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n717), .B(new_n719), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1121), .B1(KEYINPUT113), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(KEYINPUT113), .B2(new_n1123), .ZN(new_n1125));
  INV_X1    g700(.A(G2067), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n794), .B(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n754), .B(G1996), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1121), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1121), .ZN(new_n1132));
  XNOR2_X1  g707(.A(G290), .B(G1986), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1120), .A2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1121), .A2(G1986), .A3(G290), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(KEYINPUT48), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1136), .A2(KEYINPUT48), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1131), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(G1996), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1132), .A2(KEYINPUT46), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT46), .B1(new_n1132), .B2(new_n1140), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1121), .B1(new_n754), .B2(new_n1127), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT47), .ZN(new_n1145));
  INV_X1    g720(.A(new_n719), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n717), .A2(new_n1146), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1129), .A2(new_n1147), .B1(G2067), .B2(new_n794), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT127), .Z(new_n1149));
  AOI211_X1 g724(.A(new_n1139), .B(new_n1145), .C1(new_n1132), .C2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1135), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g726(.A(new_n462), .B1(new_n922), .B2(new_n924), .ZN(new_n1153));
  NOR2_X1   g727(.A1(G229), .A2(G227), .ZN(new_n1154));
  NAND4_X1  g728(.A1(new_n1153), .A2(new_n869), .A3(new_n654), .A4(new_n1154), .ZN(G225));
  INV_X1    g729(.A(G225), .ZN(G308));
endmodule


