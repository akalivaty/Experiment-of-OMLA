//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT65), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G137), .ZN(new_n461));
  INV_X1    g036(.A(G101), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(G2104), .ZN(new_n463));
  OAI22_X1  g038(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(KEYINPUT66), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n465), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n464), .B1(new_n477), .B2(G2105), .ZN(G160));
  AOI21_X1  g053(.A(new_n459), .B1(new_n472), .B2(new_n473), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n480), .B(new_n482), .C1(new_n483), .C2(new_n460), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  AND2_X1   g060(.A1(new_n459), .A2(G138), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n469), .A2(new_n474), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n458), .A2(KEYINPUT4), .A3(new_n486), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n459), .B2(G114), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n494), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  AOI211_X1 g076(.A(new_n501), .B(new_n494), .C1(new_n496), .C2(new_n498), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n458), .A2(KEYINPUT67), .A3(G126), .A4(G2105), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n493), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n507), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n510), .B(KEYINPUT70), .C1(new_n500), .C2(new_n502), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n492), .B1(new_n509), .B2(new_n511), .ZN(G164));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(G50), .ZN(new_n525));
  INV_X1    g100(.A(new_n522), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  OAI211_X1 g102(.A(G50), .B(G543), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT71), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n521), .A2(new_n522), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT5), .B(G543), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G88), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n530), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n535), .B1(new_n530), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n519), .B1(new_n536), .B2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND3_X1  g114(.A1(new_n532), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n523), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n531), .A2(new_n532), .ZN(new_n544));
  INV_X1    g119(.A(G89), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n540), .B(new_n541), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(G168));
  NAND2_X1  g125(.A1(new_n523), .A2(G52), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(new_n544), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G651), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n553), .A2(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n531), .A2(G543), .ZN(new_n560));
  XOR2_X1   g135(.A(KEYINPUT74), .B(G43), .Z(new_n561));
  OAI22_X1  g136(.A1(new_n544), .A2(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n532), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n555), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g143(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n569));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n516), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(new_n578), .A3(G651), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT9), .B1(new_n560), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n523), .A2(new_n582), .A3(G53), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n581), .A2(new_n583), .B1(G91), .B2(new_n533), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n579), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G168), .ZN(G286));
  NAND2_X1  g161(.A1(new_n523), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n531), .A2(new_n532), .A3(G87), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n516), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G48), .B2(new_n523), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n531), .A2(new_n532), .A3(G86), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT77), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n533), .A2(new_n597), .A3(G86), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n594), .A2(new_n596), .A3(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(new_n523), .A2(G47), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n544), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n555), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  OR3_X1    g182(.A1(G171), .A2(KEYINPUT78), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT78), .B1(G171), .B2(new_n607), .ZN(new_n609));
  AND3_X1   g184(.A1(new_n531), .A2(new_n532), .A3(G92), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n516), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(G54), .B2(new_n523), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n608), .B(new_n609), .C1(G868), .C2(new_n617), .ZN(G284));
  OAI211_X1 g193(.A(new_n608), .B(new_n609), .C1(G868), .C2(new_n617), .ZN(G321));
  NAND2_X1  g194(.A1(G299), .A2(new_n607), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G168), .B2(new_n607), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(G168), .B2(new_n607), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n565), .A2(new_n607), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n616), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(new_n460), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G135), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT80), .ZN(new_n634));
  AOI211_X1 g209(.A(new_n631), .B(new_n634), .C1(G123), .C2(new_n479), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n475), .A2(new_n463), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G2100), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n636), .A2(new_n642), .A3(new_n643), .ZN(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  INV_X1    g242(.A(new_n660), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n667), .B1(new_n663), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n674), .A2(new_n679), .A3(new_n677), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n679), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n682));
  AOI211_X1 g257(.A(new_n678), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT83), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  NOR2_X1   g269(.A1(G16), .A2(G19), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n566), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1341), .ZN(new_n697));
  INV_X1    g272(.A(G11), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT31), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(KEYINPUT31), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n701), .A2(G28), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n701), .B2(G28), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n699), .B(new_n700), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n635), .B2(G29), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G5), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G171), .B2(new_n707), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n617), .A2(G16), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G4), .B2(G16), .ZN(new_n711));
  INV_X1    g286(.A(G1348), .ZN(new_n712));
  OAI221_X1 g287(.A(new_n706), .B1(G1961), .B2(new_n709), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n697), .B(new_n713), .C1(G1961), .C2(new_n709), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n703), .A2(G26), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n479), .A2(G128), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT87), .Z(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n719));
  INV_X1    g294(.A(G116), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G2105), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n632), .B2(G140), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2067), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n703), .B1(new_n727), .B2(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n727), .B2(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G160), .B2(G29), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n726), .B1(G2084), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G2078), .ZN(new_n732));
  NOR2_X1   g307(.A1(G164), .A2(new_n703), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G27), .B2(new_n703), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n714), .B(new_n731), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n703), .A2(G33), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n737));
  NAND2_X1  g312(.A1(G103), .A2(G2104), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G2105), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n632), .A2(G139), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n469), .A2(new_n474), .A3(G127), .ZN(new_n742));
  NAND2_X1  g317(.A1(G115), .A2(G2104), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n459), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n745), .B2(new_n744), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n736), .B1(new_n747), .B2(new_n703), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G2072), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n734), .A2(new_n732), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n730), .A2(G2084), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT90), .Z(new_n752));
  NAND3_X1  g327(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n479), .A2(G129), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT89), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT26), .Z(new_n757));
  INV_X1    g332(.A(G105), .ZN(new_n758));
  INV_X1    g333(.A(G141), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n757), .B1(new_n758), .B2(new_n463), .C1(new_n460), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(new_n703), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n703), .B2(G32), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT27), .B(G1996), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n703), .A2(G35), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT91), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n703), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2090), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n768), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n707), .A2(G21), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G168), .B2(new_n707), .ZN(new_n774));
  INV_X1    g349(.A(G1966), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n707), .A2(G20), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT23), .Z(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G299), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1956), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n712), .A2(new_n711), .B1(new_n763), .B2(new_n764), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n772), .A2(new_n776), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n735), .A2(new_n753), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n707), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n707), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT86), .Z(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G1971), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(G1971), .ZN(new_n789));
  MUX2_X1   g364(.A(G6), .B(G305), .S(G16), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT85), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT32), .B(G1981), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(new_n793), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n707), .A2(G23), .ZN(new_n796));
  INV_X1    g371(.A(G288), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n707), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT33), .ZN(new_n799));
  INV_X1    g374(.A(G1976), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n794), .A2(new_n795), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n788), .A2(new_n789), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT34), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n788), .A2(new_n805), .A3(new_n789), .A4(new_n802), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n703), .A2(G25), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n632), .A2(G131), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n479), .A2(G119), .ZN(new_n809));
  OR2_X1    g384(.A1(G95), .A2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(new_n703), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT35), .B(G1991), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G16), .A2(G24), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n605), .B(KEYINPUT84), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G16), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G1986), .Z(new_n820));
  NAND4_X1  g395(.A1(new_n804), .A2(new_n806), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n784), .B1(new_n822), .B2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n783), .ZN(G150));
  NAND2_X1  g401(.A1(new_n565), .A2(KEYINPUT96), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT97), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n533), .A2(G93), .B1(G55), .B2(new_n523), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n532), .A2(G67), .ZN(new_n830));
  NAND2_X1  g405(.A1(G80), .A2(G543), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n555), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n829), .B1(KEYINPUT95), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(KEYINPUT95), .B2(new_n832), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(KEYINPUT96), .B2(new_n565), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n828), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n828), .A2(new_n835), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n617), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT94), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n838), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n841), .B(new_n842), .Z(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n843), .B2(KEYINPUT39), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n843), .A2(KEYINPUT98), .A3(KEYINPUT39), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n841), .B(new_n842), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n844), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G860), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n834), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(G145));
  XNOR2_X1  g429(.A(new_n747), .B(new_n723), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n761), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n479), .A2(G130), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT100), .Z(new_n859));
  INV_X1    g434(.A(G118), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(KEYINPUT101), .A3(G2105), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT101), .B1(new_n860), .B2(G2105), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n632), .A2(G142), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(new_n638), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n638), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n812), .ZN(new_n872));
  INV_X1    g447(.A(new_n494), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n497), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT68), .B1(new_n497), .B2(G2105), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n501), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n499), .A2(KEYINPUT69), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n877), .A2(new_n878), .B1(new_n506), .B2(new_n507), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n490), .B1(new_n488), .B2(new_n487), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n869), .A2(new_n813), .A3(new_n870), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n872), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n881), .B1(new_n872), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n857), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n872), .A2(new_n882), .ZN(new_n886));
  INV_X1    g461(.A(new_n881), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n872), .A2(new_n881), .A3(new_n882), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n856), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(G160), .B(KEYINPUT99), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G162), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(new_n635), .Z(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n885), .A2(new_n890), .A3(new_n894), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n896), .A2(KEYINPUT40), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT40), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(G395));
  OR2_X1    g475(.A1(new_n834), .A2(G868), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n838), .B(new_n626), .ZN(new_n902));
  XOR2_X1   g477(.A(G299), .B(new_n616), .Z(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n903), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n906), .B1(new_n907), .B2(new_n902), .ZN(new_n908));
  XNOR2_X1  g483(.A(G303), .B(G290), .ZN(new_n909));
  XOR2_X1   g484(.A(G288), .B(KEYINPUT103), .Z(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(G305), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n909), .B(new_n911), .Z(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT104), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT42), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n908), .B(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n901), .B1(new_n915), .B2(new_n607), .ZN(G295));
  OAI21_X1  g491(.A(new_n901), .B1(new_n915), .B2(new_n607), .ZN(G331));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  OAI21_X1  g493(.A(G168), .B1(new_n918), .B2(G301), .ZN(new_n919));
  NAND2_X1  g494(.A1(G301), .A2(new_n918), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n838), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n836), .A2(new_n921), .A3(new_n837), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n905), .ZN(new_n926));
  INV_X1    g501(.A(new_n912), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n903), .A3(new_n924), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n927), .B1(new_n926), .B2(new_n928), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT43), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n930), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n905), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n907), .A2(new_n936), .A3(KEYINPUT41), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n925), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n927), .B1(new_n939), .B2(new_n928), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n935), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n934), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n931), .B2(new_n933), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n935), .A2(new_n940), .A3(KEYINPUT43), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(G397));
  XNOR2_X1  g523(.A(new_n723), .B(new_n725), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT108), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n761), .ZN(new_n951));
  INV_X1    g526(.A(G1996), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(KEYINPUT107), .B(G40), .Z(new_n954));
  NAND2_X1  g529(.A1(G160), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n879), .B2(new_n880), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT45), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n951), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n952), .A3(new_n761), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n813), .A2(new_n815), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n813), .A2(new_n815), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n957), .ZN(new_n964));
  NOR2_X1   g539(.A1(G290), .A2(G1986), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G290), .A2(G1986), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(G160), .A2(new_n954), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n956), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n971), .A2(G2067), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n510), .B1(new_n500), .B2(new_n502), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n974), .B(new_n975), .C1(new_n976), .C2(new_n492), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n956), .A2(KEYINPUT109), .A3(new_n974), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n973), .A2(new_n981), .A3(new_n970), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n972), .B1(new_n982), .B2(new_n712), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n983), .A2(KEYINPUT60), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n712), .ZN(new_n985));
  INV_X1    g560(.A(new_n972), .ZN(new_n986));
  AND4_X1   g561(.A1(KEYINPUT60), .A2(new_n985), .A3(new_n616), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n616), .B1(new_n983), .B2(KEYINPUT60), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(G299), .A2(KEYINPUT57), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(G299), .A2(KEYINPUT57), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G164), .B2(G1384), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n955), .B1(KEYINPUT45), .B2(new_n956), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT56), .B(G2072), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n511), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n877), .A2(new_n878), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT70), .B1(new_n1001), .B2(new_n510), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n880), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1003), .A2(new_n974), .A3(new_n975), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n881), .A2(new_n975), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n955), .B1(new_n1005), .B2(KEYINPUT50), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1956), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n993), .B1(new_n999), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n993), .ZN(new_n1009));
  NOR3_X1   g584(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n970), .B1(new_n974), .B2(new_n956), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1009), .B(new_n998), .C1(new_n1012), .C2(G1956), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT61), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1008), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n999), .A2(new_n1007), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(KEYINPUT61), .A3(new_n1009), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n995), .A2(new_n952), .A3(new_n996), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(G1341), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n971), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n565), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT59), .ZN(new_n1025));
  XOR2_X1   g600(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1026));
  AOI211_X1 g601(.A(new_n565), .B(new_n1026), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n989), .A2(new_n1018), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n998), .B1(new_n1012), .B2(G1956), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n993), .A2(KEYINPUT117), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n991), .A2(new_n1032), .A3(new_n992), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(KEYINPUT118), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n616), .B2(new_n983), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT118), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1013), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1005), .A2(new_n994), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n956), .A2(KEYINPUT45), .ZN(new_n1040));
  NAND4_X1  g615(.A1(G160), .A2(KEYINPUT53), .A3(G40), .A4(new_n732), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n995), .A2(new_n732), .A3(new_n996), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT125), .ZN(new_n1046));
  INV_X1    g621(.A(G1961), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n982), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1046), .B1(new_n982), .B2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT127), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT127), .B(new_n1045), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(G171), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1003), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n955), .B1(new_n1005), .B2(new_n994), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n732), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1056), .A2(KEYINPUT123), .A3(new_n732), .A4(new_n1057), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT53), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n982), .A2(new_n1047), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1055), .B1(new_n1067), .B2(G301), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1029), .A2(new_n1038), .B1(new_n1054), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT126), .ZN(new_n1070));
  AND3_X1   g645(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT116), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1004), .A2(new_n1076), .A3(new_n1006), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT110), .B(G2090), .Z(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1971), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT45), .B1(new_n1003), .B2(new_n975), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n970), .B1(new_n1005), .B2(new_n994), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1074), .B1(new_n1084), .B2(G8), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n973), .A2(new_n981), .A3(new_n970), .A4(new_n1078), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(G8), .A3(new_n1074), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(G1976), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(G8), .B(new_n1091), .C1(new_n1005), .C2(new_n955), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT52), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n800), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1981), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n594), .A2(new_n598), .A3(new_n1097), .A4(new_n596), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n523), .A2(G48), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n532), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1099), .B(new_n595), .C1(new_n1100), .C2(new_n555), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G1981), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT49), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT112), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1106), .B(KEYINPUT49), .C1(new_n1098), .C2(new_n1102), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1098), .A2(KEYINPUT49), .A3(new_n1102), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n971), .A2(G8), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n971), .A2(G8), .A3(new_n1109), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT113), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1096), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1088), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1070), .B1(new_n1085), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1088), .A2(new_n1116), .ZN(new_n1119));
  AOI21_X1  g694(.A(G1971), .B1(new_n995), .B2(new_n996), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1078), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(KEYINPUT116), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1120), .B1(new_n1123), .B2(new_n1077), .ZN(new_n1124));
  INV_X1    g699(.A(G8), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1073), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1119), .A2(new_n1126), .A3(KEYINPUT126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT122), .B(KEYINPUT51), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n775), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n955), .A2(G2084), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n973), .A2(new_n981), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1125), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(G286), .A2(G8), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT121), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1128), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1132), .ZN(new_n1137));
  AOI21_X1  g712(.A(G1966), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1138));
  OAI21_X1  g713(.A(G8), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1135), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(KEYINPUT51), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1136), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1118), .A2(new_n1127), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(G171), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT124), .B(G171), .C1(new_n1063), .C2(new_n1066), .ZN(new_n1148));
  OAI211_X1 g723(.A(G301), .B(new_n1045), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1055), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1069), .A2(new_n1144), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1133), .A2(G168), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1087), .A2(G8), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1073), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1119), .A2(KEYINPUT63), .A3(new_n1154), .A4(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1085), .A2(new_n1117), .A3(new_n1153), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(KEYINPUT63), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n797), .A2(new_n800), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT115), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1098), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1125), .B1(new_n970), .B2(new_n956), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT114), .Z(new_n1165));
  INV_X1    g740(.A(new_n1088), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1163), .A2(new_n1165), .B1(new_n1166), .B2(new_n1116), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1136), .A2(new_n1141), .A3(new_n1169), .A4(new_n1142), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1143), .A2(KEYINPUT62), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1118), .A2(new_n1127), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1159), .B(new_n1167), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n969), .B1(new_n1152), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n957), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n957), .A2(new_n952), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT46), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT47), .Z(new_n1180));
  NAND3_X1  g755(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n718), .A2(new_n725), .A3(new_n722), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n964), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n965), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT48), .Z(new_n1185));
  NOR2_X1   g760(.A1(new_n963), .A2(new_n1185), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1180), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1175), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g763(.A(G319), .ZN(new_n1190));
  NOR3_X1   g764(.A1(G401), .A2(new_n1190), .A3(G227), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n693), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1192), .B1(new_n896), .B2(new_n897), .ZN(new_n1193));
  INV_X1    g767(.A(new_n940), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n931), .A2(new_n1194), .A3(new_n941), .ZN(new_n1195));
  OAI21_X1  g769(.A(KEYINPUT43), .B1(new_n935), .B2(new_n932), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AND2_X1   g771(.A1(new_n1193), .A2(new_n1197), .ZN(G308));
  NAND2_X1  g772(.A1(new_n1193), .A2(new_n1197), .ZN(G225));
endmodule


