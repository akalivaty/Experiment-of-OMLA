//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT65), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G58), .ZN(new_n208));
  INV_X1    g0008(.A(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G116), .A2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n205), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G50), .C2(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT67), .B(G68), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  NOR2_X1   g0026(.A1(new_n224), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n220), .B(new_n228), .C1(new_n211), .C2(new_n216), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI22_X1  g0036(.A1(new_n229), .A2(KEYINPUT0), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n226), .B(new_n237), .C1(KEYINPUT0), .C2(new_n229), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  XOR2_X1   g0054(.A(KEYINPUT8), .B(G58), .Z(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n230), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n256), .A2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n259), .B1(new_n264), .B2(new_n255), .ZN(new_n265));
  INV_X1    g0065(.A(new_n222), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n202), .B1(new_n266), .B2(G58), .ZN(new_n267));
  INV_X1    g0067(.A(G159), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n231), .A2(new_n269), .A3(KEYINPUT70), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT70), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G20), .B2(G33), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n267), .A2(new_n231), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT7), .ZN(new_n275));
  OR2_X1    g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n278), .B2(G20), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n274), .B1(G68), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n262), .B1(new_n285), .B2(KEYINPUT16), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT16), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n222), .B1(new_n279), .B2(new_n283), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n274), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n265), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT78), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  AND2_X1   g0092(.A1(G1), .A2(G13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G226), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G1698), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n278), .B(new_n297), .C1(G223), .C2(G1698), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G87), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G41), .ZN(new_n301));
  INV_X1    g0101(.A(G45), .ZN(new_n302));
  AOI21_X1  g0102(.A(G1), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT68), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n304), .A2(new_n305), .A3(new_n230), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT68), .B1(new_n293), .B2(new_n294), .ZN(new_n307));
  OAI211_X1 g0107(.A(G274), .B(new_n303), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n303), .ZN(new_n309));
  OAI211_X1 g0109(.A(G232), .B(new_n309), .C1(new_n306), .C2(new_n307), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT76), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT76), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n308), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n300), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT77), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n300), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n308), .A2(new_n310), .A3(new_n313), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n313), .B1(new_n308), .B2(new_n310), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n316), .B(new_n318), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n292), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(G190), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n291), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(KEYINPUT77), .ZN(new_n328));
  AOI21_X1  g0128(.A(G200), .B1(new_n328), .B2(new_n321), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n329), .A2(KEYINPUT78), .A3(new_n325), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n290), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT17), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n286), .A2(new_n289), .ZN(new_n334));
  INV_X1    g0134(.A(new_n265), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n323), .A2(new_n291), .A3(new_n326), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT78), .B1(new_n329), .B2(new_n325), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT17), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n328), .A2(new_n321), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  INV_X1    g0142(.A(G179), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(new_n315), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n336), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT18), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(KEYINPUT18), .A3(new_n336), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n305), .B1(new_n304), .B2(new_n230), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n293), .A2(KEYINPUT68), .A3(new_n294), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n303), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G244), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n278), .B1(new_n209), .B2(G1698), .ZN(new_n354));
  INV_X1    g0154(.A(G1698), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n221), .A2(new_n355), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n354), .A2(new_n356), .B1(G107), .B2(new_n278), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n308), .B(new_n353), .C1(new_n357), .C2(new_n295), .ZN(new_n358));
  INV_X1    g0158(.A(G190), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n270), .A2(new_n272), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n255), .A2(new_n361), .B1(G20), .B2(G77), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT15), .B(G87), .Z(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n231), .A2(G33), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n261), .B1(new_n205), .B2(new_n258), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n262), .A2(G77), .A3(new_n263), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n358), .A2(G200), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n360), .A2(new_n367), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n358), .A2(G179), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(new_n368), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n358), .A2(new_n342), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n333), .A2(new_n340), .A3(new_n349), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT12), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n262), .B2(new_n263), .ZN(new_n380));
  INV_X1    g0180(.A(G68), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n222), .A2(G20), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n256), .A2(KEYINPUT12), .A3(G13), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G50), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n273), .A2(new_n385), .B1(new_n205), .B2(new_n365), .ZN(new_n386));
  INV_X1    g0186(.A(new_n382), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n261), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n388), .A2(KEYINPUT11), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(KEYINPUT11), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n384), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n257), .A2(new_n379), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n296), .A2(new_n355), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n278), .B(new_n395), .C1(G232), .C2(new_n355), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G97), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n295), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT13), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n352), .A2(G238), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n308), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n308), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT13), .B1(new_n403), .B2(new_n398), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n404), .A3(G190), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT74), .ZN(new_n406));
  OR4_X1    g0206(.A1(new_n406), .A2(new_n403), .A3(KEYINPUT13), .A4(new_n398), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(new_n404), .A3(new_n406), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(G200), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n394), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n393), .A2(KEYINPUT75), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT75), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n391), .A2(new_n413), .A3(new_n392), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n407), .A2(new_n408), .A3(G169), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT14), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n402), .A2(new_n404), .A3(G179), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n407), .A2(new_n408), .A3(new_n419), .A4(G169), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n411), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT71), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n263), .A2(new_n423), .A3(G50), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n423), .B1(new_n263), .B2(G50), .ZN(new_n426));
  NOR4_X1   g0226(.A1(new_n425), .A2(new_n426), .A3(new_n258), .A4(new_n261), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n255), .A2(new_n231), .A3(G33), .ZN(new_n428));
  INV_X1    g0228(.A(G150), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n428), .B1(new_n429), .B2(new_n273), .C1(new_n204), .C2(new_n231), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n427), .B1(new_n430), .B2(new_n261), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n258), .A2(new_n385), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT72), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT9), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n436), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n431), .A2(new_n438), .A3(new_n432), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g0240(.A1(KEYINPUT69), .A2(G223), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT69), .A2(G223), .ZN(new_n442));
  OAI21_X1  g0242(.A(G1698), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n355), .A2(G222), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n278), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n295), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n446), .C1(G77), .C2(new_n278), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n352), .A2(G226), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n308), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n359), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(G200), .B2(new_n449), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT73), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT10), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n434), .A2(new_n435), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n440), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n440), .B2(new_n456), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n449), .A2(new_n342), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n433), .B(new_n460), .C1(G179), .C2(new_n449), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n378), .A2(new_n422), .A3(new_n459), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT4), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G1698), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(G244), .C1(new_n281), .C2(new_n280), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n214), .B1(new_n276), .B2(new_n277), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n465), .B(new_n466), .C1(new_n467), .C2(KEYINPUT4), .ZN(new_n468));
  OAI21_X1  g0268(.A(G250), .B1(new_n280), .B2(new_n281), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n355), .B1(new_n469), .B2(KEYINPUT4), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n446), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n350), .A2(new_n351), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n302), .A2(G1), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n301), .A2(KEYINPUT5), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G41), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n472), .A2(G274), .A3(new_n477), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT5), .B(G41), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n350), .A2(new_n351), .B1(new_n479), .B2(new_n473), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G257), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n471), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n342), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n471), .A2(new_n343), .A3(new_n478), .A4(new_n481), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n258), .A2(new_n210), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n256), .A2(G33), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n262), .A2(new_n257), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(new_n210), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT7), .B1(new_n282), .B2(new_n231), .ZN(new_n490));
  NOR4_X1   g0290(.A1(new_n280), .A2(new_n281), .A3(new_n275), .A4(G20), .ZN(new_n491));
  OAI21_X1  g0291(.A(G107), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT79), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT79), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n284), .A2(new_n494), .A3(G107), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n215), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n210), .A2(new_n215), .ZN(new_n497));
  NOR2_X1   g0297(.A1(G97), .A2(G107), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n496), .B1(new_n499), .B2(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G20), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n361), .A2(G77), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n493), .A2(new_n495), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n489), .B1(new_n503), .B2(new_n261), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n485), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n482), .A2(new_n292), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n471), .A2(new_n359), .A3(new_n478), .A4(new_n481), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n220), .A2(new_n355), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n211), .A2(G1698), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n510), .B(new_n511), .C1(new_n280), .C2(new_n281), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n480), .A2(G264), .B1(new_n514), .B2(new_n446), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n478), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n292), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(G190), .B2(new_n516), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n231), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n231), .A2(G107), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n522), .B(KEYINPUT23), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT22), .ZN(new_n524));
  AOI21_X1  g0324(.A(G20), .B1(new_n276), .B2(new_n277), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(G87), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n231), .B(G87), .C1(new_n280), .C2(new_n281), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n521), .B(new_n523), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT24), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n278), .A2(new_n524), .A3(new_n231), .A4(G87), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n531), .A2(new_n532), .B1(new_n231), .B2(new_n520), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT24), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(new_n523), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n261), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n215), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT85), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT25), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n257), .B2(G107), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n539), .B(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n488), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G107), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n518), .A2(new_n537), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(G169), .B1(new_n515), .B2(new_n478), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n514), .A2(new_n446), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n479), .A2(new_n473), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n472), .A2(G264), .A3(new_n550), .ZN(new_n551));
  AND4_X1   g0351(.A1(new_n343), .A2(new_n549), .A3(new_n478), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n262), .B1(new_n530), .B2(new_n535), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n545), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n547), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n231), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT80), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n219), .A2(new_n210), .A3(new_n215), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(KEYINPUT80), .A3(new_n231), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n525), .A2(G68), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n365), .B2(new_n210), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT81), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT81), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n569), .B(new_n566), .C1(new_n365), .C2(new_n210), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n564), .A2(new_n565), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n261), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n543), .A2(new_n363), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n363), .A2(new_n257), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n221), .A2(new_n355), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n214), .A2(G1698), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(new_n578), .C1(new_n280), .C2(new_n281), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n519), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n446), .ZN(new_n581));
  AOI21_X1  g0381(.A(G250), .B1(new_n256), .B2(G45), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n302), .A2(G1), .A3(G274), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n585), .C1(new_n306), .C2(new_n307), .ZN(new_n586));
  AOI21_X1  g0386(.A(G169), .B1(new_n581), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n582), .B(new_n584), .C1(new_n350), .C2(new_n351), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n295), .B1(new_n579), .B2(new_n519), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n589), .A2(new_n590), .A3(G179), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n576), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT82), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n574), .B1(new_n571), .B2(new_n261), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n581), .A2(new_n586), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G200), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n543), .A2(G87), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n581), .A2(G190), .A3(new_n586), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n595), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n593), .A2(new_n594), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n594), .B1(new_n593), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n216), .A2(new_n355), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n211), .A2(G1698), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n604), .A2(new_n605), .B1(new_n281), .B2(new_n280), .ZN(new_n606));
  OR2_X1    g0406(.A1(KEYINPUT83), .A2(G303), .ZN(new_n607));
  NAND2_X1  g0407(.A1(KEYINPUT83), .A2(G303), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n276), .A2(new_n607), .A3(new_n277), .A4(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT84), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n606), .A2(KEYINPUT84), .A3(new_n609), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n446), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n472), .A2(G270), .A3(new_n550), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n478), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n615), .A3(G190), .ZN(new_n616));
  INV_X1    g0416(.A(G116), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n258), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n260), .A2(new_n230), .B1(G20), .B2(new_n617), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n466), .B(new_n231), .C1(G33), .C2(new_n210), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n619), .A2(KEYINPUT20), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT20), .B1(new_n619), .B2(new_n620), .ZN(new_n622));
  OAI221_X1 g0422(.A(new_n618), .B1(new_n488), .B2(new_n617), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n478), .A2(new_n614), .ZN(new_n625));
  INV_X1    g0425(.A(new_n612), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(new_n610), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n627), .B2(new_n446), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n616), .B(new_n624), .C1(new_n628), .C2(new_n292), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n623), .A2(G169), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n630), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n628), .A2(G179), .A3(new_n623), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n613), .A2(new_n615), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(KEYINPUT21), .A3(G169), .A4(new_n623), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n629), .A2(new_n632), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n509), .A2(new_n557), .A3(new_n603), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n462), .A2(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n462), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT86), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n586), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n582), .B1(new_n350), .B2(new_n351), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT86), .B1(new_n643), .B2(new_n585), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n581), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT87), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(new_n342), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n586), .A2(new_n641), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n643), .A2(KEYINPUT86), .A3(new_n585), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n590), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT87), .B1(new_n650), .B2(G169), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n591), .B1(new_n595), .B2(new_n573), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n572), .A2(new_n575), .A3(new_n598), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n596), .A2(new_n359), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(G200), .B2(new_n645), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n652), .A2(new_n653), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n555), .A2(new_n633), .A3(new_n635), .A4(new_n632), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n509), .A2(new_n547), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n646), .B1(new_n645), .B2(new_n342), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n650), .A2(KEYINPUT87), .A3(G169), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n653), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n658), .A2(new_n664), .A3(new_n505), .ZN(new_n665));
  AOI211_X1 g0465(.A(new_n587), .B(new_n591), .C1(new_n595), .C2(new_n573), .ZN(new_n666));
  AND4_X1   g0466(.A1(new_n595), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT82), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n593), .A2(new_n594), .A3(new_n600), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n503), .A2(new_n261), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n484), .B(new_n483), .C1(new_n671), .C2(new_n489), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT26), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n660), .A2(new_n663), .A3(new_n665), .A4(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n640), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n349), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n333), .A2(new_n340), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n421), .A2(new_n415), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT88), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n374), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT88), .A4(new_n373), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n678), .B1(new_n411), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n676), .B1(new_n677), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n459), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n461), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n675), .A2(new_n686), .ZN(G369));
  INV_X1    g0487(.A(G13), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G20), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n256), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT89), .Z(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(G213), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n554), .B2(new_n545), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n557), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT90), .ZN(new_n699));
  INV_X1    g0499(.A(new_n555), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n696), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n696), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n637), .B1(new_n624), .B2(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n632), .A2(new_n635), .A3(new_n633), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n696), .A2(new_n623), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT91), .Z(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n706), .A2(new_n696), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n699), .A2(new_n714), .B1(new_n700), .B2(new_n704), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(G399));
  NOR2_X1   g0516(.A1(new_n228), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G1), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n562), .A2(G116), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n719), .A2(new_n720), .B1(new_n235), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT94), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n674), .A2(new_n724), .A3(new_n704), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n724), .B1(new_n674), .B2(new_n704), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n634), .A2(new_n343), .A3(new_n645), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n482), .A2(new_n516), .ZN(new_n729));
  OR3_X1    g0529(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT93), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT93), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND4_X1   g0532(.A1(G179), .A2(new_n613), .A3(new_n615), .A4(new_n515), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n482), .A2(new_n596), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(KEYINPUT92), .A2(KEYINPUT30), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n735), .B(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n704), .B1(new_n732), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n508), .A2(new_n504), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n504), .B2(new_n485), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n556), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n603), .A3(new_n637), .A4(new_n704), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(new_n743), .B2(KEYINPUT31), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n728), .A2(new_n729), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n745), .B(new_n704), .C1(new_n738), .C2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(G330), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n659), .A2(new_n547), .A3(new_n658), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n741), .A2(KEYINPUT95), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT95), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n672), .A2(new_n751), .A3(new_n740), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n749), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n657), .A2(new_n655), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n663), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT26), .B1(new_n755), .B2(new_n672), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n668), .A2(new_n664), .A3(new_n505), .A4(new_n669), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(new_n663), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n704), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT29), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n727), .A2(new_n748), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT96), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n722), .B1(new_n763), .B2(G1), .ZN(G364));
  AOI21_X1  g0564(.A(new_n719), .B1(G45), .B2(new_n689), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n708), .A2(G330), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n710), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n228), .A2(new_n278), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n236), .A2(new_n302), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(new_n250), .C2(new_n302), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n228), .A2(new_n282), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(G355), .B(KEYINPUT97), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n771), .B1(G116), .B2(new_n227), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n230), .B1(G20), .B2(new_n342), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n778), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n708), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n231), .A2(G190), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G179), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G329), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  NOR2_X1   g0588(.A1(new_n343), .A2(new_n292), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n784), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n282), .B1(new_n786), .B2(new_n787), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n292), .A2(G179), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT99), .Z(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n791), .B1(new_n795), .B2(G283), .ZN(new_n796));
  INV_X1    g0596(.A(new_n784), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n797), .A2(new_n343), .A3(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G311), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT100), .B(G326), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n231), .A2(new_n359), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n789), .ZN(new_n803));
  INV_X1    g0603(.A(G294), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n231), .B1(new_n785), .B2(G190), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n801), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n802), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n807), .A2(new_n343), .A3(G200), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n806), .B1(G322), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n802), .A2(new_n792), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT101), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G303), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n796), .A2(new_n799), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n794), .A2(new_n215), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n798), .A2(KEYINPUT98), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n798), .A2(KEYINPUT98), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n815), .B1(new_n819), .B2(G77), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n805), .A2(new_n210), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n385), .B2(new_n803), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G58), .B2(new_n808), .ZN(new_n824));
  INV_X1    g0624(.A(new_n786), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G159), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT32), .Z(new_n827));
  INV_X1    g0627(.A(new_n810), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n282), .B1(new_n828), .B2(G87), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n820), .A2(new_n824), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n790), .A2(new_n381), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n814), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n783), .B1(new_n779), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n768), .B1(new_n833), .B2(new_n766), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT102), .Z(G396));
  NAND4_X1  g0635(.A1(new_n680), .A2(new_n372), .A3(new_n681), .A4(new_n696), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n696), .A2(new_n372), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n375), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OR3_X1    g0640(.A1(new_n725), .A2(new_n726), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n674), .A2(new_n704), .A3(new_n840), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(new_n748), .Z(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n766), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n794), .A2(new_n219), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G311), .B2(new_n825), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT103), .ZN(new_n848));
  INV_X1    g0648(.A(G283), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n282), .B1(new_n790), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n803), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G303), .ZN(new_n852));
  INV_X1    g0652(.A(new_n808), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n822), .B(new_n852), .C1(new_n853), .C2(new_n804), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n850), .B(new_n854), .C1(G107), .C2(new_n812), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n848), .B(new_n855), .C1(new_n617), .C2(new_n818), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT104), .Z(new_n857));
  NOR2_X1   g0657(.A1(new_n794), .A2(new_n381), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n278), .B1(new_n208), .B2(new_n805), .C1(new_n811), .C2(new_n385), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n808), .A2(G143), .B1(new_n851), .B2(G137), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n860), .B1(new_n429), .B2(new_n790), .C1(new_n818), .C2(new_n268), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n858), .B(new_n859), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(G132), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n863), .B1(new_n862), .B2(new_n861), .C1(new_n864), .C2(new_n786), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n857), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT105), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n766), .B1(new_n867), .B2(new_n779), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n779), .A2(new_n776), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n868), .B1(G77), .B2(new_n870), .C1(new_n777), .C2(new_n840), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n845), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(G384));
  OAI211_X1 g0673(.A(G77), .B(new_n236), .C1(new_n222), .C2(new_n208), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT106), .ZN(new_n875));
  INV_X1    g0675(.A(new_n201), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n875), .B1(new_n381), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(G1), .A3(new_n688), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n617), .B1(new_n500), .B2(KEYINPUT35), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n234), .C1(KEYINPUT35), .C2(new_n500), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT36), .ZN(new_n881));
  INV_X1    g0681(.A(new_n345), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n290), .A2(new_n694), .ZN(new_n883));
  NOR4_X1   g0683(.A1(new_n339), .A2(new_n882), .A3(KEYINPUT37), .A4(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n286), .B1(KEYINPUT16), .B2(new_n285), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n335), .ZN(new_n887));
  INV_X1    g0687(.A(new_n694), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n887), .B1(new_n344), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n885), .B1(new_n331), .B2(new_n889), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n333), .A2(new_n340), .A3(new_n349), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n694), .B1(new_n886), .B2(new_n335), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n892), .A2(KEYINPUT107), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT107), .B1(new_n892), .B2(new_n893), .ZN(new_n895));
  OAI211_X1 g0695(.A(KEYINPUT38), .B(new_n891), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n892), .A2(new_n883), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n882), .A2(new_n883), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n885), .B1(new_n899), .B2(new_n331), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n884), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n897), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n739), .A2(KEYINPUT31), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n744), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n415), .B(new_n696), .C1(new_n411), .C2(new_n421), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n415), .A2(new_n696), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n678), .A2(new_n908), .A3(new_n410), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n906), .A2(new_n839), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n903), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n912), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n897), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n914), .B1(new_n916), .B2(new_n896), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n913), .B1(new_n917), .B2(KEYINPUT40), .ZN(new_n918));
  INV_X1    g0718(.A(new_n906), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n640), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(G330), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n462), .B1(new_n727), .B2(new_n760), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n923), .A2(new_n686), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT108), .Z(new_n925));
  NAND3_X1  g0725(.A1(new_n916), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n903), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n678), .A2(new_n696), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n676), .A2(new_n694), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n916), .A2(new_n896), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n374), .A2(new_n696), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n842), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(new_n911), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n930), .A2(new_n931), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n925), .B(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n922), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n939), .A2(KEYINPUT109), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(KEYINPUT109), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n940), .B(new_n941), .C1(new_n938), .C2(new_n922), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n689), .A2(new_n256), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n878), .B(new_n881), .C1(new_n942), .C2(new_n943), .ZN(G367));
  NAND2_X1  g0744(.A1(new_n696), .A2(new_n654), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT110), .Z(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(new_n653), .A3(new_n652), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n755), .B2(new_n946), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(new_n782), .ZN(new_n949));
  INV_X1    g0749(.A(new_n769), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n780), .B1(new_n227), .B2(new_n364), .C1(new_n246), .C2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(G317), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n282), .B1(new_n786), .B2(new_n952), .C1(new_n804), .C2(new_n790), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n819), .B2(G283), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n607), .A2(new_n608), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n853), .A2(new_n955), .B1(new_n215), .B2(new_n805), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(G311), .B2(new_n851), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT46), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n812), .B2(G116), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n810), .A2(KEYINPUT46), .A3(new_n617), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n958), .B1(new_n210), .B2(new_n793), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n805), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(G68), .ZN(new_n964));
  INV_X1    g0764(.A(G143), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n964), .B1(new_n965), .B2(new_n803), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n278), .B1(new_n853), .B2(new_n429), .ZN(new_n967));
  INV_X1    g0767(.A(new_n790), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n966), .B(new_n967), .C1(G159), .C2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n793), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G77), .A2(new_n970), .B1(new_n825), .B2(G137), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n969), .B(new_n971), .C1(new_n201), .C2(new_n818), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n810), .A2(new_n208), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n962), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n766), .B1(new_n976), .B2(new_n779), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n949), .A2(new_n951), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n750), .A2(new_n752), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n504), .B2(new_n704), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n672), .B2(new_n704), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT111), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n712), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n700), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n696), .B1(new_n986), .B2(new_n672), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n699), .A2(new_n714), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(new_n981), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT42), .Z(new_n990));
  OAI211_X1 g0790(.A(new_n984), .B(new_n985), .C1(new_n987), .C2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n985), .B1(new_n987), .B2(new_n990), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(new_n712), .A3(new_n983), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n256), .B1(new_n689), .B2(G45), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n715), .A2(new_n982), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT44), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n715), .A2(new_n982), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT45), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n713), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1002), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1004), .A2(new_n712), .A3(new_n999), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n988), .B1(new_n703), .B2(new_n714), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n709), .B(KEYINPUT112), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n709), .A2(KEYINPUT112), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1010), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n762), .B1(new_n1006), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n717), .B(KEYINPUT41), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n997), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n979), .B1(new_n996), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(G387));
  INV_X1    g0819(.A(new_n997), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1013), .A2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G322), .A2(new_n851), .B1(new_n968), .B2(G311), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n952), .B2(new_n853), .C1(new_n818), .C2(new_n955), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT48), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n849), .B2(new_n805), .C1(new_n804), .C2(new_n810), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT49), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n278), .B1(new_n970), .B2(G116), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n1026), .B2(new_n1025), .C1(new_n801), .C2(new_n786), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n810), .A2(new_n205), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n278), .B1(new_n805), .B2(new_n364), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n853), .A2(new_n385), .B1(new_n803), .B2(new_n268), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(G150), .C2(new_n825), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n798), .A2(G68), .B1(new_n968), .B2(new_n255), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n210), .C2(new_n794), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1030), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n772), .A2(new_n720), .B1(new_n215), .B2(new_n228), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n255), .A2(new_n385), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n720), .B1(new_n1039), .B2(KEYINPUT50), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n302), .C1(KEYINPUT50), .C2(new_n1039), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n381), .A2(new_n205), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n769), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT114), .Z(new_n1044));
  NOR2_X1   g0844(.A1(new_n243), .A2(new_n302), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1038), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1037), .A2(new_n779), .B1(new_n780), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n703), .B2(new_n782), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n763), .A2(new_n1013), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n717), .B1(new_n763), .B2(new_n1013), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1021), .B1(new_n766), .B2(new_n1048), .C1(new_n1050), .C2(new_n1051), .ZN(G393));
  OAI221_X1 g0852(.A(new_n780), .B1(new_n210), .B2(new_n227), .C1(new_n253), .C2(new_n950), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n808), .A2(G159), .B1(new_n851), .B2(G150), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT51), .Z(new_n1055));
  AOI21_X1  g0855(.A(new_n846), .B1(new_n819), .B2(new_n255), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n876), .A2(new_n968), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n805), .A2(new_n205), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n278), .B1(new_n786), .B2(new_n965), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n266), .C2(new_n828), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n798), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n282), .B1(new_n1062), .B2(new_n804), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1063), .B(new_n815), .C1(G116), .C2(new_n963), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n808), .A2(G311), .B1(new_n851), .B2(G317), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT52), .Z(new_n1066));
  AOI22_X1  g0866(.A1(G283), .A2(new_n828), .B1(new_n825), .B2(G322), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT115), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n790), .A2(new_n955), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1061), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n766), .B1(new_n1071), .B2(new_n779), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1053), .B(new_n1072), .C1(new_n983), .C2(new_n782), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n1049), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n717), .B1(new_n1050), .B2(new_n1006), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1073), .B1(new_n997), .B2(new_n1074), .C1(new_n1075), .C2(new_n1076), .ZN(G390));
  NOR2_X1   g0877(.A1(new_n935), .A2(new_n929), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n916), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT39), .B1(new_n896), .B2(new_n902), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n903), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n704), .B(new_n840), .C1(new_n753), .C2(new_n758), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n933), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT116), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1084), .A2(KEYINPUT116), .A3(new_n933), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1089), .A2(new_n911), .B1(new_n678), .B2(new_n696), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1083), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(G330), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n839), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n910), .B(new_n1094), .C1(new_n744), .C2(new_n747), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1082), .A2(new_n1092), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1094), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n732), .A2(new_n738), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n696), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n672), .A2(new_n547), .A3(new_n555), .A4(new_n740), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1101), .A2(new_n670), .A3(new_n636), .A4(new_n696), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1102), .B2(new_n745), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1098), .B1(new_n1103), .B2(new_n904), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n910), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1078), .B1(new_n926), .B2(new_n928), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n1091), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1097), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n459), .A2(new_n422), .A3(new_n461), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n906), .A2(new_n1109), .A3(new_n377), .A4(new_n1093), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n923), .A2(new_n1110), .A3(new_n686), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1084), .A2(KEYINPUT116), .A3(new_n933), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT116), .B1(new_n1084), .B2(new_n933), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1095), .B1(new_n1104), .B2(new_n910), .ZN(new_n1115));
  OAI21_X1  g0915(.A(KEYINPUT118), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT118), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n911), .B1(new_n906), .B2(new_n1098), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1089), .A2(new_n1117), .A3(new_n1095), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n743), .A2(KEYINPUT31), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n747), .B1(new_n1121), .B2(new_n1100), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n911), .B1(new_n1122), .B2(new_n1098), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1123), .A2(KEYINPUT117), .B1(new_n910), .B2(new_n1104), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT117), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1125), .B(new_n911), .C1(new_n1122), .C2(new_n1098), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n934), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1111), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT119), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT119), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1111), .B(new_n1130), .C1(new_n1120), .C2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1108), .A2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1108), .A2(KEYINPUT120), .A3(new_n1132), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT120), .B1(new_n1108), .B2(new_n1132), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n717), .B(new_n1133), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n777), .B1(new_n926), .B2(new_n928), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G128), .A2(new_n851), .B1(new_n968), .B2(G137), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n268), .B2(new_n805), .C1(new_n864), .C2(new_n853), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT54), .B(G143), .Z(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n819), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(G125), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n278), .B1(new_n786), .B2(new_n1142), .C1(new_n201), .C2(new_n793), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT121), .Z(new_n1144));
  NOR2_X1   g0944(.A1(new_n810), .A2(new_n429), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1141), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n282), .B1(new_n786), .B2(new_n804), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1148), .B(new_n858), .C1(G107), .C2(new_n968), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n803), .A2(new_n849), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1058), .B(new_n1150), .C1(G116), .C2(new_n808), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(new_n219), .C2(new_n811), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n818), .A2(new_n210), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1147), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n779), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n255), .B2(new_n870), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1137), .A2(new_n766), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1108), .B2(new_n1020), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1136), .A2(new_n1158), .ZN(G378));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1111), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1105), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1082), .B2(new_n1092), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1106), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1132), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT120), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1108), .A2(KEYINPUT120), .A3(new_n1132), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1161), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(G330), .B(new_n913), .C1(new_n917), .C2(KEYINPUT40), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n937), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1170), .A2(new_n931), .A3(new_n930), .A4(new_n936), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n459), .A2(new_n461), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT122), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n433), .A2(new_n888), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1178), .B(new_n1179), .Z(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1174), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1172), .A2(new_n1180), .A3(new_n1173), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1160), .B1(new_n1169), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1111), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(KEYINPUT57), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1185), .A2(new_n1188), .A3(new_n717), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1182), .A2(new_n1020), .A3(new_n1183), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n803), .A2(new_n1142), .B1(new_n805), .B2(new_n429), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G132), .A2(new_n968), .B1(new_n828), .B2(new_n1140), .ZN(new_n1192));
  INV_X1    g0992(.A(G137), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n1062), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1191), .B(new_n1194), .C1(G128), .C2(new_n808), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT59), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G41), .B1(new_n825), .B2(G124), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G33), .B1(new_n970), .B2(G159), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n964), .B1(new_n617), .B2(new_n803), .C1(new_n853), .C2(new_n215), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(new_n1200), .A2(G41), .A3(new_n278), .A4(new_n1031), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n790), .A2(new_n210), .B1(new_n793), .B2(new_n208), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G283), .B2(new_n825), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(new_n364), .C2(new_n1062), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT58), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n385), .B1(new_n280), .B2(G41), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1199), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n766), .B1(new_n1207), .B2(new_n779), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n876), .B2(new_n870), .C1(new_n1180), .C2(new_n777), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1190), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1189), .A2(new_n1211), .ZN(G375));
  OAI21_X1  g1012(.A(new_n278), .B1(new_n793), .B2(new_n208), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n853), .A2(new_n1193), .B1(new_n803), .B2(new_n864), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(G50), .C2(new_n963), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n968), .A2(new_n1140), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n812), .A2(G159), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n798), .A2(G150), .B1(G128), .B2(new_n825), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n282), .B1(new_n617), .B2(new_n790), .C1(new_n818), .C2(new_n215), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n851), .A2(G294), .B1(new_n963), .B2(new_n363), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n853), .B2(new_n849), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n794), .A2(new_n205), .B1(new_n811), .B2(new_n210), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n1220), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n825), .A2(G303), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1219), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n779), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(G68), .B2(new_n870), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n766), .B(new_n1228), .C1(new_n911), .C2(new_n776), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1120), .A2(new_n1127), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1229), .B1(new_n1231), .B2(new_n1020), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1129), .B(new_n1131), .C1(new_n1111), .C2(new_n1231), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1232), .B1(new_n1233), .B2(new_n1016), .ZN(G381));
  NAND4_X1  g1034(.A1(new_n1136), .A2(new_n1158), .A3(new_n1190), .A4(new_n1209), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1184), .B1(new_n1236), .B2(new_n1111), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n718), .B1(new_n1237), .B2(KEYINPUT57), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1235), .B1(new_n1238), .B2(new_n1185), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(G387), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1240));
  OR2_X1    g1040(.A1(G393), .A2(G396), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT123), .Z(G407));
  NAND2_X1  g1044(.A1(new_n1239), .A2(new_n695), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(G407), .A2(G213), .A3(new_n1245), .ZN(G409));
  INV_X1    g1046(.A(G396), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(G393), .B(new_n1247), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1248), .A2(KEYINPUT124), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1018), .A2(G390), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1248), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1018), .A2(G390), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1249), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1018), .A2(G390), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1248), .A2(KEYINPUT124), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1255), .A2(new_n1256), .A3(new_n1250), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1169), .A2(new_n1016), .A3(new_n1184), .ZN(new_n1260));
  INV_X1    g1060(.A(G213), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1235), .A2(new_n1260), .B1(new_n1261), .B2(G343), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G375), .B2(G378), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT60), .B1(new_n1230), .B2(new_n1161), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1233), .B2(KEYINPUT60), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n717), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1232), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n872), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(G384), .A3(new_n1232), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1261), .A2(G343), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(G2897), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1270), .A2(G2897), .A3(new_n1272), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1258), .B(new_n1259), .C1(new_n1263), .C2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT63), .B1(new_n1263), .B2(new_n1271), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1235), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1237), .A2(new_n1015), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1272), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1210), .B1(new_n1238), .B2(new_n1185), .ZN(new_n1283));
  INV_X1    g1083(.A(G378), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1282), .B(new_n1271), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT63), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT125), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1263), .A2(new_n1288), .A3(KEYINPUT63), .A4(new_n1271), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1279), .A2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1258), .A2(KEYINPUT127), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1254), .A2(new_n1257), .A3(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1284), .B1(new_n1189), .B2(new_n1211), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1274), .B(new_n1275), .C1(new_n1296), .C2(new_n1262), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1296), .A2(new_n1262), .A3(new_n1270), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT62), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1297), .B(new_n1259), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1301));
  XOR2_X1   g1101(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1302));
  NOR2_X1   g1102(.A1(new_n1285), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1295), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1291), .A2(new_n1304), .ZN(G405));
  OR3_X1    g1105(.A1(new_n1296), .A2(new_n1239), .A3(new_n1271), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1271), .B1(new_n1296), .B2(new_n1239), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1308), .B(new_n1258), .ZN(G402));
endmodule


