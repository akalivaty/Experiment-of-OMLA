//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046;
  XNOR2_X1  g000(.A(G134gat), .B(G162gat), .ZN(new_n202));
  AOI21_X1  g001(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G190gat), .B(G218gat), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT14), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G50gat), .ZN(new_n217));
  INV_X1    g016(.A(G50gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G43gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n215), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT15), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G29gat), .A2(G36gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(KEYINPUT14), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n212), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n218), .A2(G43gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n216), .A2(G50gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n221), .B1(new_n231), .B2(KEYINPUT15), .ZN(new_n232));
  AND2_X1   g031(.A1(KEYINPUT90), .A2(G85gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(KEYINPUT90), .A2(G85gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G92gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n235), .A2(new_n236), .B1(KEYINPUT8), .B2(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n237), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT91), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(KEYINPUT91), .A3(new_n237), .ZN(new_n243));
  NAND2_X1  g042(.A1(G85gat), .A2(G92gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT7), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(G85gat), .A3(G92gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n238), .A2(new_n242), .A3(new_n243), .A4(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(KEYINPUT90), .A2(G85gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(KEYINPUT90), .A2(G85gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n236), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT8), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n248), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n241), .A3(new_n240), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n232), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT93), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n256), .B(KEYINPUT92), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n224), .A2(new_n212), .B1(new_n227), .B2(new_n228), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT84), .B1(new_n227), .B2(new_n228), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n226), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT15), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT17), .ZN(new_n266));
  INV_X1    g065(.A(new_n221), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT15), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(new_n225), .B2(new_n230), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT17), .B1(new_n270), .B2(new_n221), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n261), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n207), .B1(new_n260), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n259), .A2(KEYINPUT93), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT93), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n257), .B2(new_n258), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n272), .B(new_n207), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n205), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n206), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(new_n204), .A3(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(G155gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G183gat), .B(G211gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT89), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n285), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G57gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G64gat), .ZN(new_n291));
  INV_X1    g090(.A(G64gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G57gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT9), .ZN(new_n294));
  NAND2_X1  g093(.A1(G71gat), .A2(G78gat), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n291), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT86), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(G71gat), .A2(G78gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(KEYINPUT86), .A2(G71gat), .A3(G78gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n295), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n296), .A2(KEYINPUT87), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT87), .B1(new_n296), .B2(new_n304), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G231gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n307), .A2(new_n310), .A3(new_n308), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G127gat), .ZN(new_n315));
  INV_X1    g114(.A(G1gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT16), .ZN(new_n317));
  INV_X1    g116(.A(G15gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G22gat), .ZN(new_n319));
  INV_X1    g118(.A(G22gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G15gat), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n317), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(G1gat), .B1(new_n319), .B2(new_n321), .ZN(new_n323));
  OAI21_X1  g122(.A(G8gat), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n320), .A2(G15gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n318), .A2(G22gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n316), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G8gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n317), .A2(new_n319), .A3(new_n321), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n291), .A2(new_n293), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n295), .A2(new_n294), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n304), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT87), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n296), .A2(KEYINPUT87), .A3(new_n304), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n302), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n331), .B1(new_n338), .B2(KEYINPUT21), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G127gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n312), .A2(new_n341), .A3(new_n313), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n315), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n340), .B1(new_n315), .B2(new_n342), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n289), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n345), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(new_n343), .A3(new_n288), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n283), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT94), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT94), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n283), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  XNOR2_X1  g152(.A(G120gat), .B(G148gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT96), .ZN(new_n355));
  XNOR2_X1  g154(.A(G176gat), .B(G204gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G230gat), .ZN(new_n359));
  INV_X1    g158(.A(G233gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n254), .A2(KEYINPUT95), .A3(new_n240), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n254), .A2(KEYINPUT95), .ZN(new_n364));
  INV_X1    g163(.A(new_n240), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n338), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n336), .A2(new_n337), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n368), .A2(new_n303), .B1(new_n249), .B2(new_n255), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n362), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n256), .A2(new_n338), .A3(KEYINPUT10), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n361), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n361), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n367), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n358), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT97), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n338), .A2(new_n363), .A3(new_n366), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n256), .A2(new_n307), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT10), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n371), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n373), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n374), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(new_n357), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n375), .A2(new_n376), .A3(new_n383), .ZN(new_n384));
  OAI211_X1 g183(.A(KEYINPUT97), .B(new_n358), .C1(new_n372), .C2(new_n374), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n351), .A2(new_n353), .A3(new_n386), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n387), .A2(KEYINPUT98), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(KEYINPUT98), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(KEYINPUT24), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT23), .ZN(new_n396));
  INV_X1    g195(.A(G169gat), .ZN(new_n397));
  INV_X1    g196(.A(G176gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G183gat), .ZN(new_n402));
  INV_X1    g201(.A(G190gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(KEYINPUT24), .A3(new_n393), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT25), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n395), .A2(new_n401), .A3(new_n405), .A4(KEYINPUT25), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT64), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT27), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n411), .B(new_n403), .C1(new_n412), .C2(G183gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT28), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(G190gat), .B1(new_n402), .B2(KEYINPUT27), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(G183gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n416), .A2(KEYINPUT64), .A3(new_n414), .A4(new_n417), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(G169gat), .B2(G176gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n423), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n419), .A2(new_n420), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n391), .B1(new_n410), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n394), .B1(new_n400), .B2(new_n399), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT25), .B1(new_n427), .B2(new_n405), .ZN(new_n428));
  AND4_X1   g227(.A1(KEYINPUT25), .A2(new_n395), .A3(new_n401), .A4(new_n405), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n426), .B1(new_n432), .B2(new_n391), .ZN(new_n433));
  XNOR2_X1  g232(.A(G211gat), .B(G218gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n436));
  OR2_X1    g235(.A1(G197gat), .A2(G204gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(G197gat), .A2(G204gat), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT68), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G211gat), .A2(G218gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT22), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(G197gat), .A2(G204gat), .ZN(new_n445));
  AND2_X1   g244(.A1(G197gat), .A2(G204gat), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(KEYINPUT68), .A3(new_n434), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n433), .A2(KEYINPUT70), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n391), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n430), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT29), .B1(new_n410), .B2(new_n425), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n453), .B(new_n450), .C1(new_n454), .C2(new_n452), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT70), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n420), .A2(new_n422), .A3(new_n424), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n408), .A2(new_n409), .B1(new_n458), .B2(new_n419), .ZN(new_n459));
  XOR2_X1   g258(.A(KEYINPUT69), .B(KEYINPUT29), .Z(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n391), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n450), .B1(new_n462), .B2(new_n453), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n451), .B1(new_n457), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G8gat), .B(G36gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(G64gat), .B(G92gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n465), .B(new_n466), .Z(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(KEYINPUT30), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT71), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT71), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n464), .A2(new_n470), .A3(KEYINPUT30), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT30), .B1(new_n464), .B2(new_n467), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n464), .A2(new_n467), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(G120gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(G113gat), .ZN(new_n478));
  INV_X1    g277(.A(G113gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G120gat), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT1), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(G127gat), .A2(G134gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(G127gat), .A2(G134gat), .ZN(new_n483));
  OAI22_X1  g282(.A1(new_n482), .A2(new_n483), .B1(KEYINPUT65), .B2(KEYINPUT1), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT1), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n479), .A2(G120gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n477), .A2(G113gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n490));
  INV_X1    g289(.A(G134gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n341), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G127gat), .A2(G134gat), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G148gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G141gat), .ZN(new_n497));
  INV_X1    g296(.A(G141gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G148gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G155gat), .B(G162gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(G155gat), .A2(G162gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT2), .ZN(new_n503));
  AND4_X1   g302(.A1(KEYINPUT72), .A2(new_n500), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT72), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n505), .B1(new_n497), .B2(new_n499), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n501), .B1(new_n506), .B2(new_n503), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n485), .B(new_n495), .C1(new_n504), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n501), .A3(new_n503), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n498), .A2(G148gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n496), .A2(G141gat), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT72), .B(new_n503), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n501), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n489), .A2(new_n494), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n481), .A2(new_n484), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n509), .B(new_n514), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G225gat), .A2(G233gat), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT73), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT5), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n508), .B2(new_n517), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT73), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n514), .A2(new_n509), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT3), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT3), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n514), .A2(new_n527), .A3(new_n509), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n495), .A2(new_n485), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n529), .A2(KEYINPUT4), .A3(new_n509), .A4(new_n514), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n531), .A2(new_n532), .A3(new_n534), .A4(new_n519), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n524), .A3(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n534), .A2(new_n532), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n537), .A2(new_n521), .A3(new_n519), .A4(new_n531), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G1gat), .B(G29gat), .Z(new_n540));
  XNOR2_X1  g339(.A(G57gat), .B(G85gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT40), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n537), .A2(new_n531), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT39), .ZN(new_n550));
  INV_X1    g349(.A(new_n519), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n544), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n518), .A2(new_n519), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT39), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n551), .B2(new_n549), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n548), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n549), .A2(new_n551), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT39), .A3(new_n554), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n559), .A2(KEYINPUT40), .A3(new_n544), .A4(new_n552), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n544), .B1(new_n536), .B2(new_n538), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT81), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND4_X1   g362(.A1(new_n547), .A2(new_n557), .A3(new_n560), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n476), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G228gat), .A2(G233gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n528), .A2(new_n460), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n450), .B1(new_n567), .B2(KEYINPUT79), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT79), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n528), .A2(new_n569), .A3(new_n460), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n441), .A2(new_n431), .A3(new_n448), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n441), .A2(new_n448), .A3(KEYINPUT77), .A4(new_n431), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n527), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT78), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n576), .A2(new_n577), .A3(new_n525), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n577), .B1(new_n576), .B2(new_n525), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n571), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n461), .B1(new_n447), .B2(new_n434), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT76), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n435), .A2(new_n439), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n527), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n582), .B1(new_n581), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n525), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n567), .A2(new_n449), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n566), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n580), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(G22gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT80), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n580), .A2(new_n320), .A3(new_n590), .ZN(new_n594));
  XOR2_X1   g393(.A(G78gat), .B(G106gat), .Z(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT31), .B(G50gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(KEYINPUT80), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n600), .A2(new_n597), .B1(new_n592), .B2(new_n594), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n467), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT37), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n462), .A2(new_n453), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n604), .B1(new_n605), .B2(new_n450), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n433), .A2(new_n449), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT38), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT82), .B1(new_n464), .B2(new_n604), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT82), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n452), .B1(new_n430), .B2(new_n460), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n449), .B1(new_n611), .B2(new_n426), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(new_n456), .A3(new_n455), .ZN(new_n613));
  AOI211_X1 g412(.A(new_n610), .B(KEYINPUT37), .C1(new_n613), .C2(new_n451), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n603), .B(new_n608), .C1(new_n609), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n561), .A2(KEYINPUT6), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n536), .A2(new_n544), .A3(new_n538), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT6), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n547), .A2(new_n619), .A3(new_n563), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n615), .A2(new_n616), .A3(new_n474), .A4(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT38), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n452), .B1(new_n430), .B2(new_n431), .ZN(new_n623));
  NOR4_X1   g422(.A1(new_n623), .A2(new_n426), .A3(new_n456), .A4(new_n449), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT70), .B1(new_n433), .B2(new_n450), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n624), .B1(new_n625), .B2(new_n612), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n610), .B1(new_n626), .B2(KEYINPUT37), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n464), .A2(KEYINPUT82), .A3(new_n604), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n467), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(KEYINPUT37), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n622), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n565), .B(new_n602), .C1(new_n621), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n600), .A2(new_n597), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n592), .A2(new_n594), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n598), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n618), .B(new_n617), .C1(new_n561), .C2(KEYINPUT75), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n539), .A2(KEYINPUT75), .A3(new_n545), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n616), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n475), .A3(new_n472), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(KEYINPUT67), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n430), .A2(new_n529), .ZN(new_n644));
  INV_X1    g443(.A(G227gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n360), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n410), .A2(new_n530), .A3(new_n425), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT66), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n644), .A2(KEYINPUT66), .A3(new_n646), .A4(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n644), .A2(new_n647), .ZN(new_n655));
  INV_X1    g454(.A(new_n646), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT34), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n646), .B1(new_n644), .B2(new_n647), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT34), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(G15gat), .B(G43gat), .Z(new_n663));
  XNOR2_X1  g462(.A(G71gat), .B(G99gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n654), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n659), .B(KEYINPUT34), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT33), .B1(new_n650), .B2(new_n651), .ZN(new_n668));
  INV_X1    g467(.A(new_n665), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n652), .A2(KEYINPUT32), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n666), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n666), .B2(new_n670), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n643), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n662), .B1(new_n654), .B2(new_n665), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n666), .A2(new_n670), .A3(new_n672), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT67), .B(KEYINPUT36), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n636), .A2(new_n640), .B1(new_n675), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n635), .A2(new_n678), .A3(new_n598), .A4(new_n679), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT35), .B1(new_n684), .B2(new_n640), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT35), .B1(new_n620), .B2(new_n616), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n673), .A2(new_n674), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n469), .A2(new_n471), .B1(new_n474), .B2(new_n473), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n602), .A2(new_n686), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n632), .A2(new_n683), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n322), .A2(new_n323), .A3(G8gat), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n328), .B1(new_n327), .B2(new_n329), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n271), .A2(new_n268), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT85), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n232), .B2(new_n331), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n271), .A2(new_n268), .A3(new_n695), .A4(new_n693), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(G229gat), .A2(G233gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT18), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n693), .B1(new_n270), .B2(new_n221), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n265), .A2(new_n331), .A3(new_n267), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n700), .B(KEYINPUT13), .Z(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n700), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n697), .B2(new_n698), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(KEYINPUT18), .ZN(new_n712));
  XNOR2_X1  g511(.A(G113gat), .B(G141gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT83), .B(G197gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT11), .B(G169gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT12), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n703), .A2(new_n712), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n703), .B2(new_n712), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n690), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n390), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n639), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT99), .B(G1gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1324gat));
  NOR2_X1   g525(.A1(new_n723), .A2(new_n688), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT16), .B(G8gat), .Z(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n727), .B2(new_n328), .ZN(new_n730));
  MUX2_X1   g529(.A(new_n729), .B(new_n730), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g530(.A1(new_n675), .A2(new_n682), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G15gat), .B1(new_n723), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n687), .A2(new_n318), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n723), .B2(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT101), .Z(G1326gat));
  NOR3_X1   g538(.A1(new_n690), .A2(new_n602), .A3(new_n721), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n390), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT43), .B(G22gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1327gat));
  NOR2_X1   g542(.A1(new_n690), .A2(new_n283), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n384), .A2(new_n385), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n721), .A2(new_n745), .A3(new_n349), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n639), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n208), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n632), .A2(new_n683), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n685), .A2(new_n689), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n283), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n690), .B2(new_n283), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n746), .ZN(new_n759));
  OAI21_X1  g558(.A(G29gat), .B1(new_n759), .B2(new_n639), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n750), .A2(new_n760), .ZN(G1328gat));
  NAND3_X1  g560(.A1(new_n747), .A2(new_n209), .A3(new_n476), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT102), .B(KEYINPUT46), .Z(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G36gat), .B1(new_n759), .B2(new_n688), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1329gat));
  OAI21_X1  g565(.A(G43gat), .B1(new_n759), .B2(new_n735), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n747), .A2(new_n216), .A3(new_n687), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G43gat), .B1(new_n759), .B2(new_n732), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(new_n769), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n772), .B2(new_n768), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT103), .ZN(G1330gat));
  OAI21_X1  g573(.A(G50gat), .B1(new_n759), .B2(new_n602), .ZN(new_n775));
  NOR4_X1   g574(.A1(new_n283), .A2(new_n745), .A3(new_n349), .A4(G50gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n740), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g578(.A1(new_n351), .A2(new_n721), .A3(new_n353), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n690), .A2(new_n386), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n748), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n476), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT49), .B(G64gat), .Z(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(G1333gat));
  INV_X1    g586(.A(new_n735), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n673), .A2(new_n674), .A3(G71gat), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n789), .A2(G71gat), .B1(new_n781), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g591(.A1(new_n781), .A2(new_n636), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G78gat), .ZN(G1335gat));
  INV_X1    g593(.A(new_n718), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n711), .A2(KEYINPUT18), .ZN(new_n796));
  INV_X1    g595(.A(new_n709), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n711), .A2(KEYINPUT18), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n703), .A2(new_n712), .A3(new_n718), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(new_n349), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n753), .A2(new_n754), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n744), .A2(KEYINPUT51), .A3(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n808), .A2(KEYINPUT104), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n804), .A2(KEYINPUT104), .A3(new_n805), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n748), .A2(new_n235), .A3(new_n745), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n802), .A2(new_n349), .A3(new_n386), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n758), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n639), .ZN(new_n815));
  OAI22_X1  g614(.A1(new_n811), .A2(new_n812), .B1(new_n235), .B2(new_n815), .ZN(G1336gat));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817));
  OAI21_X1  g616(.A(G92gat), .B1(new_n814), .B2(new_n688), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n476), .A2(new_n745), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(G92gat), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n817), .B(new_n818), .C1(new_n811), .C2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT105), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n823), .B1(new_n825), .B2(KEYINPUT52), .ZN(new_n826));
  AOI211_X1 g625(.A(KEYINPUT105), .B(new_n817), .C1(new_n818), .C2(new_n824), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n822), .B1(new_n826), .B2(new_n827), .ZN(G1337gat));
  OAI21_X1  g627(.A(G99gat), .B1(new_n814), .B2(new_n735), .ZN(new_n829));
  INV_X1    g628(.A(G99gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n687), .A2(new_n830), .A3(new_n745), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n811), .B2(new_n831), .ZN(G1338gat));
  NOR3_X1   g631(.A1(new_n602), .A2(G106gat), .A3(new_n386), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n809), .A2(new_n810), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n755), .A2(new_n757), .A3(new_n636), .A4(new_n813), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G106gat), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT107), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n837), .A2(KEYINPUT106), .B1(new_n808), .B2(new_n833), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT106), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n841), .A3(G106gat), .ZN(new_n842));
  AOI211_X1 g641(.A(new_n839), .B(new_n835), .C1(new_n840), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n837), .A2(KEYINPUT106), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n808), .A2(new_n833), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT107), .B1(new_n846), .B2(KEYINPUT53), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n838), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT108), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT108), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(new_n838), .C1(new_n843), .C2(new_n847), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(G1339gat));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n370), .A2(new_n361), .A3(new_n371), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n381), .A3(KEYINPUT54), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n857), .B(new_n373), .C1(new_n379), .C2(new_n380), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n358), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n853), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n855), .A2(KEYINPUT55), .A3(new_n358), .A4(new_n858), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n383), .A3(new_n861), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n697), .A2(new_n710), .A3(new_n698), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n704), .A2(new_n705), .A3(new_n708), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT109), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n717), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT110), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT109), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n864), .B(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n697), .A2(new_n710), .A3(new_n698), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(KEYINPUT110), .A3(new_n717), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n801), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n721), .A2(new_n862), .B1(new_n874), .B2(new_n386), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n283), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n383), .ZN(new_n877));
  INV_X1    g676(.A(new_n859), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT55), .B1(new_n878), .B2(new_n855), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT110), .B1(new_n872), .B2(new_n717), .ZN(new_n881));
  INV_X1    g680(.A(new_n717), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n867), .B(new_n882), .C1(new_n870), .C2(new_n871), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n754), .A2(new_n801), .A3(new_n880), .A4(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n349), .B1(new_n876), .B2(new_n885), .ZN(new_n886));
  AND4_X1   g685(.A1(new_n721), .A2(new_n351), .A3(new_n353), .A4(new_n386), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT111), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n349), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n880), .A2(new_n802), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n745), .A2(new_n884), .A3(new_n801), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n754), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n283), .A2(new_n862), .A3(new_n874), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n351), .A2(new_n721), .A3(new_n353), .A4(new_n386), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT111), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n476), .A2(new_n639), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n898), .A2(new_n602), .A3(new_n687), .A4(new_n899), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT112), .Z(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(new_n479), .A3(new_n721), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n888), .B1(new_n886), .B2(new_n887), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n895), .A2(KEYINPUT111), .A3(new_n896), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(new_n639), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n684), .A2(new_n476), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(G113gat), .B1(new_n909), .B2(new_n802), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n902), .A2(new_n910), .ZN(G1340gat));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n477), .A3(new_n745), .ZN(new_n912));
  OAI21_X1  g711(.A(G120gat), .B1(new_n901), .B2(new_n386), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT113), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(G1341gat));
  OAI21_X1  g716(.A(G127gat), .B1(new_n901), .B2(new_n890), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n909), .A2(new_n341), .A3(new_n349), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1342gat));
  OAI21_X1  g719(.A(G134gat), .B1(new_n901), .B2(new_n283), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT114), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n491), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n283), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n921), .A2(new_n927), .ZN(G1343gat));
  XOR2_X1   g727(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n929));
  NAND2_X1  g728(.A1(new_n735), .A2(new_n636), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n906), .A2(new_n688), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n802), .A2(new_n498), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n903), .A2(new_n636), .A3(new_n904), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT57), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT115), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n885), .B1(new_n893), .B2(new_n936), .ZN(new_n937));
  AOI211_X1 g736(.A(KEYINPUT115), .B(new_n754), .C1(new_n891), .C2(new_n892), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n890), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n896), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n602), .A2(new_n935), .ZN(new_n941));
  AOI22_X1  g740(.A1(new_n934), .A2(new_n935), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n732), .ZN(new_n943));
  INV_X1    g742(.A(new_n899), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n942), .A2(new_n721), .A3(new_n946), .ZN(new_n947));
  OAI221_X1 g746(.A(new_n929), .B1(new_n932), .B2(new_n933), .C1(new_n947), .C2(new_n498), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n935), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n940), .A2(new_n941), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT116), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n953), .A3(new_n945), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT116), .B1(new_n942), .B2(new_n946), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n955), .A3(new_n802), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n949), .B1(new_n956), .B2(G141gat), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT58), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n948), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT118), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g760(.A(KEYINPUT118), .B(new_n948), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1344gat));
  XNOR2_X1  g762(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n388), .A2(new_n721), .A3(new_n389), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n636), .B1(new_n965), .B2(new_n886), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(new_n935), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n898), .A2(new_n941), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n946), .A2(new_n386), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(KEYINPUT120), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G148gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT120), .B1(new_n969), .B2(new_n970), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n964), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n496), .A2(KEYINPUT59), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n954), .A2(new_n955), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n386), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n745), .A2(new_n496), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n932), .B2(new_n979), .ZN(G1345gat));
  OAI21_X1  g779(.A(G155gat), .B1(new_n976), .B2(new_n890), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n890), .A2(G155gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n932), .B2(new_n982), .ZN(G1346gat));
  INV_X1    g782(.A(G162gat), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n976), .A2(new_n984), .A3(new_n283), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n932), .A2(new_n283), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n984), .B2(new_n986), .ZN(G1347gat));
  NOR2_X1   g786(.A1(new_n748), .A2(new_n688), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT122), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n898), .A2(new_n602), .A3(new_n687), .A4(new_n989), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n990), .A2(new_n397), .A3(new_n721), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT121), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n898), .A2(new_n992), .A3(new_n639), .ZN(new_n993));
  OAI21_X1  g792(.A(KEYINPUT121), .B1(new_n905), .B2(new_n748), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n684), .A2(new_n688), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(new_n802), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n991), .B1(new_n999), .B2(new_n397), .ZN(G1348gat));
  NOR3_X1   g799(.A1(new_n990), .A2(new_n398), .A3(new_n386), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n998), .A2(new_n745), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n1001), .B1(new_n1002), .B2(new_n398), .ZN(G1349gat));
  OAI21_X1  g802(.A(G183gat), .B1(new_n990), .B2(new_n890), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n402), .A2(KEYINPUT27), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n349), .A2(new_n1005), .A3(new_n417), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1004), .B1(new_n997), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1007), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g807(.A(G190gat), .B1(new_n990), .B2(new_n283), .ZN(new_n1009));
  XNOR2_X1  g808(.A(new_n1009), .B(KEYINPUT61), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n998), .A2(new_n403), .A3(new_n754), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1351gat));
  NAND2_X1  g811(.A1(new_n735), .A2(new_n989), .ZN(new_n1013));
  XNOR2_X1  g812(.A(new_n1013), .B(KEYINPUT124), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n969), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g814(.A(G197gat), .ZN(new_n1016));
  NOR3_X1   g815(.A1(new_n1015), .A2(new_n1016), .A3(new_n721), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n995), .A2(new_n476), .A3(new_n931), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT123), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g819(.A(new_n930), .B1(new_n993), .B2(new_n994), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1021), .A2(KEYINPUT123), .A3(new_n476), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1023), .A2(new_n802), .ZN(new_n1024));
  AOI21_X1  g823(.A(new_n1017), .B1(new_n1024), .B2(new_n1016), .ZN(G1352gat));
  NOR2_X1   g824(.A1(new_n819), .A2(G204gat), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1021), .A2(new_n1026), .ZN(new_n1027));
  OR2_X1    g826(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1028));
  OAI21_X1  g827(.A(G204gat), .B1(new_n1015), .B2(new_n386), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1030));
  NAND3_X1  g829(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(G1353gat));
  INV_X1    g830(.A(G211gat), .ZN(new_n1032));
  NOR2_X1   g831(.A1(new_n1013), .A2(new_n890), .ZN(new_n1033));
  AOI21_X1  g832(.A(new_n1032), .B1(new_n969), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g833(.A(new_n1034), .B(KEYINPUT63), .ZN(new_n1035));
  NAND3_X1  g834(.A1(new_n1023), .A2(new_n1032), .A3(new_n349), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1035), .A2(new_n1036), .ZN(G1354gat));
  NAND2_X1  g836(.A1(new_n754), .A2(G218gat), .ZN(new_n1038));
  XNOR2_X1  g837(.A(new_n1038), .B(KEYINPUT126), .ZN(new_n1039));
  NOR2_X1   g838(.A1(new_n1015), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n754), .ZN(new_n1041));
  INV_X1    g840(.A(KEYINPUT125), .ZN(new_n1042));
  INV_X1    g841(.A(G218gat), .ZN(new_n1043));
  NAND3_X1  g842(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g843(.A(new_n283), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1045));
  OAI21_X1  g844(.A(KEYINPUT125), .B1(new_n1045), .B2(G218gat), .ZN(new_n1046));
  AOI21_X1  g845(.A(new_n1040), .B1(new_n1044), .B2(new_n1046), .ZN(G1355gat));
endmodule


